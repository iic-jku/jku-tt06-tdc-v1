** sch_path: /foss/designs/sim/tb_tt06_tdc.sch
**.subckt tb_tt06_tdc
x1 start stop res[0] res[14] res[16] res[19] res[20] res[21] res[22] res[23] res[24] res[25] res[26] res[27] res[28] res[2]
+ res[32] res[35] res[37] res[38] res[3] res[40] res[41] res[42] res[43] res[44] res[45] res[49] res[50] res[51] res[53] res[54] res[56]
+ res[57] res[59] res[5] res[60] res[61] res[62] res[6] res[7] res[8] res[46] res[11] res[48] res[29] res[34] res[31] res[13] res[18]
+ res[10] res[58] res[63] res[55] res[47] res[52] res[39] res[36] res[33] res[30] res[15] res[12] res[17] res[4] res[9] VDD res[1] GND tdc
VDAC start GND 0 pwl(0 0 500n 0 500.1n 1.8)
.save v(start)
VDAC1 stop GND 0 pwl(0 0 508n 0 508.1n 1.8)
.save v(stop)
Cload[65] res[65] GND 10f m=1
Cload[64] res[64] GND 10f m=1
Cload[63] res[63] GND 10f m=1
Cload[62] res[62] GND 10f m=1
Cload[61] res[61] GND 10f m=1
Cload[60] res[60] GND 10f m=1
Cload[59] res[59] GND 10f m=1
Cload[58] res[58] GND 10f m=1
Cload[57] res[57] GND 10f m=1
Cload[56] res[56] GND 10f m=1
Cload[55] res[55] GND 10f m=1
Cload[54] res[54] GND 10f m=1
Cload[53] res[53] GND 10f m=1
Cload[52] res[52] GND 10f m=1
Cload[51] res[51] GND 10f m=1
Cload[50] res[50] GND 10f m=1
Cload[49] res[49] GND 10f m=1
Cload[48] res[48] GND 10f m=1
Cload[47] res[47] GND 10f m=1
Cload[46] res[46] GND 10f m=1
Cload[45] res[45] GND 10f m=1
Cload[44] res[44] GND 10f m=1
Cload[43] res[43] GND 10f m=1
Cload[42] res[42] GND 10f m=1
Cload[41] res[41] GND 10f m=1
Cload[40] res[40] GND 10f m=1
Cload[39] res[39] GND 10f m=1
Cload[38] res[38] GND 10f m=1
Cload[37] res[37] GND 10f m=1
Cload[36] res[36] GND 10f m=1
Cload[35] res[35] GND 10f m=1
Cload[34] res[34] GND 10f m=1
Cload[33] res[33] GND 10f m=1
Cload[32] res[32] GND 10f m=1
Cload[31] res[31] GND 10f m=1
Cload[30] res[30] GND 10f m=1
Cload[29] res[29] GND 10f m=1
Cload[28] res[28] GND 10f m=1
Cload[27] res[27] GND 10f m=1
Cload[26] res[26] GND 10f m=1
Cload[25] res[25] GND 10f m=1
Cload[24] res[24] GND 10f m=1
Cload[23] res[23] GND 10f m=1
Cload[22] res[22] GND 10f m=1
Cload[21] res[21] GND 10f m=1
Cload[20] res[20] GND 10f m=1
Cload[19] res[19] GND 10f m=1
Cload[18] res[18] GND 10f m=1
Cload[17] res[17] GND 10f m=1
Cload[16] res[16] GND 10f m=1
Cload[15] res[15] GND 10f m=1
Cload[14] res[14] GND 10f m=1
Cload[13] res[13] GND 10f m=1
Cload[12] res[12] GND 10f m=1
Cload[11] res[11] GND 10f m=1
Cload[10] res[10] GND 10f m=1
Cload[9] res[9] GND 10f m=1
Cload[8] res[8] GND 10f m=1
Cload[7] res[7] GND 10f m=1
Cload[6] res[6] GND 10f m=1
Cload[5] res[5] GND 10f m=1
Cload[4] res[4] GND 10f m=1
Cload[3] res[3] GND 10f m=1
Cload[2] res[2] GND 10f m=1
Cload[1] res[1] GND 10f m=1
Cload[0] res[0] GND 10f m=1
.save v(res[65])
.save v(res[64])
.save v(res[63])
.save v(res[62])
.save v(res[61])
.save v(res[60])
.save v(res[59])
.save v(res[58])
.save v(res[57])
.save v(res[56])
.save v(res[55])
.save v(res[54])
.save v(res[53])
.save v(res[52])
.save v(res[51])
.save v(res[50])
.save v(res[49])
.save v(res[48])
.save v(res[47])
.save v(res[46])
.save v(res[45])
.save v(res[44])
.save v(res[43])
.save v(res[42])
.save v(res[41])
.save v(res[40])
.save v(res[39])
.save v(res[38])
.save v(res[37])
.save v(res[36])
.save v(res[35])
.save v(res[34])
.save v(res[33])
.save v(res[32])
.save v(res[31])
.save v(res[30])
.save v(res[29])
.save v(res[28])
.save v(res[27])
.save v(res[26])
.save v(res[25])
.save v(res[24])
.save v(res[23])
.save v(res[22])
.save v(res[21])
.save v(res[20])
.save v(res[19])
.save v(res[18])
.save v(res[17])
.save v(res[16])
.save v(res[15])
.save v(res[14])
.save v(res[13])
.save v(res[12])
.save v(res[11])
.save v(res[10])
.save v(res[9])
.save v(res[8])
.save v(res[7])
.save v(res[6])
.save v(res[5])
.save v(res[4])
.save v(res[3])
.save v(res[2])
.save v(res[1])
.save v(res[0])
.save v(vdd)
VDAC2 VDD GND 0 pwl(0 0 100n 1.8)
**** begin user architecture code



* ngspice commands
****************

.save v(x1.w_dly_sig[0])
.save v(x1.w_dly_sig[1])
.save v(x1.w_dly_sig[2])
.save v(x1.w_dly_sig[3])
.save v(x1.w_dly_sig[4])
.save v(x1.w_dly_sig[5])
.save v(x1.w_dly_sig[6])
.save v(x1.w_dly_sig[7])
.save v(x1.w_dly_sig[8])
.save v(x1.w_dly_sig[9])
.save v(x1.w_dly_sig[10])
.save v(x1.w_dly_sig[11])
.save v(x1.w_dly_sig[12])
.save v(x1.w_dly_sig[13])
.save v(x1.w_dly_sig[14])
.save v(x1.w_dly_sig[15])
.save v(x1.w_dly_sig[16])
.save v(x1.w_dly_sig[17])
.save v(x1.w_dly_sig[18])
.save v(x1.w_dly_sig[19])
.save v(x1.w_dly_sig[20])
.save v(x1.w_dly_sig[21])

****************
* Misc
****************
.param fclk=10MEG
.options method=gear maxord=2
.temp 30

.control
set num_threads=6
tran 0.01n 600n

write tb_tt06_tdc.raw

*exit
.endc




** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  tdc.sym # of pins=5
** sym_path: /foss/designs/sim/tdc.sym
.include tdc.pex.spice
.GLOBAL VDD
.GLOBAL GND
.end
