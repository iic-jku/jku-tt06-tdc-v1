* PEX produced on Thu Mar 14 08:36:32 AM CET 2024 using /foss/tools/osic-multitool/iic-pex.sh with m=1 and s=1
* NGSPICE file created from tt_um_hpretl_tt06_tdc.ext - technology: sky130A

.subckt tt_um_hpretl_tt06_tdc clk ena rst_n ui_in[1] ui_in[2] ui_in[5] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[1]
+ uio_oe[3] uio_oe[4] uio_oe[6] uio_oe[7] uio_out[3] uio_out[4] uio_out[6] uio_out[7]
+ uo_out[4] ui_in[0] ui_in[4] uio_oe[0] ui_in[6] uio_out[1] uio_out[0] uo_out[3] uio_out[5]
+ uio_oe[5] uio_out[2] uo_out[2] uio_oe[2] uo_out[1] uo_out[0] uo_out[7] ui_in[3]
+ uo_out[6] uo_out[5] VGND VPWR
X0 a_9135_5487# _028_ a_9217_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR a_7470_17732# a_7399_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2 VGND tdc0.w_dly_sig\[38\] tdc0.w_dly_sig_n\[38\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_12134_6549# _010_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND _054_ a_10883_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 VPWR tdc0.w_dly_sig_n\[0\] tdc0.w_dly_sig\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_8879_11989# a_8795_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7 a_10774_15101# a_10527_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X8 a_8561_9129# a_7571_8757# a_8435_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9 VGND a_17555_6807# tdc0.o_result\[116\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 VGND tdc0.w_dly_sig_n\[33\] tdc0.w_dly_sig_n\[35\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_2290_2879# a_2122_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12 tdc0.w_dly_sig\[51\] tdc0.w_dly_sig_n\[50\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 tdc0.w_dly_sig_n\[67\] tdc0.w_dly_sig_n\[65\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_13353_8207# a_13176_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X16 tdc0.o_result\[82\] a_2715_1109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 tdc0.w_dly_sig_n\[68\] tdc0.w_dly_sig_n\[66\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X18 a_17033_8751# tdc0.w_dly_sig\[118\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X19 a_15374_13103# a_15127_13481# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X21 VPWR clknet_4_3_0_clk a_7019_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X22 VGND tdc0.w_dly_sig_n\[69\] tdc0.w_dly_sig_n\[71\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_13817_9545# tdc0.o_result\[28\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X24 tdc0.w_dly_sig_n\[7\] tdc0.w_dly_sig\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X25 a_15462_15101# a_15189_14735# a_15377_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X27 a_1573_6581# a_1407_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X29 a_10759_8181# _004_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X30 a_17739_4631# a_17835_4631# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X31 net3 a_10423_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X32 VGND a_16733_5461# _064_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X33 a_12117_8457# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X34 tdc0.w_dly_sig\[40\] tdc0.w_dly_sig_n\[39\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 clknet_4_11_0_clk a_16762_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 a_16762_8207# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X37 a_11504_11445# _056_ a_11892_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 VGND a_3698_12559# clknet_4_4_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X40 a_9374_14165# a_9206_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X41 a_15561_17999# tdc0.w_dly_sig\[23\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X42 a_7553_7663# a_7019_7669# a_7458_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X43 a_3686_18365# a_3413_17999# a_3601_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X44 _053_ a_10975_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X45 VGND _005_ a_12210_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X46 VGND tdc0.w_dly_sig\[28\] tdc0.w_dly_sig_n\[28\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X48 tdc0.w_dly_sig\[27\] tdc0.w_dly_sig_n\[26\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X51 a_6173_8207# a_6007_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X52 tdc0.w_dly_sig_n\[93\] tdc0.w_dly_sig\[93\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X53 a_8228_11305# a_7829_10933# a_8102_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X54 VPWR a_7074_15935# a_7001_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X55 a_11610_13380# a_11410_13225# a_11759_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X56 a_13947_5487# a_13165_5493# a_13863_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X57 tdc0.w_dly_sig\[76\] tdc0.w_dly_sig_n\[75\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X58 VPWR a_15887_15101# a_16055_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X59 _095_ a_14747_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X60 tdc0.w_dly_sig\[10\] tdc0.w_dly_sig\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X61 VPWR _002_ a_9319_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X62 a_10401_7369# _001_ a_10147_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X63 tdc0.w_dly_sig\[64\] tdc0.w_dly_sig_n\[63\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X64 a_10883_11721# _055_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X65 tdc0.w_dly_sig_n\[55\] tdc0.w_dly_sig\[55\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X66 tdc0.w_dly_sig\[122\] tdc0.w_dly_sig_n\[121\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X67 VPWR tdc0.w_dly_sig_n\[43\] tdc0.w_dly_sig\[44\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X68 a_4421_11305# a_3431_10933# a_4295_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X69 VPWR a_7856_14165# clknet_4_7_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X70 VPWR a_4755_4399# a_4923_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X71 a_16301_6031# _012_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X72 tdc0.w_dly_sig\[128\] tdc0.w_dly_sig_n\[127\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X73 a_12642_7271# net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X74 VGND tdc0.w_dly_sig\[24\] tdc0.w_dly_sig_n\[24\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X75 tdc0.w_dly_sig\[69\] tdc0.w_dly_sig_n\[68\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X76 a_12118_9295# _081_ a_12284_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X77 VGND tdc0.w_dly_sig\[96\] tdc0.w_dly_sig_n\[96\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X78 _026_ a_11490_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X79 tdc0.w_dly_sig\[11\] tdc0.w_dly_sig\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X80 a_2029_9295# a_1039_9295# a_1903_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X81 clknet_4_9_0_clk a_14664_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X82 a_10945_14735# a_10391_14709# a_10598_14709# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X83 a_10931_2919# a_11027_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X84 a_6177_12015# tdc0.w_dly_sig\[58\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X86 a_2858_17455# a_2585_17461# a_2773_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X88 a_4571_14013# a_3873_13647# a_4314_13759# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X89 tdc0.w_dly_sig\[15\] tdc0.w_dly_sig_n\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X90 _011_ a_13459_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X91 VPWR a_7286_7119# clknet_4_3_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X92 VPWR tdc0.w_dly_sig\[81\] tdc0.w_dly_sig\[83\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X93 a_16578_13103# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X95 a_17199_4917# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X96 a_17647_12247# a_17743_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X97 VPWR a_11122_7637# _029_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X98 VGND tdc0.w_dly_sig\[42\] tdc0.w_dly_sig_n\[42\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X99 VPWR tdc0.w_dly_sig\[12\] tdc0.w_dly_sig_n\[12\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X100 VGND a_4774_17429# a_4732_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X101 a_16915_10357# a_17206_10657# a_17157_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X102 a_13082_12292# a_12882_12137# a_13231_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X103 a_10598_14709# a_10391_14709# a_10774_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X104 a_17493_9295# tdc0.w_dly_sig\[120\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X105 VGND tdc0.o_result\[45\] a_10241_17775# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X106 tdc0.w_dly_sig\[116\] tdc0.w_dly_sig_n\[115\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X107 tdc0.w_dly_sig_n\[73\] tdc0.w_dly_sig_n\[71\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X108 VPWR a_5786_5055# a_5713_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X109 a_3509_5487# tdc0.w_dly_sig\[72\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X110 a_10873_16073# tdc0.o_result\[39\] a_10791_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X111 VPWR _086_ a_14944_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X112 a_13541_9071# tdc0.o_result\[84\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X113 VGND tdc0.w_dly_sig\[117\] a_18489_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X114 tdc0.w_dly_sig_n\[104\] tdc0.w_dly_sig_n\[102\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X115 VPWR tdc0.w_dly_sig\[25\] tdc0.w_dly_sig\[27\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X116 VPWR clknet_4_4_0_clk a_947_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X117 a_10527_14735# a_10391_14709# a_10107_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X118 VPWR a_16155_17687# _047_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X119 VPWR a_14783_2223# a_14951_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X120 a_14592_12809# _005_ a_14676_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X121 a_15198_13380# a_14991_13321# a_15374_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X122 a_16332_9839# _096_ a_16166_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X123 tdc0.o_result\[98\] a_13479_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X124 VPWR a_2363_10927# a_2531_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X125 tdc0.w_dly_sig\[4\] tdc0.w_dly_sig_n\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X126 VPWR a_14991_13321# a_14998_13225# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X127 tdc0.w_dly_sig_n\[49\] tdc0.w_dly_sig_n\[47\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X128 a_16248_9839# tdc0.o_result\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X129 VPWR tdc0.w_dly_sig\[44\] tdc0.w_dly_sig_n\[44\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X130 VGND a_12651_4123# a_12609_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X131 a_13990_8573# a_13551_8207# a_13905_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X132 tdc0.w_dly_sig_n\[1\] tdc0.w_dly_sig\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X133 a_10689_12809# _060_ a_10607_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X134 a_7274_6397# a_6835_6031# a_7189_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X135 a_12771_11159# a_12867_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X136 a_15127_13481# a_14991_13321# a_14707_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X137 VPWR net28 a_10321_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X138 tdc0.w_dly_sig_n\[23\] tdc0.w_dly_sig_n\[21\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X139 a_15220_8751# _018_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X140 VPWR a_14676_12809# uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X141 _010_ a_12134_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X142 a_14546_18365# a_14299_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X143 VGND tdc0.w_dly_sig_n\[15\] tdc0.w_dly_sig\[16\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X144 a_6633_15823# a_6467_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X145 tdc0.o_result\[53\] a_4279_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X146 a_2858_17455# a_2419_17461# a_2773_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X147 a_8481_8457# tdc0.o_result\[44\] a_8399_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X148 VPWR a_16331_1947# a_16247_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X149 VPWR _022_ a_7561_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X151 a_10931_2919# a_11027_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X152 a_16823_17973# a_17107_17973# a_17042_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X153 a_14729_15285# a_14563_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X154 net2 a_12999_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X155 a_8302_4765# a_7987_4631# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X156 VPWR a_12518_7119# _012_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X157 a_13705_11305# a_13151_11145# a_13358_11204# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X158 VGND a_18326_4676# a_18255_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X159 tdc0.o_result\[59\] a_7223_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X161 VGND clknet_0_clk a_14664_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X162 a_8941_6031# tdc0.o_result\[108\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X163 a_8565_15823# a_8399_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X165 a_13809_14197# a_13643_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X166 a_7783_6397# a_7001_6031# a_7699_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X167 a_11957_12393# a_11410_12137# a_11610_12292# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X169 a_18255_4777# a_18126_4521# a_17835_4631# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X171 tdc0.w_dly_sig\[35\] tdc0.w_dly_sig\[33\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X172 tdc0.o_result\[12\] a_14675_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X173 VPWR a_15162_5095# _086_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X174 a_14163_17973# clknet_4_13_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X175 tdc0.w_dly_sig\[114\] tdc0.w_dly_sig_n\[113\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X176 VGND tdc0.w_dly_sig\[102\] tdc0.w_dly_sig\[104\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X177 tdc0.w_dly_sig\[52\] tdc0.w_dly_sig\[50\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X178 VPWR tdc0.w_dly_sig_n\[119\] tdc0.w_dly_sig\[120\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X179 clknet_4_0_0_clk a_4176_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X180 a_9503_11043# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X181 VPWR a_11610_12292# a_11539_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X182 tdc0.w_dly_sig_n\[58\] tdc0.w_dly_sig_n\[56\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X183 VGND a_4923_1947# a_4881_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X185 _046_ a_11987_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X186 a_4237_17999# a_3247_17999# a_4111_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X188 VPWR net3 a_9779_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X189 tdc0.w_dly_sig_n\[123\] tdc0.w_dly_sig\[123\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X190 a_5169_9545# tdc0.o_result\[70\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X191 a_2087_9839# a_1223_9845# a_1830_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X192 VGND clknet_4_8_0_clk a_12447_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X193 tdc0.w_dly_sig_n\[99\] tdc0.w_dly_sig_n\[97\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X194 a_3593_12335# tdc0.o_result\[50\] a_3247_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X196 uo_out[5] a_11456_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 a_8872_17833# a_8473_17461# a_8746_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X198 tdc0.w_dly_sig\[99\] tdc0.w_dly_sig\[97\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X199 a_5713_5309# a_5179_4943# a_5618_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X200 a_2363_10927# a_1499_10933# a_2106_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X201 a_14121_18365# a_13783_18151# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X202 VGND a_11610_13380# a_11539_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X203 clknet_4_2_0_clk a_8500_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X204 VGND clknet_0_clk a_14388_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X205 _091_ a_6835_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X206 VGND tdc0.w_dly_sig\[124\] a_18121_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X207 a_9834_3285# a_9666_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X208 a_4314_5055# a_4146_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X209 VGND tdc0.w_dly_sig\[6\] tdc0.w_dly_sig_n\[6\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X210 VGND tdc0.w_dly_sig_n\[43\] tdc0.w_dly_sig_n\[45\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X211 a_17283_16599# a_17567_16585# a_17502_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X212 a_9319_12015# _013_ a_9401_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X213 tdc0.w_dly_sig_n\[0\] net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X214 VGND tdc0.w_dly_sig_n\[61\] tdc0.w_dly_sig_n\[63\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X215 tdc0.w_dly_sig_n\[23\] tdc0.w_dly_sig\[23\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X216 a_14358_2223# a_14085_2229# a_14273_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X217 a_6169_5807# tdc0.o_result\[83\] a_5823_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X218 VPWR a_7423_2223# a_7591_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X219 _033_ a_9595_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X220 a_5993_13647# tdc0.w_dly_sig\[37\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X221 a_7423_2223# a_6725_2229# a_7166_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X222 a_2033_10927# a_1499_10933# a_1938_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X223 a_13817_9295# tdc0.o_result\[60\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X224 a_4701_17455# a_4167_17461# a_4606_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X225 tdc0.w_dly_sig\[23\] tdc0.w_dly_sig_n\[22\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X226 VGND _000_ _019_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X227 a_4314_13759# a_4146_14013# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X228 VPWR clknet_4_13_0_clk a_14563_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X229 VPWR _037_ a_11685_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X230 tdc0.w_dly_sig\[33\] tdc0.w_dly_sig_n\[32\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X231 _037_ a_10239_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X232 a_3686_10749# a_3413_10383# a_3601_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X233 a_7139_10927# a_6357_10933# a_7055_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X234 a_11582_1791# a_11414_2045# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X236 a_12376_8751# _051_ a_12644_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X237 a_6906_16189# a_6467_15823# a_6821_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X238 VGND tdc0.w_dly_sig_n\[76\] tdc0.w_dly_sig\[77\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X239 a_14370_17973# a_14163_17973# a_14546_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X240 a_2125_3317# a_1959_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X241 clknet_4_10_0_clk a_16412_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X242 a_7198_17821# a_6883_17687# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X243 VPWR tdc0.w_dly_sig\[106\] tdc0.w_dly_sig_n\[106\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X244 a_7400_6031# a_7001_6031# a_7274_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X245 VGND tdc0.w_dly_sig_n\[95\] tdc0.w_dly_sig_n\[97\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X246 VGND tdc0.w_dly_sig_n\[98\] tdc0.w_dly_sig\[99\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X247 VGND tdc0.w_dly_sig\[63\] tdc0.w_dly_sig\[65\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X248 a_15465_10383# a_15299_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X249 a_9959_10633# _016_ a_9741_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X250 VGND tdc0.w_dly_sig\[16\] tdc0.w_dly_sig\[18\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X251 a_11473_4943# _001_ a_11359_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.137 ps=1.07 w=0.65 l=0.15
X252 VPWR clknet_4_1_0_clk a_1591_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X253 VPWR a_17567_17673# a_17574_17577# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X254 VPWR clknet_4_4_0_clk a_3431_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X255 VPWR _006_ a_14195_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X256 VPWR _015_ a_11609_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X257 VPWR tdc0.w_dly_sig_n\[91\] tdc0.w_dly_sig\[92\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X258 a_11057_17455# tdc0.o_result\[47\] a_10975_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X259 a_8201_12015# tdc0.w_dly_sig\[64\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X260 a_7286_7119# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X261 VPWR clknet_0_clk a_16412_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X262 a_17199_10357# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X263 VGND a_9747_8181# _007_ VGND sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.26 as=0.107 ps=0.98 w=0.65 l=0.15
X264 VPWR tdc0.w_dly_sig_n\[122\] tdc0.w_dly_sig_n\[124\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X265 a_3229_8757# a_3063_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X267 a_16155_14423# tdc0.o_result\[122\] a_16301_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X268 tdc0.w_dly_sig_n\[100\] tdc0.w_dly_sig_n\[98\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X269 VGND a_18027_3529# a_18034_3433# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X270 VGND clknet_4_1_0_clk a_4995_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X271 a_9493_12809# tdc0.o_result\[31\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X272 VPWR tdc0.w_dly_sig_n\[55\] tdc0.w_dly_sig\[56\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X273 VPWR clknet_4_5_0_clk a_3247_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X274 tdc0.w_dly_sig\[113\] tdc0.w_dly_sig_n\[112\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X275 a_14085_2229# a_13919_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X276 VPWR tdc0.w_dly_sig_n\[0\] tdc0.w_dly_sig\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X278 a_3698_12559# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X279 tdc0.w_dly_sig\[111\] tdc0.w_dly_sig\[109\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X280 VGND a_14675_14165# a_14633_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X281 VGND tdc0.w_dly_sig_n\[12\] tdc0.w_dly_sig\[13\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X282 VGND a_17774_2741# a_17703_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X283 a_7571_17161# _029_ a_7653_17161# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X284 VGND tdc0.w_dly_sig\[120\] tdc0.w_dly_sig\[122\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X285 a_7277_3311# a_6743_3317# a_7182_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X286 a_17555_10071# a_17651_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X287 VPWR tdc0.w_dly_sig_n\[24\] tdc0.w_dly_sig\[25\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X288 tdc0.w_dly_sig\[45\] tdc0.w_dly_sig_n\[44\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X289 tdc0.w_dly_sig\[48\] tdc0.w_dly_sig\[46\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X290 a_7423_2223# a_6559_2229# a_7166_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X291 a_16727_18151# a_16823_17973# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X293 a_9907_9661# a_9209_9295# a_9650_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X295 VPWR a_17314_17973# a_17243_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X296 a_11504_11445# _061_ a_11892_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X297 tdc0.o_result\[49\] a_3175_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X298 tdc0.w_dly_sig_n\[108\] tdc0.w_dly_sig\[108\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X299 tdc0.w_dly_sig\[127\] tdc0.w_dly_sig_n\[126\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X300 VPWR a_2106_10901# a_2033_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X302 a_14115_14735# a_13986_15009# a_13695_14709# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X303 VGND tdc0.w_dly_sig\[13\] tdc0.w_dly_sig_n\[13\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X304 a_9240_13481# a_8841_13109# a_9114_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X306 VPWR a_4774_17429# a_4701_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X309 a_16819_10535# a_16915_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X310 VPWR a_14031_5461# a_13947_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X311 VGND clknet_4_4_0_clk a_1131_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X312 tdc0.w_dly_sig_n\[29\] tdc0.w_dly_sig\[29\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X313 VGND tdc0.w_dly_sig\[73\] tdc0.w_dly_sig_n\[73\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X314 a_7090_9661# a_6817_9295# a_7005_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X315 VPWR tdc0.w_dly_sig\[52\] tdc0.w_dly_sig_n\[52\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X316 VGND _007_ a_10493_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X317 VPWR a_16332_9839# uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X318 VGND _010_ a_10401_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X319 a_3689_15285# a_3523_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X320 a_15035_9295# a_14899_9269# a_14615_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X321 a_15772_17999# a_15373_17999# a_15646_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X322 tdc0.w_dly_sig\[105\] tdc0.w_dly_sig_n\[104\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X323 a_14747_7663# _015_ a_14829_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X325 a_18291_6941# a_18071_6953# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X326 VPWR clknet_4_0_0_clk a_3891_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X327 a_6354_6575# a_6081_6581# a_6269_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X328 VPWR a_1903_11837# a_2071_11739# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X329 VGND tdc0.w_dly_sig_n\[37\] tdc0.w_dly_sig_n\[39\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X330 tdc0.w_dly_sig\[107\] tdc0.w_dly_sig_n\[106\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X331 VPWR a_16578_13103# clknet_4_15_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X332 VPWR a_4176_6005# clknet_4_0_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X333 VGND _080_ a_9366_10071# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X334 a_15807_12711# a_15903_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X336 VPWR tdc0.w_dly_sig_n\[111\] tdc0.w_dly_sig_n\[113\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X337 tdc0.o_result\[60\] a_7683_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X338 VPWR a_16394_12533# a_16323_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X339 VGND tdc0.w_dly_sig\[36\] tdc0.w_dly_sig_n\[36\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X340 a_14093_6281# _020_ a_13947_6183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X341 net8 a_12171_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X342 a_2398_3311# a_1959_3317# a_2313_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X343 VGND a_2290_1109# a_2248_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X344 VPWR clknet_4_11_0_clk a_16679_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X345 VPWR a_8500_4917# clknet_4_2_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X346 VPWR tdc0.w_dly_sig_n\[44\] tdc0.w_dly_sig\[45\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X347 tdc0.o_result\[101\] a_17527_1109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X348 VGND tdc0.w_dly_sig\[29\] tdc0.w_dly_sig\[31\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X349 VGND a_14491_1109# a_14449_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X350 VPWR tdc0.w_dly_sig\[78\] tdc0.w_dly_sig_n\[78\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X352 a_9661_7119# _003_ a_9589_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X353 VGND a_7883_7663# a_8051_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X354 a_14415_8573# a_13717_8207# a_14158_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X355 VGND a_12548_4917# clknet_4_8_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X356 tdc0.w_dly_sig_n\[38\] tdc0.w_dly_sig_n\[36\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X358 VPWR clknet_4_3_0_clk a_5915_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X359 a_12792_6549# _001_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.176 ps=1.68 w=0.42 l=0.15
X361 tdc0.o_result\[73\] a_2623_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X362 VGND a_13605_4917# _074_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X363 VPWR tdc0.w_dly_sig\[34\] tdc0.w_dly_sig_n\[34\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X364 a_10239_12015# _026_ a_10321_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X365 tdc0.w_dly_sig\[28\] tdc0.w_dly_sig\[26\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X366 a_9043_8751# _028_ a_9125_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X367 tdc0.w_dly_sig\[60\] tdc0.w_dly_sig_n\[59\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X368 VGND tdc0.w_dly_sig_n\[88\] tdc0.w_dly_sig_n\[90\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X369 VGND tdc0.w_dly_sig\[125\] a_17477_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X370 VPWR tdc0.w_dly_sig_n\[29\] tdc0.w_dly_sig\[30\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X371 tdc0.w_dly_sig_n\[48\] tdc0.w_dly_sig_n\[46\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X372 VGND a_15170_15253# a_15128_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X373 VPWR a_2255_9813# a_2171_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X374 VGND tdc0.w_dly_sig\[72\] tdc0.w_dly_sig\[74\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X375 VPWR tdc0.w_dly_sig\[26\] tdc0.w_dly_sig_n\[26\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X376 tdc0.w_dly_sig\[69\] tdc0.w_dly_sig\[67\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X377 _025_ a_9650_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X378 VGND a_16412_6549# clknet_4_10_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X379 clknet_4_7_0_clk a_7856_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X380 tdc0.w_dly_sig\[129\] tdc0.w_dly_sig_n\[128\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X381 VPWR net10 a_6181_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X383 a_9263_16189# a_8399_15823# a_9006_15935# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X384 VGND a_9006_15935# a_8964_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X385 VPWR a_14526_2197# a_14453_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X386 a_9839_4617# clknet_4_8_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X387 a_9459_4631# a_9555_4631# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X389 VPWR tdc0.w_dly_sig_n\[68\] tdc0.w_dly_sig\[69\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X390 a_6078_14013# a_5805_13647# a_5993_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X391 a_7829_10933# a_7663_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X392 a_7883_5487# a_7185_5493# a_7626_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X393 VGND a_15198_13380# a_15127_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X394 tdc0.o_result\[66\] a_5199_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X395 VGND a_6855_11989# a_6813_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X396 VGND tdc0.w_dly_sig\[58\] tdc0.w_dly_sig\[60\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X397 a_1577_14735# tdc0.w_dly_sig\[49\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X398 VGND tdc0.w_dly_sig\[79\] tdc0.w_dly_sig\[81\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X399 VGND tdc0.w_dly_sig\[110\] tdc0.w_dly_sig\[112\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X400 a_17283_2741# a_17567_2741# a_17502_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X401 tdc0.w_dly_sig_n\[92\] tdc0.w_dly_sig_n\[90\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X402 a_17187_17687# a_17283_17687# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X403 VPWR a_18171_9563# a_18087_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X404 _066_ a_15575_6281# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X405 _006_ a_11386_6652# a_11745_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.52 pd=3.04 as=0.135 ps=1.27 w=1 l=0.15
X406 _030_ a_8399_8457# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X407 a_14158_8319# a_13990_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X408 a_13753_9839# a_13415_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X409 VGND tdc0.w_dly_sig_n\[5\] tdc0.w_dly_sig\[6\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X410 a_7074_15935# a_6906_16189# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X411 a_9205_6031# tdc0.o_result\[68\] a_8859_6281# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X412 a_18291_10205# a_18071_10217# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X413 VPWR tdc0.w_dly_sig\[36\] tdc0.w_dly_sig\[38\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X414 net4 a_12631_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X415 a_7369_6397# a_6835_6031# a_7274_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X416 VGND a_3698_12559# clknet_4_4_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X417 tdc0.o_result\[64\] a_6027_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X418 a_2524_3689# a_2125_3317# a_2398_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X419 tdc0.w_dly_sig_n\[41\] tdc0.w_dly_sig_n\[39\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X420 tdc0.w_dly_sig_n\[5\] tdc0.w_dly_sig_n\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X421 VGND a_12318_7637# _015_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X423 a_3594_5487# a_3155_5493# a_3509_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X424 tdc0.w_dly_sig_n\[113\] tdc0.w_dly_sig\[113\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 VPWR tt_um_hpretl_tt06_tdc_22.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X425 VGND _052_ a_10883_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X426 a_5985_7119# a_4995_7119# a_5859_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X427 tdc0.w_dly_sig\[51\] tdc0.w_dly_sig\[49\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X428 a_9907_2045# a_9209_1679# a_9650_1791# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X429 tdc0.w_dly_sig\[54\] tdc0.w_dly_sig\[52\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X430 a_2271_6575# a_1573_6581# a_2014_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X431 VPWR tdc0.w_dly_sig\[125\] tdc0.w_dly_sig_n\[125\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X432 a_15327_13799# tdc0.o_result\[124\] a_15473_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X433 tdc0.w_dly_sig\[127\] tdc0.w_dly_sig\[125\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X434 VPWR clknet_4_9_0_clk a_12999_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X435 VGND tdc0.w_dly_sig\[30\] tdc0.w_dly_sig\[32\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X437 VGND tdc0.w_dly_sig\[120\] tdc0.w_dly_sig_n\[120\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X438 VPWR tdc0.w_dly_sig\[59\] tdc0.w_dly_sig\[61\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X439 tdc0.w_dly_sig_n\[99\] tdc0.w_dly_sig\[99\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X440 VGND tdc0.w_dly_sig_n\[34\] tdc0.w_dly_sig\[35\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X441 VGND a_13606_3285# a_13564_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X442 VGND a_11214_7093# _022_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X444 tdc0.w_dly_sig\[44\] tdc0.w_dly_sig_n\[43\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X445 a_10321_12015# tdc0.o_result\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X446 a_17950_14013# a_17703_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X447 VGND a_5694_14847# a_5652_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X449 a_18071_6953# a_17935_6793# a_17651_6807# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X450 a_14453_2223# a_13919_2229# a_14358_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X451 VGND clknet_4_0_0_clk a_5179_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X452 tdc0.w_dly_sig_n\[24\] tdc0.w_dly_sig\[24\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X453 VPWR a_7591_2197# a_7507_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X454 a_2581_4777# a_1591_4405# a_2455_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X455 VPWR a_7286_7119# clknet_4_3_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X456 tdc0.o_result\[60\] a_7683_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X457 a_9631_14191# a_8767_14197# a_9374_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X458 a_10321_10383# tdc0.o_result\[77\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X459 tdc0.w_dly_sig\[7\] tdc0.w_dly_sig_n\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X460 a_12875_12233# clknet_4_12_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X461 a_6826_17973# a_6626_18273# a_6975_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X462 tdc0.w_dly_sig_n\[117\] tdc0.w_dly_sig\[117\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X463 tdc0.w_dly_sig\[83\] tdc0.w_dly_sig_n\[82\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X464 VPWR _092_ a_16377_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X465 a_14829_7663# tdc0.o_result\[99\] a_14747_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X466 VPWR tdc0.w_dly_sig\[92\] tdc0.w_dly_sig_n\[92\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X467 VPWR a_9006_15935# a_8933_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X468 VPWR tdc0.w_dly_sig_n\[41\] tdc0.w_dly_sig_n\[43\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X469 VPWR tdc0.w_dly_sig\[71\] tdc0.w_dly_sig_n\[71\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X470 tdc0.w_dly_sig_n\[42\] tdc0.w_dly_sig\[42\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X471 VGND a_10259_3285# a_10217_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X474 a_13173_7779# _050_ a_13091_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X475 _021_ a_8859_6281# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X476 VGND a_12771_11159# tdc0.o_result\[5\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X477 a_4571_5309# a_3707_4943# a_4314_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X478 VGND a_2363_10927# a_2531_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X479 tdc0.w_dly_sig_n\[17\] tdc0.w_dly_sig\[17\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X480 VGND tdc0.w_dly_sig_n\[108\] tdc0.w_dly_sig\[109\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X481 VPWR tdc0.w_dly_sig\[107\] tdc0.w_dly_sig\[109\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X482 VPWR clknet_4_10_0_clk a_16495_1141# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X483 a_10585_9071# tdc0.o_result\[30\] a_10239_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X484 net11 a_14195_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X485 VGND _005_ a_14786_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X486 VPWR a_1979_11989# a_1895_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X487 VGND _002_ _019_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X488 tdc0.w_dly_sig_n\[114\] tdc0.w_dly_sig_n\[112\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X489 a_14676_12809# _005_ a_14592_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X490 tdc0.w_dly_sig\[77\] tdc0.w_dly_sig_n\[76\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X491 a_6813_7119# tdc0.o_result\[80\] a_6467_7369# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X492 VGND tdc0.w_dly_sig_n\[82\] tdc0.w_dly_sig_n\[84\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X493 VGND tdc0.w_dly_sig\[87\] tdc0.w_dly_sig_n\[87\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X494 tdc0.w_dly_sig_n\[50\] tdc0.w_dly_sig\[50\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X495 _013_ a_11159_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.213 ps=1.3 w=0.65 l=0.15
X496 a_6127_5309# a_5345_4943# a_6043_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X497 VPWR a_6522_6549# a_6449_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X498 a_4774_6549# a_4606_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X499 clknet_4_6_0_clk a_6550_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X500 VPWR a_17719_8359# _052_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X501 a_14081_9295# tdc0.o_result\[28\] a_13735_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X503 a_11119_12247# a_11403_12233# a_11338_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X504 VPWR tdc0.w_dly_sig_n\[63\] tdc0.w_dly_sig\[64\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X505 VPWR tdc0.w_dly_sig_n\[31\] tdc0.w_dly_sig\[32\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X506 a_15098_16189# a_14851_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X507 VPWR tdc0.w_dly_sig\[115\] a_18673_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X508 _006_ _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X509 VPWR tdc0.w_dly_sig_n\[51\] tdc0.w_dly_sig_n\[53\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X510 a_3854_10495# a_3686_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X511 a_1846_6575# a_1573_6581# a_1761_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X512 tdc0.o_result\[59\] a_7223_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X513 a_13905_8207# tdc0.w_dly_sig\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X514 _075_ a_11251_8457# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X515 VPWR clknet_4_7_0_clk a_6467_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X516 a_2547_5309# a_1849_4943# a_2290_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X517 a_3720_5865# a_3321_5493# a_3594_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X518 a_9501_9955# _077_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X520 a_17774_17732# a_17567_17673# a_17950_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X521 a_13599_4007# a_13695_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X522 tdc0.w_dly_sig_n\[85\] tdc0.w_dly_sig_n\[83\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X523 a_15393_5193# _083_ a_15297_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
R1 uio_out[2] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X524 VGND tdc0.w_dly_sig_n\[61\] tdc0.w_dly_sig\[62\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X525 a_8987_16367# a_8123_16373# a_8730_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X526 VPWR tdc0.w_dly_sig\[106\] tdc0.w_dly_sig\[108\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X527 a_9389_1513# a_8399_1141# a_9263_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X528 VGND a_4130_15253# a_4088_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X529 a_17635_2045# a_16771_1679# a_17378_1791# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X530 tdc0.w_dly_sig_n\[71\] tdc0.w_dly_sig_n\[69\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X531 a_17627_8751# a_16845_8757# a_17543_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X532 _058_ a_9411_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X533 VPWR ui_in[0] a_18187_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X534 VPWR a_10075_1947# a_9991_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X535 a_2037_1135# tdc0.w_dly_sig\[83\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X536 VGND tdc0.o_result\[117\] a_18613_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X537 a_12591_12247# a_12882_12137# a_12833_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X538 tdc0.w_dly_sig\[12\] tdc0.w_dly_sig_n\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X539 a_9393_3317# a_9227_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X540 a_5985_6031# tdc0.o_result\[82\] a_5639_6281# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X541 a_7001_6031# a_6835_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X542 a_11333_8207# tdc0.o_result\[73\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X543 tdc0.w_dly_sig_n\[51\] tdc0.w_dly_sig\[51\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X544 a_8657_16367# a_8123_16373# a_8562_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X546 tdc0.w_dly_sig_n\[119\] tdc0.w_dly_sig\[119\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X548 a_4176_6005# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X549 tdc0.w_dly_sig_n\[61\] tdc0.w_dly_sig\[61\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X550 a_3601_14735# tdc0.w_dly_sig\[47\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X551 tdc0.w_dly_sig_n\[56\] tdc0.w_dly_sig_n\[54\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X552 a_4314_5055# a_4146_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X553 tdc0.w_dly_sig_n\[62\] tdc0.w_dly_sig_n\[60\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X554 VPWR tdc0.o_result\[0\] a_16248_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X555 a_11372_10927# tdc0.o_result\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X556 VPWR tdc0.w_dly_sig_n\[67\] tdc0.w_dly_sig\[68\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 _054_ a_10226_11247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X558 VPWR a_6430_11989# a_6357_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X559 VGND _025_ a_17036_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X561 tdc0.w_dly_sig\[120\] tdc0.w_dly_sig_n\[119\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X562 tdc0.o_result\[87\] a_6395_1947# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X563 a_6273_17775# tdc0.o_result\[42\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X564 VGND tdc0.w_dly_sig_n\[107\] tdc0.w_dly_sig\[108\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X565 VGND a_18179_8983# _039_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X566 VGND tdc0.w_dly_sig\[54\] tdc0.w_dly_sig_n\[54\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X567 VGND a_3790_7119# clknet_4_1_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X568 a_5602_7231# a_5434_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X569 tdc0.w_dly_sig_n\[75\] tdc0.w_dly_sig\[75\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X570 a_15553_4777# a_14563_4405# a_15427_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X571 tdc0.w_dly_sig\[115\] tdc0.w_dly_sig\[113\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X572 a_7653_16911# tdc0.o_result\[40\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X573 VGND clknet_4_0_0_clk a_1683_1141# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X574 VPWR _000_ a_10975_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X575 VPWR a_11456_10927# uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X576 tdc0.o_result\[100\] a_14031_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X577 a_17567_16585# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X578 VGND tdc0.w_dly_sig\[85\] tdc0.w_dly_sig_n\[85\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X579 _071_ a_7755_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X580 VPWR tdc0.w_dly_sig_n\[28\] tdc0.w_dly_sig\[29\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X581 VPWR tdc0.w_dly_sig\[22\] tdc0.w_dly_sig\[24\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X582 tdc0.w_dly_sig_n\[45\] tdc0.w_dly_sig_n\[43\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X583 tdc0.w_dly_sig_n\[6\] tdc0.w_dly_sig\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X584 tdc0.w_dly_sig_n\[96\] tdc0.w_dly_sig\[96\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X585 VPWR a_4019_5487# a_4187_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X586 VPWR tdc0.o_result\[5\] a_11372_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X587 a_11246_2767# a_10931_2919# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X588 VPWR a_8543_7093# _020_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.143 pd=1.33 as=0.153 ps=1.3 w=1 l=0.15
X589 a_13599_4007# a_13695_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X590 tdc0.w_dly_sig_n\[126\] tdc0.w_dly_sig_n\[124\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X591 tdc0.w_dly_sig\[88\] tdc0.w_dly_sig_n\[87\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X592 VPWR tdc0.w_dly_sig_n\[96\] tdc0.w_dly_sig\[97\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X593 _067_ a_6467_7369# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X594 VPWR tdc0.w_dly_sig_n\[1\] tdc0.w_dly_sig_n\[3\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X595 a_13931_10217# a_13795_10057# a_13511_10071# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X597 VPWR clknet_4_11_0_clk a_17139_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X598 VGND a_17935_6793# a_17942_6697# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X599 a_16122_12559# a_15807_12711# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X600 a_8491_5487# _028_ a_8573_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X601 VGND _062_ a_15575_6281# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X602 VPWR a_12495_12247# tdc0.o_result\[7\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X603 a_6099_16367# _029_ a_6181_16687# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X604 VPWR tdc0.w_dly_sig\[62\] tdc0.w_dly_sig\[64\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X605 tdc0.w_dly_sig\[21\] tdc0.w_dly_sig\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X606 a_7699_4221# a_7001_3855# a_7442_3967# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X607 tdc0.w_dly_sig_n\[14\] tdc0.w_dly_sig\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X608 VGND tdc0.o_result\[6\] a_12210_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X609 VGND tdc0.w_dly_sig_n\[102\] tdc0.w_dly_sig\[103\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X611 clknet_4_12_0_clk a_12548_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X612 VGND a_8270_10901# a_8228_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X613 VPWR a_9366_10071# _081_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X614 tdc0.w_dly_sig\[109\] tdc0.w_dly_sig\[107\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X615 VPWR clknet_4_3_0_clk a_7571_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X616 a_15170_15253# a_15002_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X617 VGND a_7626_7637# a_7584_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X618 VGND _027_ a_9043_8457# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X619 VGND net5 a_14287_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X620 VPWR a_16762_8207# clknet_4_11_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X621 tdc0.w_dly_sig_n\[57\] tdc0.w_dly_sig\[57\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X622 VGND a_17567_2741# a_17574_3041# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X623 VGND a_12483_4221# a_12651_4123# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X625 VGND tdc0.w_dly_sig_n\[123\] tdc0.w_dly_sig_n\[125\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X626 a_4057_4405# a_3891_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X627 clknet_0_clk a_11058_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X628 VPWR tdc0.w_dly_sig\[103\] tdc0.w_dly_sig\[105\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X629 tdc0.o_result\[53\] a_4279_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X631 a_4038_10901# a_3870_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X632 a_8481_6895# tdc0.o_result\[91\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X633 VPWR tdc0.w_dly_sig_n\[4\] tdc0.w_dly_sig\[5\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X634 _077_ a_4535_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X635 a_13735_9545# _013_ a_13817_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X636 tdc0.w_dly_sig\[97\] tdc0.w_dly_sig_n\[96\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X638 tdc0.w_dly_sig_n\[102\] tdc0.w_dly_sig\[102\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X639 tdc0.w_dly_sig\[66\] tdc0.w_dly_sig\[64\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X641 tdc0.w_dly_sig_n\[50\] tdc0.w_dly_sig_n\[48\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X642 tdc0.w_dly_sig\[56\] tdc0.w_dly_sig\[54\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X643 a_9666_3311# a_9227_3317# a_9581_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X645 tdc0.w_dly_sig\[122\] tdc0.w_dly_sig\[120\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X646 VPWR a_17774_13621# a_17703_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
R2 tt_um_hpretl_tt06_tdc_12.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X647 tdc0.w_dly_sig_n\[2\] tdc0.w_dly_sig_n\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X648 a_13353_3311# tdc0.w_dly_sig\[101\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X649 VPWR a_17102_1109# a_17029_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X650 a_5433_9295# tdc0.o_result\[70\] a_5087_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X651 _012_ a_12518_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X652 a_17555_10071# a_17651_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X653 VGND tdc0.w_dly_sig\[21\] tdc0.w_dly_sig\[23\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X654 VPWR tdc0.w_dly_sig\[15\] tdc0.w_dly_sig_n\[15\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X655 a_14633_14569# a_13643_14197# a_14507_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X656 VGND tdc0.w_dly_sig_n\[90\] tdc0.w_dly_sig\[91\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X657 a_1393_9295# tdc0.w_dly_sig\[76\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X658 a_11892_11471# _061_ a_11504_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X659 VGND clknet_4_4_0_clk a_4259_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X660 VGND a_3007_14191# a_3175_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X661 VGND tdc0.w_dly_sig\[124\] tdc0.w_dly_sig\[126\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X662 a_14633_6953# a_13643_6581# a_14507_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X663 VPWR net3 a_12171_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X664 tdc0.w_dly_sig_n\[13\] tdc0.w_dly_sig\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X665 VGND tdc0.w_dly_sig_n\[78\] tdc0.w_dly_sig\[79\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X666 VPWR tdc0.w_dly_sig\[14\] a_11957_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X667 VPWR tdc0.w_dly_sig_n\[12\] tdc0.w_dly_sig_n\[14\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X668 a_10423_5193# _020_ a_10505_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X669 a_17778_14557# a_17463_14423# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X670 VGND a_9171_17455# a_9339_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X671 tdc0.w_dly_sig_n\[26\] tdc0.w_dly_sig\[26\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X672 clknet_4_3_0_clk a_7286_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X673 a_8611_10927# a_7829_10933# a_8527_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
R3 VGND uio_out[6] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X674 VPWR a_8995_7093# a_8543_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X675 a_18325_8751# _025_ a_18179_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X676 VPWR tdc0.w_dly_sig\[126\] a_18121_16745# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X677 a_2547_1135# a_1683_1141# a_2290_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X678 a_15427_15279# a_14729_15285# a_15170_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X679 VGND tdc0.w_dly_sig\[88\] tdc0.w_dly_sig\[90\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X680 VGND tdc0.w_dly_sig\[65\] tdc0.w_dly_sig\[67\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X681 a_17935_10057# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X682 VGND a_4866_13077# a_4824_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X683 a_6154_17023# a_5986_17277# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X684 tdc0.w_dly_sig\[58\] tdc0.w_dly_sig_n\[57\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X685 tdc0.w_dly_sig_n\[52\] tdc0.w_dly_sig\[52\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X686 VPWR tdc0.w_dly_sig\[114\] tdc0.w_dly_sig\[116\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X687 VPWR tdc0.w_dly_sig\[55\] tdc0.w_dly_sig_n\[55\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X688 VPWR tdc0.w_dly_sig_n\[121\] tdc0.w_dly_sig\[122\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X689 _010_ a_12134_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X690 VPWR a_2163_13077# a_2079_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X691 VPWR a_16578_13103# clknet_4_15_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X692 a_18489_10217# a_17935_10057# a_18142_10116# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X693 a_12376_8751# _046_ a_12210_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X694 a_18071_10217# a_17942_9961# a_17651_10071# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X695 VPWR a_15327_13799# _008_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X696 a_6181_16367# tdc0.o_result\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X697 a_7181_11305# a_6191_10933# a_7055_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X698 a_9482_9661# a_9043_9295# a_9397_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X699 a_4881_9071# tdc0.o_result\[81\] a_4535_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X700 VPWR tdc0.w_dly_sig\[15\] tdc0.w_dly_sig\[17\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X701 a_10229_16073# tdc0.o_result\[125\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X703 a_10791_16073# net6 a_10873_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X704 a_4866_13077# a_4698_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X705 VPWR net4 a_11159_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.22 ps=1.44 w=1 l=0.15
X707 tdc0.w_dly_sig_n\[36\] tdc0.w_dly_sig\[36\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X708 tdc0.w_dly_sig_n\[77\] tdc0.w_dly_sig\[77\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X709 a_1301_12015# tdc0.w_dly_sig\[75\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X710 clknet_4_4_0_clk a_3698_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X712 a_14066_1109# a_13898_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X713 a_1662_9839# a_1223_9845# a_1577_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X714 tdc0.w_dly_sig\[14\] tdc0.w_dly_sig_n\[13\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X715 VPWR a_17803_1947# a_17719_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X717 a_9171_17455# a_8307_17461# a_8914_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X718 a_4698_13103# a_4425_13109# a_4613_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X719 VPWR tdc0.w_dly_sig_n\[109\] tdc0.w_dly_sig\[110\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X720 VGND tdc0.w_dly_sig\[98\] tdc0.w_dly_sig\[100\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X721 VPWR a_17567_2741# a_17574_3041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X722 a_9774_4765# a_9459_4631# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X723 VGND tdc0.w_dly_sig_n\[117\] tdc0.w_dly_sig\[118\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X724 _072_ a_11251_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X725 VGND tdc0.w_dly_sig\[45\] tdc0.w_dly_sig\[47\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X726 tdc0.w_dly_sig\[75\] tdc0.w_dly_sig_n\[74\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X727 VPWR clknet_4_0_0_clk a_3707_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X729 VPWR tdc0.w_dly_sig\[56\] tdc0.w_dly_sig\[58\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X730 a_12810_7119# net3 a_12696_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.137 ps=1.07 w=0.65 l=0.15
X731 VPWR tdc0.w_dly_sig\[122\] a_18489_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X732 a_9792_3689# a_9393_3317# a_9666_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
R4 VGND uio_oe[0] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X734 tdc0.w_dly_sig_n\[87\] tdc0.w_dly_sig_n\[85\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X735 VPWR _012_ a_16117_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X736 tdc0.o_result\[91\] a_7959_1109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X738 VGND tdc0.w_dly_sig_n\[31\] tdc0.w_dly_sig_n\[33\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X740 tdc0.o_result\[42\] a_5199_17429# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X741 VGND a_13863_5487# a_14031_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X742 a_2949_12335# tdc0.o_result\[48\] a_2603_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X743 a_2198_17023# a_2030_17277# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X744 tdc0.w_dly_sig_n\[81\] tdc0.w_dly_sig_n\[79\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X745 tdc0.w_dly_sig\[115\] tdc0.w_dly_sig_n\[114\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X746 VGND a_12171_5487# net8 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X747 _088_ a_6191_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X748 VGND a_14783_2223# a_14951_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X749 a_17835_7895# a_18126_7785# a_18077_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X750 a_5997_13103# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X752 VPWR tdc0.w_dly_sig\[115\] tdc0.w_dly_sig_n\[115\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X753 VGND a_5583_18365# a_5751_18267# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X754 tdc0.o_result\[42\] a_5199_17429# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X755 VGND a_12284_9545# uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X756 tdc0.w_dly_sig_n\[64\] tdc0.w_dly_sig_n\[62\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X757 clknet_4_15_0_clk a_16578_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X758 a_17187_13799# a_17283_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X759 VPWR a_14952_8751# uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X760 tdc0.o_result\[40\] a_6579_17179# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X762 VPWR a_8500_4917# clknet_4_2_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X763 tdc0.w_dly_sig_n\[12\] tdc0.w_dly_sig\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X764 tdc0.w_dly_sig\[36\] tdc0.w_dly_sig_n\[35\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X765 VPWR tdc0.w_dly_sig_n\[48\] tdc0.w_dly_sig\[49\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X766 clknet_4_11_0_clk a_16762_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X767 _062_ a_8491_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X768 tdc0.w_dly_sig\[92\] tdc0.w_dly_sig_n\[91\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X769 a_10977_4399# tdc0.o_result\[86\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X770 VGND tdc0.w_dly_sig_n\[112\] tdc0.w_dly_sig\[113\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X771 a_5786_5055# a_5618_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X772 tdc0.w_dly_sig\[73\] tdc0.w_dly_sig\[71\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X773 tdc0.o_result\[30\] a_10075_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X774 a_9121_3855# tdc0.w_dly_sig\[110\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X775 VGND a_17187_17687# tdc0.o_result\[127\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X777 VGND tdc0.w_dly_sig_n\[120\] tdc0.w_dly_sig\[121\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X778 a_15373_17999# a_15207_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X779 a_3601_17999# tdc0.w_dly_sig\[44\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X780 tdc0.w_dly_sig_n\[43\] tdc0.w_dly_sig_n\[41\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X781 a_1941_6575# a_1407_6581# a_1846_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X782 VPWR tdc0.w_dly_sig_n\[63\] tdc0.w_dly_sig_n\[65\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X783 a_16166_10159# tdc0.o_result\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X784 VPWR tdc0.w_dly_sig\[43\] tdc0.w_dly_sig\[45\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X785 a_11403_13321# clknet_4_12_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X786 VGND tdc0.w_dly_sig\[18\] tdc0.w_dly_sig_n\[18\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X788 tdc0.w_dly_sig\[6\] tdc0.w_dly_sig_n\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X789 VGND tdc0.w_dly_sig\[61\] tdc0.w_dly_sig\[63\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X790 VPWR a_9531_5095# _035_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X791 a_9493_12559# tdc0.o_result\[63\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X792 a_11023_13335# a_11119_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X793 net9 a_9227_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X794 VGND tdc0.w_dly_sig_n\[59\] tdc0.w_dly_sig_n\[61\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X795 a_8573_5807# tdc0.o_result\[88\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X796 a_7001_16189# a_6467_15823# a_6906_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X797 tdc0.w_dly_sig_n\[110\] tdc0.w_dly_sig_n\[108\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X798 a_9493_2543# tdc0.o_result\[93\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X799 a_9608_9295# a_9209_9295# a_9482_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X800 a_6081_6581# a_5915_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X801 a_11839_2045# a_10975_1679# a_11582_1791# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X802 tdc0.w_dly_sig_n\[73\] tdc0.w_dly_sig\[73\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X803 VGND tdc0.w_dly_sig_n\[25\] tdc0.w_dly_sig\[26\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X804 VGND a_16412_6549# clknet_4_10_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X805 a_9959_10633# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X806 VPWR clknet_0_clk a_6550_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X807 a_5345_4943# a_5179_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X808 a_5115_17455# a_4333_17461# a_5031_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X810 a_8519_8751# a_7737_8757# a_8435_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X811 a_7458_5487# a_7019_5493# a_7373_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X812 _065_ a_14563_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X814 _048_ a_5087_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X815 a_2773_17455# tdc0.w_dly_sig\[46\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X816 a_8921_4777# a_8374_4521# a_8574_4676# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X817 VGND tdc0.w_dly_sig_n\[94\] tdc0.w_dly_sig_n\[96\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X818 VPWR clknet_0_clk a_7286_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X819 a_7373_7663# tdc0.w_dly_sig\[36\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X822 VGND tdc0.w_dly_sig_n\[67\] tdc0.w_dly_sig_n\[69\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X823 tdc0.w_dly_sig\[32\] tdc0.w_dly_sig\[30\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X824 tdc0.w_dly_sig_n\[103\] tdc0.w_dly_sig\[103\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X825 a_6549_7119# tdc0.o_result\[64\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X826 VGND a_7423_2223# a_7591_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X828 VGND a_16732_11445# _356_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X829 _025_ a_9650_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X830 tdc0.o_result\[70\] a_4095_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X831 VGND _001_ a_9761_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=1 as=0.0619 ps=0.715 w=0.42 l=0.15
X832 a_16727_18151# a_16823_17973# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X833 VPWR tdc0.w_dly_sig_n\[53\] tdc0.w_dly_sig_n\[55\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X834 tdc0.o_result\[36\] a_6671_13915# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X835 a_11027_2741# a_11311_2741# a_11246_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
R5 VPWR tt_um_hpretl_tt06_tdc_18.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X836 clknet_4_14_0_clk a_17314_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X837 VPWR a_12875_12233# a_12882_12137# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X838 a_4111_15101# a_3413_14735# a_3854_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X840 a_15377_14735# tdc0.w_dly_sig\[28\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X841 _044_ a_11146_4719# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X842 a_15002_4399# a_14729_4405# a_14917_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X843 tdc0.w_dly_sig\[85\] tdc0.w_dly_sig\[83\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X844 a_4245_1679# tdc0.w_dly_sig\[86\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X845 a_12297_8457# _003_ a_12201_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X846 a_6554_17999# a_6239_18151# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X847 VPWR a_12483_4221# a_12651_4123# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X848 VPWR a_12642_7271# a_12518_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X849 a_9029_13103# tdc0.w_dly_sig\[32\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X850 a_14362_15101# a_14115_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
R6 tt_um_hpretl_tt06_tdc_25.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X851 VPWR clknet_4_4_0_clk a_6191_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X852 VPWR a_2715_1109# a_2631_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X853 a_15002_15279# a_14563_15285# a_14917_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X854 VPWR tdc0.w_dly_sig_n\[110\] tdc0.w_dly_sig\[111\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X855 a_9482_2045# a_9043_1679# a_9397_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X856 a_9631_14191# a_8933_14197# a_9374_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X858 tdc0.w_dly_sig\[68\] tdc0.w_dly_sig\[66\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X862 VPWR a_16181_5461# _084_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X863 tdc0.w_dly_sig\[41\] tdc0.w_dly_sig_n\[40\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X864 VPWR a_9741_10357# _034_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X865 a_5951_15101# a_5087_14735# a_5694_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X866 a_6246_13759# a_6078_14013# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X867 VPWR tdc0.w_dly_sig_n\[28\] tdc0.w_dly_sig_n\[30\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X868 a_5349_7119# tdc0.w_dly_sig\[65\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X869 a_17283_13621# a_17567_13621# a_17502_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X870 VPWR net2 a_11386_6652# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X871 VGND a_2163_13077# a_2121_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X872 a_1662_15101# a_1223_14735# a_1577_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X873 clknet_4_6_0_clk a_6550_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X874 VGND a_14664_6005# clknet_4_9_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X875 a_16127_7779# _095_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X876 tdc0.w_dly_sig_n\[114\] tdc0.w_dly_sig\[114\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X877 _003_ a_14287_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X878 a_3247_12015# _026_ a_3329_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X879 VGND tdc0.w_dly_sig_n\[91\] tdc0.w_dly_sig_n\[93\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X880 tdc0.w_dly_sig\[116\] tdc0.w_dly_sig\[114\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X881 VPWR a_18187_10901# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X882 a_11403_12233# clknet_4_12_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X883 VPWR tdc0.w_dly_sig\[69\] tdc0.w_dly_sig_n\[69\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X884 tdc0.w_dly_sig\[4\] tdc0.w_dly_sig\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X886 tdc0.w_dly_sig\[81\] tdc0.w_dly_sig\[79\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X887 VGND a_9650_9407# a_9608_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X888 a_18234_3588# a_18034_3433# a_18383_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X889 VPWR tdc0.w_dly_sig\[46\] tdc0.w_dly_sig\[48\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X890 a_4521_6575# tdc0.w_dly_sig\[67\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X891 VGND tdc0.w_dly_sig_n\[103\] tdc0.w_dly_sig\[104\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X892 VPWR a_13479_2197# a_13395_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X893 tdc0.w_dly_sig_n\[105\] tdc0.w_dly_sig_n\[103\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X894 tdc0.w_dly_sig\[117\] tdc0.w_dly_sig_n\[116\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X895 a_14944_12809# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X896 VPWR tdc0.w_dly_sig_n\[34\] tdc0.w_dly_sig_n\[36\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X897 tdc0.w_dly_sig\[59\] tdc0.w_dly_sig\[57\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X898 a_15198_13380# a_14998_13225# a_15347_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X899 tdc0.w_dly_sig_n\[53\] tdc0.w_dly_sig_n\[51\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X900 VPWR _000_ a_11159_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.135 ps=1.27 w=1 l=0.15
X901 a_10785_12809# _059_ a_10689_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X902 VGND a_14066_1109# a_14024_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X903 VPWR a_12548_14165# clknet_4_12_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X904 VPWR _021_ a_9293_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X905 a_7584_5865# a_7185_5493# a_7458_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X906 _016_ _000_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X907 a_16301_14511# _007_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X908 _101_ a_6467_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X910 tdc0.w_dly_sig_n\[98\] tdc0.w_dly_sig_n\[96\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X911 tdc0.w_dly_sig\[62\] tdc0.w_dly_sig_n\[61\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X912 a_7032_15823# a_6633_15823# a_6906_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X913 a_16187_12533# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X914 a_4697_13647# a_3707_13647# a_4571_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X915 clknet_4_2_0_clk a_8500_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X917 VPWR tdc0.w_dly_sig_n\[72\] tdc0.w_dly_sig_n\[74\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X918 VGND tdc0.w_dly_sig\[5\] tdc0.w_dly_sig_n\[5\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X919 a_2037_4943# tdc0.w_dly_sig\[80\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X920 a_18187_10901# ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X921 a_14533_14735# a_13979_14709# a_14186_14709# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X922 tdc0.w_dly_sig_n\[91\] tdc0.w_dly_sig_n\[89\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X923 clknet_4_4_0_clk a_3698_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X924 a_8764_7119# _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.104 ps=1 w=0.42 l=0.15
X925 a_3689_5487# a_3155_5493# a_3594_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X926 VPWR clknet_4_9_0_clk a_13551_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X927 a_15575_6281# _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X928 a_9043_6575# _026_ a_9125_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X929 VGND a_7856_14165# clknet_4_7_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X931 VGND tdc0.w_dly_sig\[70\] tdc0.w_dly_sig_n\[70\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X932 a_16248_12015# _005_ a_16332_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X933 VGND tdc0.w_dly_sig\[3\] tdc0.w_dly_sig\[5\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X934 VGND a_12007_1947# a_11965_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X935 a_14115_3855# a_13979_3829# a_13695_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X936 tdc0.o_result\[95\] a_10075_1947# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X937 VGND a_11058_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X938 VPWR a_6395_12827# a_6311_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X939 a_17283_13621# a_17574_13921# a_17525_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X941 VGND tdc0.w_dly_sig\[34\] tdc0.w_dly_sig\[36\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X942 VGND _034_ a_9503_11043# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X943 a_11759_13469# a_11539_13481# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X944 a_14186_14709# a_13979_14709# a_14362_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X945 VGND tdc0.w_dly_sig_n\[17\] tdc0.w_dly_sig\[18\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X946 tdc0.w_dly_sig_n\[54\] tdc0.w_dly_sig\[54\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X947 a_3601_10383# tdc0.w_dly_sig\[54\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X948 tdc0.w_dly_sig_n\[75\] tdc0.w_dly_sig_n\[73\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X949 VGND a_6550_13103# clknet_4_6_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X950 a_13606_3285# a_13438_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X951 VPWR tdc0.w_dly_sig_n\[10\] tdc0.w_dly_sig_n\[12\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X952 VPWR tdc0.w_dly_sig_n\[57\] tdc0.w_dly_sig_n\[59\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X953 a_17406_4917# a_17199_4917# a_17582_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X954 a_2122_5309# a_1683_4943# a_2037_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X955 clknet_4_10_0_clk a_16412_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X956 a_13898_1135# a_13459_1141# a_13813_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X957 a_5441_3855# tdc0.w_dly_sig\[87\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X958 tdc0.w_dly_sig\[37\] tdc0.w_dly_sig\[35\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X959 a_14115_14735# a_13979_14709# a_13695_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X960 tdc0.w_dly_sig\[29\] tdc0.w_dly_sig_n\[28\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X961 VPWR a_17107_17973# a_17114_18273# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X962 a_9608_1679# a_9209_1679# a_9482_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X963 tdc0.w_dly_sig_n\[15\] tdc0.w_dly_sig\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X964 VGND tdc0.w_dly_sig_n\[20\] tdc0.w_dly_sig_n\[22\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X965 VGND tdc0.w_dly_sig_n\[71\] tdc0.w_dly_sig\[72\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X966 VPWR a_2823_3311# a_2991_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X967 a_17651_6807# a_17942_6697# a_17893_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X969 a_17923_17821# a_17703_17833# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X970 a_10493_15823# tdc0.o_result\[125\] a_10147_16073# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X971 VPWR clknet_4_6_0_clk a_5639_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X973 VPWR ui_in[6] a_11711_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X974 tdc0.w_dly_sig_n\[3\] tdc0.w_dly_sig_n\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X976 a_10595_7369# _003_ _016_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X977 tdc0.o_result\[101\] a_17527_1109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X978 VGND a_4176_6005# clknet_4_0_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X979 a_13429_12393# a_12875_12233# a_13082_12292# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X980 VGND _057_ a_10607_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X981 tdc0.o_result\[61\] a_8695_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X982 VPWR tdc0.w_dly_sig\[1\] tdc0.w_dly_sig\[3\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X983 VGND tdc0.w_dly_sig_n\[45\] tdc0.w_dly_sig\[46\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X984 VPWR tdc0.w_dly_sig_n\[36\] tdc0.w_dly_sig\[37\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X985 a_11724_10927# _041_ a_11456_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X986 a_14066_1109# a_13898_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X987 a_2121_13481# a_1131_13109# a_1995_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X988 VPWR tdc0.w_dly_sig\[26\] a_15269_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X989 a_18581_3689# a_18027_3529# a_18234_3588# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X990 VPWR a_3927_8751# a_4095_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X991 tdc0.w_dly_sig\[64\] tdc0.w_dly_sig\[62\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X992 a_1738_13077# a_1570_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X995 a_2907_3311# a_2125_3317# a_2823_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X996 VGND _072_ a_11619_8867# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X997 a_12200_9545# tdc0.o_result\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X998 VGND tdc0.w_dly_sig\[82\] tdc0.w_dly_sig_n\[82\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X999 a_18119_7881# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1000 tdc0.w_dly_sig_n\[56\] tdc0.w_dly_sig\[56\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1001 a_15269_15823# a_14715_15797# a_14922_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1002 VGND clknet_4_3_0_clk a_7019_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1003 tdc0.w_dly_sig\[109\] tdc0.w_dly_sig_n\[108\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1004 tdc0.w_dly_sig\[55\] tdc0.w_dly_sig\[53\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1006 a_1573_6581# a_1407_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1007 VPWR tdc0.w_dly_sig_n\[53\] tdc0.w_dly_sig\[54\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1008 clknet_4_5_0_clk a_3348_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1009 VPWR tdc0.w_dly_sig_n\[120\] tdc0.w_dly_sig_n\[122\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1010 net9 a_9227_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1011 tdc0.w_dly_sig\[104\] tdc0.w_dly_sig\[102\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1013 a_1570_13103# a_1297_13109# a_1485_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1015 VPWR a_17130_14709# a_17059_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1016 VGND tdc0.w_dly_sig_n\[126\] tdc0.w_dly_sig\[127\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1017 _023_ a_10446_6549# a_10226_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1018 VGND tdc0.w_dly_sig\[97\] tdc0.w_dly_sig\[99\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1019 a_17555_10383# a_17335_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1021 tdc0.w_dly_sig_n\[31\] tdc0.w_dly_sig\[31\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1023 VGND a_14611_13335# tdc0.o_result\[2\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1025 a_13989_5865# a_12999_5493# a_13863_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1026 a_9466_18111# a_9298_18365# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1027 a_12612_6895# net5 a_12516_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.107 ps=0.98 w=0.65 l=0.15
X1028 a_14611_13335# a_14707_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1030 a_11149_9545# tdc0.o_result\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1032 VGND tdc0.w_dly_sig_n\[9\] tdc0.w_dly_sig_n\[11\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1033 VPWR a_4111_10749# a_4279_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1034 a_14082_14191# a_13643_14197# a_13997_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1035 tdc0.o_result\[57\] a_6855_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1036 VGND tdc0.w_dly_sig\[119\] a_18673_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1037 tdc0.o_result\[66\] a_5199_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1038 a_17582_5309# a_17335_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1039 a_13914_3855# a_13599_4007# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1040 VGND tdc0.w_dly_sig\[69\] tdc0.w_dly_sig\[71\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1041 a_7308_10217# a_6909_9845# a_7182_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1042 a_3962_15279# a_3523_15285# a_3877_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1043 VGND a_14031_5461# a_13989_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1044 a_5970_12671# a_5802_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1045 a_16305_7779# _094_ a_16209_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1046 tdc0.w_dly_sig_n\[104\] tdc0.w_dly_sig\[104\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1047 a_3686_15101# a_3247_14735# a_3601_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1048 tdc0.o_result\[48\] a_2255_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1049 VGND a_17555_10071# tdc0.o_result\[121\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1050 a_10321_8751# tdc0.o_result\[30\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1051 tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1053 clknet_4_3_0_clk a_7286_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1054 VGND a_1830_9813# a_1788_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1055 a_2248_4943# a_1849_4943# a_2122_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1056 VPWR tdc0.w_dly_sig\[101\] tdc0.w_dly_sig_n\[101\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1057 tdc0.o_result\[83\] a_4647_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1058 a_11759_12381# a_11539_12393# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1059 a_3812_17999# a_3413_17999# a_3686_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1060 VGND a_7534_1109# a_7492_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1061 tdc0.w_dly_sig\[126\] tdc0.w_dly_sig\[124\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1062 a_12345_4719# _015_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X1063 a_14024_1513# a_13625_1141# a_13898_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1064 a_7967_5487# a_7185_5493# a_7883_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1065 VGND _003_ a_13690_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X1066 VGND a_9650_1791# a_9608_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1067 tdc0.w_dly_sig_n\[14\] tdc0.w_dly_sig_n\[12\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1068 tdc0.w_dly_sig_n\[80\] tdc0.w_dly_sig\[80\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1069 a_8527_10927# a_7663_10933# a_8270_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1071 a_7479_13103# net6 a_7561_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1072 VPWR tdc0.w_dly_sig\[123\] a_18397_14569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1073 VGND tdc0.w_dly_sig\[18\] tdc0.w_dly_sig\[20\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1074 tdc0.w_dly_sig\[108\] tdc0.w_dly_sig_n\[107\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1075 VPWR tdc0.w_dly_sig_n\[40\] tdc0.w_dly_sig_n\[42\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1076 a_13258_12015# a_13011_12393# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1077 a_1113_12021# a_947_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1079 a_14563_5487# _015_ a_14645_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1080 a_8197_10927# a_7663_10933# a_8102_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1081 VGND a_6522_6549# a_6480_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1082 a_4295_10927# a_3597_10933# a_4038_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1083 VGND tdc0.w_dly_sig\[4\] tdc0.w_dly_sig_n\[4\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1084 a_17525_16367# a_17187_16599# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1085 VGND a_2271_6575# a_2439_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1086 uo_out[7] a_11504_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1087 a_15565_7663# _025_ a_15419_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X1088 a_5667_18365# a_4885_17999# a_5583_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1089 a_9135_5487# _028_ a_9217_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1090 VGND tdc0.w_dly_sig\[74\] tdc0.w_dly_sig_n\[74\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1091 a_12552_9545# _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X1094 VGND a_5851_13335# _042_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1095 a_2497_14191# tdc0.w_dly_sig\[50\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1097 a_11057_17455# tdc0.o_result\[23\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1098 tdc0.o_result\[39\] a_9155_16341# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1099 a_9125_6575# tdc0.o_result\[76\] a_9043_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1100 VGND net10 a_7917_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1101 VPWR tdc0.w_dly_sig\[23\] tdc0.w_dly_sig\[25\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1102 a_17525_3133# a_17187_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1103 a_11892_11471# tdc0.o_result\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1104 a_2581_16911# a_1591_16911# a_2455_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1105 tdc0.w_dly_sig\[17\] tdc0.w_dly_sig\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1106 a_9397_9295# tdc0.w_dly_sig\[31\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1107 a_10137_2223# tdc0.o_result\[87\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1108 VGND tdc0.w_dly_sig\[105\] tdc0.w_dly_sig_n\[105\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1110 tdc0.w_dly_sig\[57\] tdc0.w_dly_sig\[55\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1111 a_5851_13335# tdc0.o_result\[38\] a_5997_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1113 tdc0.w_dly_sig_n\[107\] tdc0.w_dly_sig_n\[105\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1115 a_2355_6575# a_1573_6581# a_2271_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1117 tdc0.w_dly_sig\[59\] tdc0.w_dly_sig_n\[58\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1118 tdc0.w_dly_sig\[55\] tdc0.w_dly_sig_n\[54\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1119 VPWR tdc0.w_dly_sig_n\[93\] tdc0.w_dly_sig_n\[95\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1120 a_4881_4777# a_3891_4405# a_4755_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1121 tdc0.w_dly_sig\[43\] tdc0.w_dly_sig_n\[42\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1122 tdc0.w_dly_sig_n\[69\] tdc0.w_dly_sig_n\[67\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1123 tdc0.w_dly_sig_n\[19\] tdc0.w_dly_sig\[19\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1124 a_7515_9661# a_6817_9295# a_7258_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1125 a_13809_14197# a_13643_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1126 a_2539_17277# a_1757_16911# a_2455_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1127 VPWR tdc0.w_dly_sig_n\[77\] tdc0.w_dly_sig_n\[79\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1128 VPWR a_7331_16189# a_7499_16091# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1129 VPWR clknet_0_clk a_4176_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1130 tdc0.w_dly_sig\[58\] tdc0.w_dly_sig\[56\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1131 VPWR tdc0.w_dly_sig\[127\] tdc0.w_dly_sig\[129\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1132 clknet_4_0_0_clk a_4176_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1133 VGND tdc0.w_dly_sig\[50\] tdc0.w_dly_sig_n\[50\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1134 a_7534_1109# a_7366_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1135 _027_ a_9043_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1136 VGND tdc0.w_dly_sig_n\[2\] tdc0.w_dly_sig\[3\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1137 VPWR tdc0.w_dly_sig_n\[11\] tdc0.w_dly_sig_n\[13\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1138 a_5802_2045# a_5363_1679# a_5717_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1139 a_5786_5055# a_5618_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1140 a_16163_2045# a_15465_1679# a_15906_1791# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1141 a_17134_4943# a_16819_5095# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1142 tdc0.o_result\[62\] a_7775_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1143 clknet_4_15_0_clk a_16578_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1145 a_9677_11721# tdc0.o_result\[29\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1146 VGND a_2290_5055# a_2248_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1147 tdc0.w_dly_sig\[21\] tdc0.w_dly_sig_n\[20\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1148 a_14868_8751# tdc0.o_result\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X1150 VPWR tdc0.w_dly_sig_n\[6\] tdc0.w_dly_sig_n\[8\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1151 VGND a_17187_13799# tdc0.o_result\[123\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1152 a_10769_4943# tdc0.o_result\[71\] a_10423_5193# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1153 VGND tdc0.w_dly_sig_n\[72\] tdc0.w_dly_sig\[73\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1154 a_12867_11159# a_13151_11145# a_13086_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1155 VPWR a_12548_4917# clknet_4_8_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1156 a_14645_5487# tdc0.o_result\[96\] a_14563_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1157 tdc0.w_dly_sig\[49\] tdc0.w_dly_sig_n\[48\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1158 a_6262_12015# a_5823_12021# a_6177_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1159 VPWR tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1160 VPWR tdc0.w_dly_sig\[68\] tdc0.w_dly_sig_n\[68\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1161 a_6285_13423# net6 a_5851_13335# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1162 tdc0.o_result\[24\] a_15595_17429# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1163 a_18187_10901# ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1165 VPWR tdc0.w_dly_sig_n\[11\] tdc0.w_dly_sig\[12\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1166 tdc0.w_dly_sig_n\[112\] tdc0.w_dly_sig\[112\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1167 tdc0.w_dly_sig\[98\] tdc0.w_dly_sig_n\[97\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1168 a_11122_7637# a_10975_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X1169 tdc0.w_dly_sig\[16\] tdc0.w_dly_sig_n\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1170 tdc0.w_dly_sig\[121\] tdc0.w_dly_sig_n\[120\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1171 a_13511_10071# a_13795_10057# a_13730_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1172 VGND clknet_4_15_0_clk a_15207_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1174 VGND clknet_4_13_0_clk a_14563_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1175 VGND _005_ a_16166_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1176 tdc0.w_dly_sig\[45\] tdc0.w_dly_sig\[43\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1177 tdc0.w_dly_sig_n\[95\] tdc0.w_dly_sig_n\[93\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1178 VGND _083_ a_15162_5095# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1179 VPWR a_4463_10901# a_4379_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1180 VGND a_11403_13321# a_11410_13225# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1181 tdc0.w_dly_sig_n\[18\] tdc0.w_dly_sig\[18\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1182 VPWR a_14323_1135# a_14491_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1183 a_14323_1135# a_13625_1141# a_14066_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1184 VPWR tdc0.w_dly_sig_n\[29\] tdc0.w_dly_sig_n\[31\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1185 tdc0.w_dly_sig\[92\] tdc0.w_dly_sig\[90\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1186 a_18119_4617# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1187 a_7258_9407# a_7090_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1188 VGND a_5951_15101# a_6119_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1190 a_4054_3311# a_3781_3317# a_3969_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1191 a_16187_12533# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1192 VGND tdc0.w_dly_sig\[10\] tdc0.w_dly_sig_n\[10\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1193 a_8367_4617# clknet_4_2_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1194 a_10093_7983# _000_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.213 ps=1.3 w=0.65 l=0.15
X1195 _005_ a_10759_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1196 tdc0.w_dly_sig\[93\] tdc0.w_dly_sig_n\[92\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1198 tdc0.w_dly_sig\[67\] tdc0.w_dly_sig\[65\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1199 VPWR tdc0.w_dly_sig\[12\] tdc0.w_dly_sig\[14\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1200 a_11527_4399# _026_ a_11609_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1201 uo_out[4] a_14952_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1202 tdc0.w_dly_sig\[26\] tdc0.w_dly_sig_n\[25\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1203 a_10857_12809# _058_ a_10785_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1204 VPWR a_14287_7119# _003_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1205 VGND clknet_4_9_0_clk a_13551_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1206 VGND a_17567_17673# a_17574_17577# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1207 VPWR a_7286_7119# clknet_4_3_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1208 tdc0.w_dly_sig\[9\] tdc0.w_dly_sig\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1209 a_9715_4221# a_8933_3855# a_9631_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1210 tdc0.o_result\[46\] a_4279_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1211 VPWR a_15170_15253# a_15097_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1212 clknet_4_11_0_clk a_16762_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1213 VGND a_14157_4917# _017_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1214 tdc0.w_dly_sig_n\[58\] tdc0.w_dly_sig\[58\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1216 VGND _016_ a_10226_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X1217 tdc0.o_result\[100\] a_14031_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1218 VGND tdc0.w_dly_sig\[65\] tdc0.w_dly_sig_n\[65\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1220 a_3870_1135# a_3597_1141# a_3785_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1221 a_13863_3311# a_12999_3317# a_13606_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1222 tdc0.w_dly_sig_n\[68\] tdc0.w_dly_sig\[68\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1223 VGND a_2455_17277# a_2623_17179# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1224 a_8933_16189# a_8399_15823# a_8838_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1225 a_17753_4943# a_17206_5217# a_17406_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1226 tdc0.w_dly_sig_n\[70\] tdc0.w_dly_sig\[70\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1227 VPWR a_10598_14709# a_10527_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1228 VGND a_7442_3967# a_7400_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1229 VGND a_17102_1109# a_17060_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1230 a_1478_9661# a_1205_9295# a_1393_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1231 VGND tdc0.w_dly_sig_n\[16\] tdc0.w_dly_sig_n\[18\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1233 a_14926_13469# a_14611_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1234 a_5928_1679# a_5529_1679# a_5802_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1236 a_6169_4943# a_5179_4943# a_6043_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1237 _016_ _002_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1238 VGND tdc0.w_dly_sig\[11\] tdc0.w_dly_sig\[13\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1239 tdc0.w_dly_sig\[100\] tdc0.w_dly_sig\[98\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1240 a_18475_8029# a_18255_8041# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1241 a_15653_1679# tdc0.w_dly_sig\[105\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1242 VGND a_16727_18151# tdc0.o_result\[126\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1243 tdc0.w_dly_sig_n\[97\] tdc0.w_dly_sig_n\[95\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1244 tdc0.w_dly_sig\[22\] tdc0.w_dly_sig\[20\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1245 VGND a_17199_10357# a_17206_10657# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1246 a_8083_4631# a_8367_4617# a_8302_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1247 VGND clknet_4_6_0_clk a_5639_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1248 net6 a_8819_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1249 tdc0.w_dly_sig\[110\] tdc0.w_dly_sig_n\[109\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1250 VGND _010_ a_5985_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1251 a_11968_6031# net5 a_11872_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.107 ps=0.98 w=0.65 l=0.15
X1252 VPWR tdc0.w_dly_sig_n\[80\] tdc0.w_dly_sig\[81\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1253 VPWR tdc0.w_dly_sig\[85\] tdc0.w_dly_sig\[87\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1255 VPWR tdc0.w_dly_sig\[113\] tdc0.w_dly_sig_n\[113\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1256 _057_ a_10239_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1257 VGND ui_in[3] a_12999_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X1258 a_5802_12925# a_5529_12559# a_5717_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1259 VPWR a_4279_15003# a_4195_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1260 a_14323_1135# a_13459_1141# a_14066_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1261 VGND a_5291_13077# a_5249_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1262 a_5989_12021# a_5823_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1263 VPWR a_4095_8725# a_4011_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1264 tdc0.w_dly_sig_n\[0\] net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1265 VGND tdc0.w_dly_sig\[116\] tdc0.w_dly_sig\[118\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1266 _024_ a_7479_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1267 tdc0.w_dly_sig_n\[121\] tdc0.w_dly_sig\[121\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1268 a_7281_1135# tdc0.w_dly_sig\[92\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1269 a_9397_1679# tdc0.w_dly_sig\[96\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1270 VPWR a_13603_7093# net10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1271 a_17703_17833# a_17574_17577# a_17283_17687# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1272 a_15807_12711# a_15903_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1273 a_13783_18151# a_13879_17973# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1275 VGND tdc0.w_dly_sig\[75\] tdc0.w_dly_sig\[77\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1276 a_17950_17455# a_17703_17833# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1277 tdc0.w_dly_sig_n\[30\] tdc0.w_dly_sig_n\[28\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R7 VPWR tt_um_hpretl_tt06_tdc_14.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1278 a_7925_8751# tdc0.w_dly_sig\[34\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1279 tdc0.o_result\[72\] a_2071_11739# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1280 a_17210_2045# a_16937_1679# a_17125_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1281 a_3329_12015# tdc0.o_result\[74\] a_3247_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1282 VGND a_13479_2197# a_13437_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1283 VGND a_15906_10495# a_15864_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1284 VGND a_11403_12233# a_11410_12137# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1285 clknet_4_0_0_clk a_4176_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1286 a_8841_13109# a_8675_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1287 VGND tdc0.w_dly_sig_n\[64\] tdc0.w_dly_sig\[65\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R8 VGND uio_out[1] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1288 a_6269_6575# tdc0.w_dly_sig\[59\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1289 a_9113_16745# a_8123_16373# a_8987_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1291 VGND tdc0.w_dly_sig_n\[7\] tdc0.w_dly_sig_n\[9\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1292 tdc0.w_dly_sig\[39\] tdc0.w_dly_sig_n\[38\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1293 a_14093_6281# _013_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X1294 VPWR _012_ a_10321_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1295 a_6798_10901# a_6630_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1296 tdc0.w_dly_sig_n\[36\] tdc0.w_dly_sig_n\[34\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1297 a_17703_2767# a_17567_2741# a_17283_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1298 tdc0.w_dly_sig_n\[77\] tdc0.w_dly_sig_n\[75\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1299 tdc0.w_dly_sig\[13\] tdc0.w_dly_sig_n\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1300 VGND tdc0.w_dly_sig_n\[86\] tdc0.w_dly_sig\[87\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1301 VPWR tdc0.w_dly_sig\[76\] tdc0.w_dly_sig_n\[76\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1302 VPWR net1 tdc0.w_dly_sig_n\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1303 a_16155_14423# tdc0.o_result\[26\] a_16301_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1304 VGND a_3790_7119# clknet_4_1_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1305 VPWR a_8051_5461# a_7967_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1306 a_14250_14165# a_14082_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1307 VPWR tdc0.w_dly_sig\[112\] tdc0.w_dly_sig\[114\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1308 a_4732_17833# a_4333_17461# a_4606_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1309 VGND a_15235_5719# _085_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1310 a_7005_9295# tdc0.w_dly_sig\[61\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1311 clknet_4_4_0_clk a_3698_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1312 clknet_4_8_0_clk a_12548_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1313 VPWR tdc0.w_dly_sig\[117\] tdc0.w_dly_sig\[119\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1314 VPWR a_3348_13077# clknet_4_5_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1315 VPWR tdc0.w_dly_sig\[95\] tdc0.w_dly_sig_n\[95\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1316 tdc0.o_result\[11\] a_14583_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1317 tdc0.w_dly_sig_n\[5\] tdc0.w_dly_sig\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1318 VPWR tdc0.w_dly_sig\[128\] tdc0.w_dly_sig_n\[128\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1319 a_14082_14191# a_13809_14197# a_13997_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1320 VGND a_7856_14165# clknet_4_7_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1321 VGND clknet_4_3_0_clk a_5915_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1322 tdc0.o_result\[32\] a_7867_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1323 VGND a_11058_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1324 a_8286_12015# a_7847_12021# a_8201_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1325 tdc0.o_result\[107\] a_15595_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1326 VPWR tdc0.w_dly_sig\[108\] tdc0.w_dly_sig\[110\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1327 VPWR tdc0.w_dly_sig_n\[112\] tdc0.w_dly_sig_n\[114\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1328 VPWR tdc0.w_dly_sig_n\[86\] tdc0.w_dly_sig_n\[88\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1329 VGND tdc0.w_dly_sig_n\[56\] tdc0.w_dly_sig\[57\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1330 clknet_4_13_0_clk a_14388_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1331 a_10091_3311# a_9393_3317# a_9834_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1332 VPWR tdc0.w_dly_sig_n\[117\] tdc0.w_dly_sig_n\[119\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1333 tdc0.w_dly_sig\[93\] tdc0.w_dly_sig\[91\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1334 VGND a_12284_9545# uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1335 tdc0.w_dly_sig_n\[79\] tdc0.w_dly_sig_n\[77\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1336 VGND a_5970_1791# a_5928_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1337 VGND a_2198_8725# a_2156_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1338 VPWR tdc0.w_dly_sig\[76\] tdc0.w_dly_sig\[78\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1339 a_7825_6031# a_6835_6031# a_7699_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1341 VGND tdc0.w_dly_sig\[11\] tdc0.w_dly_sig_n\[11\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1342 tdc0.w_dly_sig_n\[21\] tdc0.w_dly_sig\[21\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1343 tdc0.w_dly_sig\[36\] tdc0.w_dly_sig\[34\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1344 a_18489_6953# a_17935_6793# a_18142_6852# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1346 tdc0.o_result\[93\] a_9431_1109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1347 tdc0.o_result\[56\] a_6395_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1348 a_16332_12015# _071_ a_16600_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1349 tdc0.w_dly_sig\[30\] tdc0.w_dly_sig\[28\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1350 VGND tdc0.o_result\[98\] a_15669_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1351 VGND tdc0.w_dly_sig\[116\] a_17385_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1352 a_16915_4917# a_17199_4917# a_17134_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1353 a_11023_14423# a_11119_14423# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1354 tdc0.w_dly_sig\[91\] tdc0.w_dly_sig\[89\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1355 a_1478_11837# a_1205_11471# a_1393_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1356 a_11539_12393# a_11410_12137# a_11119_12247# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1357 VGND tdc0.w_dly_sig_n\[109\] tdc0.w_dly_sig_n\[111\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1358 VGND a_14250_14165# a_14208_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1359 VGND a_7499_16091# a_7457_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1360 tdc0.w_dly_sig_n\[63\] tdc0.w_dly_sig_n\[61\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1361 a_2037_4943# tdc0.w_dly_sig\[80\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1362 a_6227_2045# a_5529_1679# a_5970_1791# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1363 VGND _097_ a_6467_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1364 _073_ a_10975_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1365 a_12118_9295# _076_ a_12284_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1366 VPWR tdc0.w_dly_sig\[31\] tdc0.w_dly_sig\[33\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1367 a_15462_15101# a_15023_14735# a_15377_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1368 VPWR tdc0.w_dly_sig_n\[104\] tdc0.w_dly_sig_n\[106\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1369 VGND a_10011_14887# tdc0.o_result\[15\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1370 VGND _067_ a_7755_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1371 VPWR a_16762_8207# clknet_4_11_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1372 VGND tdc0.w_dly_sig_n\[83\] tdc0.w_dly_sig_n\[85\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1373 a_16399_5487# net8 a_16181_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1374 tdc0.w_dly_sig\[70\] tdc0.w_dly_sig\[68\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1375 VGND a_8500_4917# clknet_4_2_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1376 VPWR _002_ a_9747_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X1377 tdc0.o_result\[73\] a_2623_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1378 VPWR tdc0.w_dly_sig_n\[4\] tdc0.w_dly_sig_n\[6\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1380 VPWR a_4130_15253# a_4057_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1381 a_10607_12809# _058_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1382 tdc0.w_dly_sig_n\[47\] tdc0.w_dly_sig\[47\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1383 VPWR a_4222_3285# a_4149_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1384 tdc0.w_dly_sig\[3\] tdc0.w_dly_sig\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1385 a_12058_4221# a_11785_3855# a_11973_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1386 a_8325_4399# a_7987_4631# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1387 a_11456_10927# _041_ a_11724_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1389 VPWR a_11122_7637# _029_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1390 a_10291_7983# _002_ a_10177_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.137 ps=1.07 w=0.65 l=0.15
X1391 a_8481_8457# tdc0.o_result\[92\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1392 VPWR tdc0.w_dly_sig\[53\] tdc0.w_dly_sig_n\[53\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1393 a_18234_3588# a_18027_3529# a_18410_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1394 tdc0.w_dly_sig_n\[88\] tdc0.w_dly_sig_n\[86\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1395 a_18318_6575# a_18071_6953# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1397 VPWR a_16331_10651# a_16247_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1398 a_3762_5461# a_3594_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1399 clknet_4_5_0_clk a_3348_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1400 tdc0.w_dly_sig\[111\] tdc0.w_dly_sig_n\[110\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1401 VGND clknet_4_0_0_clk a_1683_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1402 VPWR a_18027_12233# a_18034_12137# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1403 _022_ a_11214_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X1404 VPWR a_14163_17973# a_14170_18273# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1405 VGND tdc0.w_dly_sig_n\[88\] tdc0.w_dly_sig\[89\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1406 VPWR tdc0.w_dly_sig\[113\] tdc0.w_dly_sig\[115\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1407 uo_out[6] a_12376_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1408 tdc0.o_result\[19\] a_5751_18267# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1409 tdc0.o_result\[67\] a_4923_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1410 VGND a_14388_13621# clknet_4_13_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1411 tdc0.w_dly_sig_n\[122\] tdc0.w_dly_sig_n\[120\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1412 a_4606_6575# a_4167_6581# a_4521_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1413 a_6204_13647# a_5805_13647# a_6078_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1414 tdc0.w_dly_sig\[100\] tdc0.w_dly_sig_n\[99\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1415 tdc0.o_result\[91\] a_7959_1109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1416 a_13353_5487# tdc0.w_dly_sig\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1417 a_4521_17455# tdc0.w_dly_sig\[43\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1419 tdc0.w_dly_sig_n\[24\] tdc0.w_dly_sig_n\[22\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1420 tdc0.w_dly_sig\[76\] tdc0.w_dly_sig\[74\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1421 a_7791_1135# a_6927_1141# a_7534_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1422 a_2030_4399# a_1757_4405# a_1945_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1423 a_16248_9839# _005_ a_16332_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1424 a_8933_3855# a_8767_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1425 tdc0.w_dly_sig\[25\] tdc0.w_dly_sig\[23\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1426 VGND a_18234_3588# a_18163_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1427 a_13070_8207# a_12893_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1428 a_7515_9661# a_6651_9295# a_7258_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1429 a_6335_17973# a_6626_18273# a_6577_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1430 VPWR tdc0.w_dly_sig\[24\] tdc0.w_dly_sig\[26\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1431 VPWR a_6687_12015# a_6855_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1432 VGND tdc0.w_dly_sig_n\[39\] tdc0.w_dly_sig\[40\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1433 tdc0.w_dly_sig\[2\] tdc0.w_dly_sig_n\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1434 a_2603_12015# _026_ a_2685_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1435 a_7415_16189# a_6633_15823# a_7331_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1436 tdc0.w_dly_sig_n\[76\] tdc0.w_dly_sig\[76\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1437 VPWR a_1646_9407# a_1573_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1438 a_8013_12021# a_7847_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1440 tdc0.o_result\[8\] a_14675_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1441 VGND a_6687_12015# a_6855_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1442 tdc0.w_dly_sig_n\[113\] tdc0.w_dly_sig_n\[111\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1443 a_9389_6895# tdc0.o_result\[116\] a_9043_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1444 VPWR a_13151_11145# a_13158_11049# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1445 a_2122_1135# a_1849_1141# a_2037_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1446 VPWR tdc0.w_dly_sig_n\[44\] tdc0.w_dly_sig_n\[46\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1447 VGND clknet_4_6_0_clk a_7663_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1448 a_8723_4765# a_8503_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1449 _061_ a_10607_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1450 VGND a_11023_14423# tdc0.o_result\[14\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1451 a_18163_3689# a_18034_3433# a_17743_3543# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1452 VPWR tdc0.w_dly_sig\[105\] tdc0.w_dly_sig\[107\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1453 VPWR tdc0.w_dly_sig\[121\] a_18581_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1455 VPWR tdc0.w_dly_sig\[111\] tdc0.w_dly_sig\[113\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1456 tdc0.w_dly_sig_n\[76\] tdc0.w_dly_sig_n\[74\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1457 a_6779_6575# a_5915_6581# a_6522_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1458 VGND tdc0.w_dly_sig\[29\] a_14533_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1460 tdc0.w_dly_sig_n\[80\] tdc0.w_dly_sig_n\[78\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1461 tdc0.w_dly_sig\[19\] tdc0.w_dly_sig_n\[18\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1462 VGND tdc0.w_dly_sig_n\[60\] tdc0.w_dly_sig\[61\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1463 a_7189_3855# tdc0.w_dly_sig\[93\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1464 VGND a_17286_8725# a_17244_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1465 a_4061_13647# tdc0.w_dly_sig\[53\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1466 VPWR tdc0.w_dly_sig_n\[16\] tdc0.w_dly_sig\[17\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1467 VPWR tdc0.w_dly_sig\[78\] tdc0.w_dly_sig\[80\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1468 a_16071_18365# a_15207_17999# a_15814_18111# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1469 VGND clknet_4_5_0_clk a_1223_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1470 a_8953_7119# _001_ a_8853_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X1471 clknet_4_14_0_clk a_17314_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1472 VPWR a_14002_10116# a_13931_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1474 VGND tdc0.w_dly_sig\[49\] tdc0.w_dly_sig_n\[49\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1475 VPWR a_14491_1109# a_14407_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1476 tdc0.w_dly_sig\[104\] tdc0.w_dly_sig_n\[103\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1477 VGND a_3348_13077# clknet_4_5_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1478 tdc0.w_dly_sig_n\[30\] tdc0.w_dly_sig\[30\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1479 VGND tdc0.w_dly_sig\[126\] tdc0.w_dly_sig_n\[126\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1480 tdc0.w_dly_sig\[101\] tdc0.w_dly_sig_n\[100\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1481 a_12783_8029# net4 a_12692_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X1482 VGND tdc0.w_dly_sig_n\[49\] tdc0.w_dly_sig_n\[51\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1483 a_6619_17973# clknet_4_7_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1484 VGND tdc0.w_dly_sig\[90\] tdc0.w_dly_sig_n\[90\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1485 VGND tdc0.w_dly_sig\[93\] tdc0.w_dly_sig_n\[93\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1486 a_5943_7485# a_5161_7119# a_5859_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1487 VGND tdc0.w_dly_sig_n\[102\] tdc0.w_dly_sig_n\[104\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1488 tdc0.w_dly_sig\[20\] tdc0.w_dly_sig\[18\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1489 a_18410_3311# a_18163_3689# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1490 a_15511_4399# a_14729_4405# a_15427_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1491 a_17582_10749# a_17335_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1492 tdc0.w_dly_sig_n\[42\] tdc0.w_dly_sig_n\[40\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1493 a_7442_6143# a_7274_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1494 VPWR tdc0.w_dly_sig\[6\] a_13705_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1495 VGND clknet_4_3_0_clk a_6835_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1496 VGND clknet_4_10_0_clk a_16495_1141# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1497 VPWR tdc0.w_dly_sig_n\[23\] tdc0.w_dly_sig\[24\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1498 a_2603_12015# _026_ a_2685_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1499 a_1577_9839# tdc0.w_dly_sig\[78\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1500 a_12649_7814# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X1501 tdc0.w_dly_sig_n\[4\] tdc0.w_dly_sig\[4\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1502 tdc0.w_dly_sig\[2\] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1503 a_13165_5493# a_12999_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1504 a_10883_11721# _053_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1505 a_4613_13103# tdc0.w_dly_sig\[55\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1506 a_14664_6005# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1507 VGND a_11504_11445# uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1509 tdc0.w_dly_sig_n\[125\] tdc0.w_dly_sig\[125\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1510 a_15936_7119# _025_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1511 VPWR clknet_4_4_0_clk a_1039_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1512 VPWR tdc0.w_dly_sig_n\[50\] tdc0.w_dly_sig\[51\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1513 _070_ a_2603_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1514 a_11957_14569# a_11403_14409# a_11610_14468# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1515 VGND a_6430_11989# a_6388_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1516 tdc0.w_dly_sig\[35\] tdc0.w_dly_sig_n\[34\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1517 a_3870_10927# a_3597_10933# a_3785_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1518 a_12082_6031# a_11343_6031# a_11968_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.137 ps=1.07 w=0.65 l=0.15
X1519 a_4732_6953# a_4333_6581# a_4606_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1521 a_2631_5309# a_1849_4943# a_2547_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1522 a_1573_9661# a_1039_9295# a_1478_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1523 a_17493_9295# tdc0.w_dly_sig\[120\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1524 a_16600_9839# _101_ a_16332_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1525 a_5997_13103# net6 a_5851_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X1526 a_11333_8457# tdc0.o_result\[121\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1527 _098_ a_6099_16367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1528 a_11413_9295# tdc0.o_result\[14\] a_11067_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1529 VGND a_6211_5211# a_6169_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1530 tdc0.w_dly_sig_n\[38\] tdc0.w_dly_sig\[38\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1531 uo_out[2] a_14676_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1532 tdc0.w_dly_sig_n\[32\] tdc0.w_dly_sig\[32\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1533 VPWR _010_ a_4617_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1534 VGND tdc0.w_dly_sig_n\[26\] tdc0.w_dly_sig\[27\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1535 VPWR tdc0.w_dly_sig\[16\] a_10945_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1536 a_8933_3855# a_8767_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1537 tdc0.w_dly_sig\[7\] tdc0.w_dly_sig\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1538 a_18581_12393# a_18027_12233# a_18234_12292# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1540 a_10321_12335# tdc0.o_result\[79\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1541 a_6035_15101# a_5253_14735# a_5951_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1543 VGND a_16155_6183# _063_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1544 tdc0.o_result\[27\] a_16055_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1545 VGND tdc0.w_dly_sig_n\[46\] tdc0.w_dly_sig\[47\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1546 tdc0.w_dly_sig_n\[90\] tdc0.w_dly_sig_n\[88\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1547 VGND a_4222_3285# a_4180_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1548 tdc0.w_dly_sig_n\[84\] tdc0.w_dly_sig_n\[82\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1549 tdc0.w_dly_sig_n\[120\] tdc0.w_dly_sig_n\[118\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1550 VPWR tdc0.w_dly_sig\[2\] tdc0.w_dly_sig_n\[2\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1551 a_17187_2919# a_17283_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1552 a_8399_6575# _028_ a_8481_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1553 tdc0.w_dly_sig\[3\] tdc0.w_dly_sig_n\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1554 tdc0.w_dly_sig_n\[41\] tdc0.w_dly_sig\[41\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1555 VPWR tdc0.w_dly_sig\[127\] tdc0.w_dly_sig_n\[127\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1556 a_11785_3855# a_11619_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1557 VGND ui_in[5] a_12631_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X1558 VGND tdc0.w_dly_sig\[80\] tdc0.w_dly_sig_n\[80\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1559 a_3413_17999# a_3247_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1560 a_14151_10205# a_13931_10217# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1561 VPWR a_2198_4373# a_2125_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1562 VPWR tdc0.o_result\[58\] a_14093_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X1563 a_13603_7093# _009_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X1564 a_5717_1679# tdc0.w_dly_sig\[88\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1565 a_1903_11837# a_1205_11471# a_1646_11583# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1567 tdc0.w_dly_sig_n\[62\] tdc0.w_dly_sig\[62\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1568 VPWR clknet_4_5_0_clk a_1223_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1569 tdc0.w_dly_sig_n\[107\] tdc0.w_dly_sig\[107\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1571 VGND tdc0.w_dly_sig\[75\] tdc0.w_dly_sig_n\[75\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1572 a_1389_9845# a_1223_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1575 a_17406_10357# a_17199_10357# a_17582_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1576 VPWR tdc0.w_dly_sig_n\[19\] tdc0.w_dly_sig\[20\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1577 VGND a_16412_6549# clknet_4_10_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1578 VGND a_16394_12533# a_16323_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1579 a_11414_2045# a_11141_1679# a_11329_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1580 a_10595_7369# _002_ a_10401_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1581 VGND tdc0.w_dly_sig_n\[10\] tdc0.w_dly_sig\[11\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1582 VPWR tdc0.w_dly_sig\[8\] a_13429_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1583 a_17647_12247# a_17743_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1584 VPWR a_5031_6575# a_5199_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1585 tdc0.w_dly_sig_n\[1\] tdc0.w_dly_sig\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1586 _076_ a_11619_8867# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1588 a_17187_7119# a_16967_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1589 a_6706_4373# a_6538_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1590 VGND tdc0.o_result\[104\] a_16589_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1591 a_14591_6575# a_13809_6581# a_14507_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1592 a_17335_10383# a_17199_10357# a_16915_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1593 a_14917_15279# tdc0.w_dly_sig\[27\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1594 VPWR tdc0.w_dly_sig\[111\] tdc0.w_dly_sig_n\[111\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1595 a_14909_5807# tdc0.o_result\[8\] a_14563_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1596 a_6913_2223# tdc0.w_dly_sig\[90\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1598 VGND _074_ a_11619_8867# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1599 a_8503_4777# a_8367_4617# a_8083_4631# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1600 a_10791_16073# net6 a_10873_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1601 VPWR a_12226_3967# a_12153_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1602 VGND clknet_4_1_0_clk a_1591_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1603 a_3686_15101# a_3413_14735# a_3601_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1604 VPWR clknet_4_3_0_clk a_6835_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1606 VPWR a_11027_6005# net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1607 a_18489_6953# a_17942_6697# a_18142_6852# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1608 VGND tdc0.w_dly_sig\[110\] tdc0.w_dly_sig_n\[110\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1609 VGND a_17314_12559# clknet_4_14_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X1610 VPWR a_2750_14165# a_2677_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1611 VPWR a_9891_18267# a_9807_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1612 VPWR tdc0.o_result\[2\] a_14592_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1613 a_8841_17455# a_8307_17461# a_8746_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1614 a_15128_15657# a_14729_15285# a_15002_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1615 a_17463_17999# a_17243_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1616 VGND a_8711_12015# a_8879_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1617 a_17359_1135# a_16495_1141# a_17102_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1618 a_10029_6575# _003_ a_10226_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1619 clknet_4_2_0_clk a_8500_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X1620 a_16166_10159# _101_ a_16332_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1621 tdc0.o_result\[51\] a_2531_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1622 VPWR tdc0.w_dly_sig_n\[3\] tdc0.w_dly_sig\[4\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1623 a_15465_5193# _084_ a_15393_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1624 a_3229_8757# a_3063_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1626 VPWR tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1627 clknet_4_7_0_clk a_7856_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1628 a_17187_2919# a_17283_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1629 a_6963_4399# a_6265_4405# a_6706_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1630 tdc0.w_dly_sig_n\[85\] tdc0.w_dly_sig\[85\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1631 a_11957_13481# a_11403_13321# a_11610_13380# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1632 VGND tdc0.w_dly_sig\[84\] tdc0.w_dly_sig_n\[84\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1633 a_17187_13799# a_17283_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1634 VGND tdc0.w_dly_sig_n\[21\] tdc0.w_dly_sig_n\[23\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1635 a_5823_5487# net7 a_5905_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1636 VPWR a_4111_15101# a_4279_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1637 clknet_4_12_0_clk a_12548_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1638 a_17107_17973# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1639 tdc0.w_dly_sig_n\[74\] tdc0.w_dly_sig\[74\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1640 VPWR clknet_4_3_0_clk a_9043_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1641 VGND a_7867_6299# a_7825_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
R9 tt_um_hpretl_tt06_tdc_13.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1642 VPWR a_5951_4221# a_6119_4123# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1643 tdc0.o_result\[65\] a_7039_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1644 VPWR a_7683_9563# a_7599_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1645 VPWR tdc0.w_dly_sig_n\[27\] tdc0.w_dly_sig_n\[29\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1646 tdc0.w_dly_sig\[118\] tdc0.w_dly_sig_n\[117\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1647 VPWR a_2290_1109# a_2217_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1648 a_2125_4399# a_1591_4405# a_2030_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1649 VGND a_2715_1109# a_2673_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1650 a_17065_18365# a_16727_18151# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1651 a_6871_8573# a_6173_8207# a_6614_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1653 VGND tdc0.w_dly_sig_n\[94\] tdc0.w_dly_sig\[95\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1655 VGND a_2823_3311# a_2991_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1656 VPWR a_6947_6549# a_6863_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1657 tdc0.w_dly_sig_n\[0\] net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1658 VGND a_9631_4221# a_9799_4123# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1660 a_2217_3133# a_1683_2767# a_2122_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1661 VPWR a_17774_16644# a_17703_16745# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1662 VPWR _028_ a_8481_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1663 clknet_4_7_0_clk a_7856_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1664 a_11372_10927# _005_ a_11456_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1665 VGND a_14664_6005# clknet_4_9_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1667 tdc0.w_dly_sig\[13\] tdc0.w_dly_sig\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1668 tdc0.w_dly_sig\[103\] tdc0.w_dly_sig_n\[102\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1669 VPWR tdc0.w_dly_sig\[87\] tdc0.w_dly_sig\[89\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1670 VPWR tdc0.w_dly_sig\[9\] tdc0.w_dly_sig_n\[9\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1671 clknet_0_clk a_11058_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1672 a_11785_3855# a_11619_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1673 a_11311_2741# clknet_4_8_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1674 VGND tdc0.w_dly_sig_n\[56\] tdc0.w_dly_sig_n\[58\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1675 VPWR a_5583_18365# a_5751_18267# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1676 VGND a_17774_17732# a_17703_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1677 a_13534_10927# a_13287_11305# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1678 VGND tdc0.w_dly_sig\[112\] tdc0.w_dly_sig_n\[112\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1679 a_13947_6183# tdc0.o_result\[58\] a_14093_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X1681 clknet_4_3_0_clk a_7286_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1682 a_17743_3543# a_18034_3433# a_17985_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1684 a_18325_8751# _015_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X1685 a_2447_10927# a_1665_10933# a_2363_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1686 a_10975_17455# _029_ a_11057_17775# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1687 tdc0.w_dly_sig\[63\] tdc0.w_dly_sig_n\[62\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1688 a_17033_8751# tdc0.w_dly_sig\[118\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1689 VGND a_8454_11989# a_8412_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1690 a_12153_4221# a_11619_3855# a_12058_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1692 a_11504_11445# _005_ a_12326_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1693 a_17038_7093# a_16838_7393# a_17187_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1694 VPWR tdc0.w_dly_sig_n\[18\] tdc0.w_dly_sig_n\[20\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1695 VGND tdc0.w_dly_sig_n\[98\] tdc0.w_dly_sig_n\[100\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1696 a_5583_18365# a_4885_17999# a_5326_18111# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1697 a_17962_3677# a_17647_3543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1698 VPWR net1 tdc0.w_dly_sig_n\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1699 VPWR a_13082_12292# a_13011_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1700 VPWR a_8914_17429# a_8841_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1701 VGND tdc0.w_dly_sig_n\[49\] tdc0.w_dly_sig\[50\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1704 a_1646_11583# a_1478_11837# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1705 VGND a_15807_12711# tdc0.o_result\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1706 VGND tdc0.w_dly_sig\[103\] a_11865_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1707 a_12633_4719# _025_ a_12199_4631# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1708 VPWR a_9006_1109# a_8933_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1709 a_16145_12925# a_15807_12711# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1710 _100_ a_2511_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1711 a_2984_17833# a_2585_17461# a_2858_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1713 VGND tdc0.w_dly_sig\[103\] tdc0.w_dly_sig_n\[103\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1714 VPWR tdc0.w_dly_sig_n\[99\] tdc0.w_dly_sig_n\[101\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1715 VPWR clknet_4_7_0_clk a_8675_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1716 VGND clknet_4_11_0_clk a_16679_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1717 a_11119_14423# a_11410_14313# a_11361_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1718 tdc0.o_result\[84\] a_4463_1109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1719 VPWR tdc0.w_dly_sig_n\[5\] tdc0.w_dly_sig_n\[7\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1720 a_8491_5487# _028_ a_8573_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1721 _097_ a_5823_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1722 VGND tdc0.w_dly_sig_n\[64\] tdc0.w_dly_sig_n\[66\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1723 tdc0.w_dly_sig_n\[111\] tdc0.w_dly_sig\[111\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1725 a_9411_2223# _028_ a_9493_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1726 VPWR a_9539_13103# a_9707_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1727 VGND a_18187_10901# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1728 tdc0.w_dly_sig\[80\] tdc0.w_dly_sig_n\[79\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1729 tdc0.w_dly_sig\[89\] tdc0.w_dly_sig\[87\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1730 a_5031_6575# a_4167_6581# a_4774_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1731 VGND a_9539_13103# a_9707_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1732 VPWR a_3348_13077# clknet_4_5_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1733 a_9677_11471# tdc0.o_result\[61\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1734 a_17567_17673# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1735 a_3597_10933# a_3431_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1737 VGND _023_ a_9481_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1738 tdc0.w_dly_sig_n\[16\] tdc0.w_dly_sig\[16\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1739 tdc0.w_dly_sig\[103\] tdc0.w_dly_sig\[101\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1740 VGND clk a_11058_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1741 a_4237_14735# a_3247_14735# a_4111_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1742 tdc0.o_result\[83\] a_4647_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1743 clknet_4_13_0_clk a_14388_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1744 tdc0.w_dly_sig\[32\] tdc0.w_dly_sig_n\[31\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1746 a_16639_14709# a_16923_14709# a_16858_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1748 VPWR tdc0.w_dly_sig_n\[93\] tdc0.w_dly_sig\[94\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1749 VPWR net4 a_11214_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X1750 tdc0.o_result\[21\] a_9891_18267# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1751 a_9757_14569# a_8767_14197# a_9631_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1752 a_16035_8457# _020_ a_16117_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1753 a_17059_14735# a_16930_15009# a_16639_14709# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1754 VPWR tdc0.w_dly_sig\[74\] tdc0.w_dly_sig\[76\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1755 tdc0.w_dly_sig_n\[119\] tdc0.w_dly_sig_n\[117\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1756 a_9485_7485# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X1757 a_7055_10927# a_6357_10933# a_6798_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1758 a_15097_4399# a_14563_4405# a_15002_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1759 a_16127_7779# _093_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1760 VGND a_8178_8725# a_8136_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1761 VPWR tdc0.w_dly_sig\[64\] tdc0.w_dly_sig_n\[64\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1762 a_13358_11204# a_13151_11145# a_13534_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1763 tdc0.w_dly_sig_n\[32\] tdc0.w_dly_sig_n\[30\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1764 tdc0.w_dly_sig\[26\] tdc0.w_dly_sig\[24\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1765 VGND tdc0.w_dly_sig\[63\] tdc0.w_dly_sig_n\[63\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1766 VGND a_4176_6005# clknet_4_0_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1768 tdc0.w_dly_sig_n\[11\] tdc0.w_dly_sig\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1769 VGND tdc0.w_dly_sig\[82\] tdc0.w_dly_sig\[84\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1771 a_17647_3543# a_17743_3543# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1772 _092_ a_8399_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1773 a_11361_13103# a_11023_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1774 a_3877_15279# tdc0.w_dly_sig\[45\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1775 VGND tdc0.w_dly_sig_n\[58\] tdc0.w_dly_sig_n\[60\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1776 a_11311_2741# clknet_4_8_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1777 a_17635_2045# a_16937_1679# a_17378_1791# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1778 VPWR tdc0.w_dly_sig\[6\] tdc0.w_dly_sig\[8\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1779 VPWR a_11582_1791# a_11509_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1780 VPWR clknet_4_10_0_clk a_15299_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1781 VGND tdc0.w_dly_sig_n\[90\] tdc0.w_dly_sig_n\[92\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1782 VGND a_16762_8207# clknet_4_11_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1783 VPWR a_11023_14423# tdc0.o_result\[14\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1784 a_1849_4943# a_1683_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1785 VPWR _007_ a_11333_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1786 a_8477_16367# tdc0.w_dly_sig\[40\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1787 a_4088_15657# a_3689_15285# a_3962_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1788 tdc0.w_dly_sig\[17\] tdc0.w_dly_sig_n\[16\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1789 a_17385_7119# a_16831_7093# a_17038_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1790 a_9539_13103# a_8675_13109# a_9282_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1791 a_6467_10633# _098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1792 a_12199_4631# tdc0.o_result\[113\] a_12345_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1793 tdc0.w_dly_sig\[119\] tdc0.w_dly_sig_n\[118\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1794 VPWR a_17314_12559# clknet_4_14_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1795 VGND tdc0.w_dly_sig\[94\] tdc0.w_dly_sig_n\[94\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1796 a_3601_10383# tdc0.w_dly_sig\[54\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1797 VPWR clknet_0_clk a_3790_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1798 a_6353_12559# a_5363_12559# a_6227_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1799 tdc0.w_dly_sig\[78\] tdc0.w_dly_sig\[76\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1801 a_1297_13109# a_1131_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1802 VGND tdc0.w_dly_sig\[29\] tdc0.w_dly_sig_n\[29\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1803 VGND clknet_4_0_0_clk a_3615_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1804 VGND tdc0.w_dly_sig_n\[114\] tdc0.w_dly_sig_n\[116\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1805 VPWR tdc0.w_dly_sig_n\[14\] tdc0.w_dly_sig_n\[16\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1806 VGND a_7883_5487# a_8051_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1807 tdc0.w_dly_sig_n\[117\] tdc0.w_dly_sig_n\[115\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1808 VGND tdc0.w_dly_sig\[72\] tdc0.w_dly_sig_n\[72\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1809 a_6181_16687# tdc0.o_result\[43\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1810 VGND a_14186_3829# a_14115_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1811 tdc0.w_dly_sig\[78\] tdc0.w_dly_sig_n\[77\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1813 VPWR net10 a_9401_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1814 a_17283_17687# a_17574_17577# a_17525_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1815 a_15575_6281# _063_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1816 VGND a_15595_15253# a_15553_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1817 VPWR a_17527_1109# a_17443_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1818 tdc0.w_dly_sig_n\[53\] tdc0.w_dly_sig\[53\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1819 VPWR a_12199_4631# _080_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X1821 a_7917_16911# tdc0.o_result\[16\] a_7571_17161# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1822 tdc0.w_dly_sig\[47\] tdc0.w_dly_sig\[45\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1823 VPWR tdc0.w_dly_sig_n\[23\] tdc0.w_dly_sig_n\[25\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1824 a_9374_3967# a_9206_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1825 VGND a_10759_8181# _005_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1826 a_15853_7369# tdc0.o_result\[115\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1827 uo_out[1] a_12284_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1828 tdc0.o_result\[72\] a_2071_11739# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1829 tdc0.w_dly_sig\[6\] tdc0.w_dly_sig\[4\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1831 VPWR tdc0.w_dly_sig_n\[65\] tdc0.w_dly_sig\[66\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1832 a_13415_10071# a_13511_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1833 VPWR tdc0.w_dly_sig\[114\] a_17753_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1834 a_14707_13335# a_14991_13321# a_14926_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1835 clknet_4_3_0_clk a_7286_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1836 tdc0.w_dly_sig\[125\] tdc0.w_dly_sig_n\[124\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1837 VGND tdc0.w_dly_sig\[81\] tdc0.w_dly_sig_n\[81\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1838 a_5905_5807# tdc0.o_result\[67\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1839 tdc0.w_dly_sig_n\[109\] tdc0.w_dly_sig_n\[107\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1840 a_6549_7369# tdc0.o_result\[80\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1841 a_12613_2229# a_12447_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1842 a_15127_13481# a_14998_13225# a_14707_13335# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1843 a_9114_13103# a_8841_13109# a_9029_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1844 VGND a_5031_17455# a_5199_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1846 VGND clknet_4_1_0_clk a_1039_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1847 a_3413_10383# a_3247_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1848 a_15738_2045# a_15465_1679# a_15653_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1849 VGND a_5859_7485# a_6027_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1851 a_15347_13469# a_15127_13481# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1852 tdc0.w_dly_sig\[40\] tdc0.w_dly_sig_n\[39\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1853 a_1386_12015# a_947_12021# a_1301_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1854 VGND clknet_4_6_0_clk a_7847_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1857 a_14917_17455# tdc0.w_dly_sig\[25\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1858 a_18397_14569# a_17850_14313# a_18050_14468# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1859 tdc0.w_dly_sig\[63\] tdc0.w_dly_sig\[61\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1860 tdc0.w_dly_sig_n\[46\] tdc0.w_dly_sig_n\[44\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1861 VPWR net28 a_12893_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X1862 VGND a_6826_17973# a_6755_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1863 a_4881_1679# a_3891_1679# a_4755_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1865 tdc0.w_dly_sig_n\[13\] tdc0.w_dly_sig_n\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1866 tdc0.w_dly_sig_n\[33\] tdc0.w_dly_sig\[33\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1867 VPWR a_7223_10901# a_7139_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1868 VGND tdc0.w_dly_sig\[26\] tdc0.w_dly_sig\[28\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1869 a_14177_6575# a_13643_6581# a_14082_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1870 VPWR a_5199_6549# a_5115_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1871 VPWR tdc0.w_dly_sig_n\[59\] tdc0.w_dly_sig\[60\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1872 a_13011_12393# a_12882_12137# a_12591_12247# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1873 VPWR tdc0.w_dly_sig\[118\] tdc0.w_dly_sig_n\[118\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1874 VPWR clknet_4_7_0_clk a_8123_16373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1875 a_6871_8573# a_6007_8207# a_6614_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1876 uo_out[4] a_14952_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1877 a_14991_13321# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1878 VPWR a_18050_14468# a_17979_14569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1879 VGND a_14323_1135# a_14491_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1880 a_14349_10217# a_13795_10057# a_14002_10116# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1882 VGND tdc0.w_dly_sig_n\[70\] tdc0.w_dly_sig\[71\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1883 VPWR tdc0.w_dly_sig\[97\] tdc0.w_dly_sig_n\[97\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1884 a_14917_4399# tdc0.w_dly_sig\[108\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1885 VPWR a_13415_10071# tdc0.o_result\[6\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1886 a_7549_2601# a_6559_2229# a_7423_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1888 a_9555_4631# a_9839_4617# a_9774_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1889 VGND a_6671_13915# a_6629_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1890 tdc0.w_dly_sig_n\[49\] tdc0.w_dly_sig\[49\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1891 tdc0.w_dly_sig_n\[109\] tdc0.w_dly_sig\[109\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1892 a_14163_17973# clknet_4_13_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1893 a_14851_15823# a_14722_16097# a_14431_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1894 a_11149_9295# tdc0.o_result\[62\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1895 VPWR a_14675_14165# a_14591_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1896 VPWR tdc0.w_dly_sig_n\[128\] tdc0.w_dly_sig\[129\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1897 a_14375_5193# net8 a_14157_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1898 a_9347_16189# a_8565_15823# a_9263_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1899 tdc0.w_dly_sig_n\[96\] tdc0.w_dly_sig_n\[94\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1900 tdc0.w_dly_sig_n\[51\] tdc0.w_dly_sig_n\[49\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1901 VPWR tdc0.w_dly_sig_n\[100\] tdc0.w_dly_sig\[101\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1902 VGND a_15814_18111# a_15772_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1903 VGND _006_ a_14195_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X1904 VPWR tdc0.w_dly_sig\[51\] tdc0.w_dly_sig\[53\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1905 tdc0.w_dly_sig\[72\] tdc0.w_dly_sig_n\[71\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1906 a_17893_9839# a_17555_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1907 VGND a_13054_2197# a_13012_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1908 a_8753_1135# tdc0.w_dly_sig\[94\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1909 a_8933_14197# a_8767_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1910 a_5031_17455# a_4167_17461# a_4774_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1911 a_11225_5487# _001_ a_10975_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1912 VPWR tdc0.w_dly_sig_n\[17\] tdc0.w_dly_sig_n\[19\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1915 tdc0.w_dly_sig_n\[31\] tdc0.w_dly_sig_n\[29\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1916 a_17835_4631# a_18126_4521# a_18077_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1917 tdc0.w_dly_sig_n\[111\] tdc0.w_dly_sig_n\[109\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1918 _007_ a_9747_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X1919 tdc0.w_dly_sig_n\[34\] tdc0.w_dly_sig\[34\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1920 VGND tdc0.w_dly_sig\[109\] a_8921_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1921 a_11667_2767# a_11447_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1922 VGND _000_ a_8995_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1923 tdc0.w_dly_sig_n\[59\] tdc0.w_dly_sig\[59\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1924 VPWR a_6550_13103# clknet_4_6_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1925 tdc0.w_dly_sig\[14\] tdc0.w_dly_sig\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1926 clknet_4_0_0_clk a_4176_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X1927 a_12620_8029# a_12171_7663# a_12318_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1929 a_10873_15823# tdc0.o_result\[39\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1930 VGND a_6227_12925# a_6395_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1931 a_8730_16341# a_8562_16367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1934 VPWR a_13863_5487# a_14031_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1935 a_9213_17999# tdc0.w_dly_sig\[22\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1936 _038_ a_9411_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1937 VPWR tdc0.o_result\[101\] a_18325_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X1938 a_10140_11247# _022_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1939 VGND tdc0.w_dly_sig_n\[39\] tdc0.w_dly_sig_n\[41\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1940 VGND tdc0.w_dly_sig\[121\] tdc0.w_dly_sig_n\[121\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1941 tdc0.w_dly_sig\[85\] tdc0.w_dly_sig_n\[84\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1942 tdc0.w_dly_sig\[89\] tdc0.w_dly_sig_n\[88\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1943 tdc0.w_dly_sig\[102\] tdc0.w_dly_sig_n\[101\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1944 VGND a_13070_8207# a_13176_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1945 a_2106_10901# a_1938_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1946 VGND tdc0.w_dly_sig_n\[105\] tdc0.w_dly_sig\[106\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1947 VPWR a_12548_4917# clknet_4_8_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1948 a_12226_3967# a_12058_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1949 VPWR tdc0.w_dly_sig\[49\] tdc0.w_dly_sig\[51\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1950 VPWR tdc0.w_dly_sig\[52\] tdc0.w_dly_sig\[54\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1951 VGND tdc0.w_dly_sig_n\[55\] tdc0.w_dly_sig_n\[57\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1953 tdc0.o_result\[31\] a_9707_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1954 a_6265_4405# a_6099_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1955 a_9953_17455# net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X1957 a_11403_14409# clknet_4_12_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1958 VGND clknet_4_13_0_clk a_15023_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1959 VPWR tdc0.w_dly_sig_n\[110\] tdc0.w_dly_sig_n\[112\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1960 tdc0.w_dly_sig_n\[93\] tdc0.w_dly_sig_n\[91\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1961 a_7182_3311# a_6909_3317# a_7097_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1963 a_1830_14847# a_1662_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1964 tdc0.o_result\[31\] a_9707_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1965 tdc0.w_dly_sig_n\[67\] tdc0.w_dly_sig\[67\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1966 tdc0.w_dly_sig\[71\] tdc0.w_dly_sig\[69\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1967 tdc0.w_dly_sig_n\[2\] tdc0.w_dly_sig\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1968 tdc0.w_dly_sig\[95\] tdc0.w_dly_sig\[93\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1969 a_6771_12015# a_5989_12021# a_6687_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1970 _036_ a_9503_11043# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1971 VGND clknet_4_5_0_clk a_3247_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1972 VPWR tdc0.o_result\[4\] a_14868_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1973 VGND a_9366_10071# _081_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X1975 tdc0.w_dly_sig_n\[26\] tdc0.w_dly_sig_n\[24\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1976 VGND tdc0.w_dly_sig_n\[6\] tdc0.w_dly_sig\[7\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1977 VPWR tdc0.w_dly_sig\[104\] tdc0.w_dly_sig\[106\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1980 VPWR tdc0.w_dly_sig_n\[105\] tdc0.w_dly_sig_n\[107\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1981 a_13997_6575# tdc0.w_dly_sig\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1983 clknet_4_4_0_clk a_3698_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1984 VGND a_15162_5095# _086_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X1985 a_4146_14013# a_3707_13647# a_4061_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1986 tdc0.w_dly_sig\[11\] tdc0.w_dly_sig_n\[10\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1987 VGND a_9263_16189# a_9431_16091# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1988 clknet_4_6_0_clk a_6550_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1989 VGND a_17647_12247# tdc0.o_result\[120\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1990 a_9531_5095# tdc0.o_result\[109\] a_9677_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1991 a_4498_1791# a_4330_2045# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1992 clknet_4_2_0_clk a_8500_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1995 tdc0.w_dly_sig_n\[97\] tdc0.w_dly_sig\[97\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1997 VPWR a_2087_9839# a_2255_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1998 VPWR clknet_4_0_0_clk a_5363_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1999 VGND tdc0.w_dly_sig_n\[92\] tdc0.w_dly_sig_n\[94\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2000 clknet_4_2_0_clk a_8500_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2001 a_12771_11159# a_12867_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2002 VPWR tdc0.w_dly_sig_n\[68\] tdc0.w_dly_sig_n\[70\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2003 VPWR tdc0.w_dly_sig\[124\] a_18121_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2004 VGND a_9799_14165# a_9757_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2005 VGND tdc0.w_dly_sig_n\[32\] tdc0.w_dly_sig\[33\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2006 uo_out[6] a_12376_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2007 VGND clknet_4_3_0_clk a_7571_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2008 tdc0.o_result\[51\] a_2531_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2009 VGND tdc0.w_dly_sig\[17\] tdc0.w_dly_sig_n\[17\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2010 VGND a_18234_12292# a_18163_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2011 VPWR a_16187_12533# a_16194_12833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2012 VPWR tdc0.w_dly_sig_n\[15\] tdc0.w_dly_sig_n\[17\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2013 a_13438_5487# a_13165_5493# a_13353_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2014 a_5993_13647# tdc0.w_dly_sig\[37\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2015 tdc0.w_dly_sig_n\[90\] tdc0.w_dly_sig\[90\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2016 a_11518_2741# a_11318_3041# a_11667_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2017 a_8711_12015# a_8013_12021# a_8454_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2018 a_9797_4399# a_9459_4631# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2019 tdc0.w_dly_sig\[101\] tdc0.w_dly_sig\[99\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2020 VGND tdc0.w_dly_sig\[115\] tdc0.w_dly_sig\[117\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2021 VGND tdc0.w_dly_sig\[28\] tdc0.w_dly_sig\[30\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2022 VGND tdc0.w_dly_sig\[22\] tdc0.w_dly_sig_n\[22\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2023 VGND a_16543_14887# tdc0.o_result\[124\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2024 tdc0.w_dly_sig\[19\] tdc0.w_dly_sig\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2025 VPWR _016_ a_12171_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2026 VGND tdc0.w_dly_sig\[94\] tdc0.w_dly_sig\[96\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2027 a_16332_12015# _005_ a_16248_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2028 VPWR _057_ a_10857_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2029 tdc0.w_dly_sig\[67\] tdc0.w_dly_sig_n\[66\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2030 tdc0.w_dly_sig_n\[66\] tdc0.w_dly_sig\[66\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2031 VGND clknet_4_6_0_clk a_6651_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2033 a_12376_8751# _051_ a_12210_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2034 tdc0.o_result\[93\] a_9431_1109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2035 a_9319_12015# _013_ a_9401_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2036 VPWR a_15906_1791# a_15833_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2037 a_7097_9839# tdc0.w_dly_sig\[63\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2038 VGND _047_ a_13091_7779# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X2040 a_16543_12559# a_16323_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2041 a_14519_17999# a_14299_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2042 tdc0.w_dly_sig_n\[29\] tdc0.w_dly_sig_n\[27\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2043 a_13287_11305# a_13158_11049# a_12867_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2044 VPWR a_4038_1109# a_3965_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2045 VGND tdc0.w_dly_sig\[88\] tdc0.w_dly_sig_n\[88\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2046 a_2290_1109# a_2122_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2047 tdc0.w_dly_sig_n\[127\] tdc0.w_dly_sig_n\[125\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2048 a_11839_2045# a_11141_1679# a_11582_1791# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2049 _094_ a_16022_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X2050 VGND clknet_4_10_0_clk a_15299_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2051 a_11058_9839# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2052 a_6467_10633# _100_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2053 tdc0.w_dly_sig\[86\] tdc0.w_dly_sig\[84\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2054 VPWR tdc0.w_dly_sig\[51\] tdc0.w_dly_sig_n\[51\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2055 a_7173_17999# a_6619_17973# a_6826_17973# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2056 a_13599_14887# a_13695_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2057 VGND _085_ a_15162_5095# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X2058 VGND a_3927_8751# a_4095_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2059 VGND a_16163_10749# a_16331_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2060 VPWR tdc0.w_dly_sig_n\[54\] tdc0.w_dly_sig_n\[56\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2061 tdc0.w_dly_sig_n\[34\] tdc0.w_dly_sig_n\[32\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2062 VGND a_6550_13103# clknet_4_6_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X2063 VPWR clknet_4_13_0_clk a_15023_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2064 VPWR tdc0.w_dly_sig_n\[92\] tdc0.w_dly_sig\[93\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2065 a_6227_2045# a_5363_1679# a_5970_1791# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2066 tdc0.w_dly_sig\[41\] tdc0.w_dly_sig\[39\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2067 VGND a_6043_5309# a_6211_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2068 VPWR _018_ a_15220_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2069 VGND a_8695_10901# a_8653_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2070 a_11456_10927# _005_ a_11372_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2071 VPWR tdc0.o_result\[126\] a_16301_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X2072 VPWR a_13183_6583# _002_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2073 VPWR clknet_4_3_0_clk a_7019_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
R10 tt_um_hpretl_tt06_tdc_21.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2074 VPWR tdc0.w_dly_sig\[40\] tdc0.w_dly_sig\[42\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2075 a_6538_4399# a_6099_4405# a_6453_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2076 VGND tdc0.w_dly_sig_n\[66\] tdc0.w_dly_sig_n\[68\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2077 _050_ a_11527_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2078 a_8009_5865# a_7019_5493# a_7883_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2079 VGND a_16762_8207# clknet_4_11_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X2080 VGND a_13919_7119# _001_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2081 tdc0.w_dly_sig\[37\] tdc0.w_dly_sig_n\[36\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2082 VGND a_2255_15003# a_2213_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2083 a_6826_17973# a_6619_17973# a_7002_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2084 a_12326_11721# tdc0.o_result\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X2085 a_17502_2767# a_17187_2919# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2086 VPWR tdc0.w_dly_sig_n\[85\] tdc0.w_dly_sig\[86\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2087 VGND a_8051_5461# a_8009_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2088 a_5694_3967# a_5526_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2089 a_1849_1141# a_1683_1141# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2090 a_6446_8573# a_6007_8207# a_6361_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2091 tdc0.w_dly_sig\[50\] tdc0.w_dly_sig_n\[49\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2093 tdc0.w_dly_sig\[127\] tdc0.w_dly_sig_n\[126\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2094 a_15565_7663# _020_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2095 a_13151_11145# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2096 a_11338_13469# a_11023_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2097 VPWR tdc0.w_dly_sig_n\[124\] tdc0.w_dly_sig_n\[126\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2099 tdc0.w_dly_sig\[79\] tdc0.w_dly_sig_n\[78\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2100 a_11865_2767# a_11311_2741# a_11518_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2101 a_17578_9661# a_17305_9295# a_17493_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2102 VGND _001_ _023_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2103 _020_ a_8543_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X2104 a_7274_6397# a_7001_6031# a_7189_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2105 VGND a_12495_12247# tdc0.o_result\[7\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2106 a_11027_6005# _019_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2107 a_4330_4399# a_4057_4405# a_4245_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2108 a_4111_10749# a_3413_10383# a_3854_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2109 VGND a_1811_12015# a_1979_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2110 _029_ a_11122_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2111 a_15833_2045# a_15299_1679# a_15738_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2112 VGND tdc0.w_dly_sig\[14\] tdc0.w_dly_sig_n\[14\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2113 tdc0.w_dly_sig\[90\] tdc0.w_dly_sig\[88\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2114 net1 a_18187_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2115 a_17502_17821# a_17187_17687# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2116 tdc0.w_dly_sig_n\[70\] tdc0.w_dly_sig_n\[68\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2117 tdc0.w_dly_sig_n\[55\] tdc0.w_dly_sig_n\[53\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2118 a_8914_17429# a_8746_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2119 a_2397_6953# a_1407_6581# a_2271_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2120 clknet_4_13_0_clk a_14388_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2121 VPWR a_14186_14709# a_14115_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2122 a_13979_3829# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2123 a_11141_1679# a_10975_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2124 tdc0.w_dly_sig\[70\] tdc0.w_dly_sig_n\[69\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2125 VPWR a_18119_7881# a_18126_7785# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2126 a_3321_5493# a_3155_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2127 a_13054_2197# a_12886_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2128 a_9401_12015# tdc0.o_result\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2129 a_13690_7895# _002_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X2130 _018_ a_14195_8867# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X2131 a_16377_7779# _093_ a_16305_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2132 a_1393_11471# tdc0.w_dly_sig\[73\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2133 tdc0.o_result\[52\] a_4739_13915# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2134 a_10401_2543# tdc0.o_result\[87\] a_10055_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2135 tdc0.w_dly_sig_n\[84\] tdc0.w_dly_sig\[84\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2136 VGND a_4176_6005# clknet_4_0_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2138 VPWR a_7350_3285# a_7277_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2139 VPWR tdc0.w_dly_sig\[8\] tdc0.w_dly_sig_n\[8\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2141 VPWR _010_ a_10977_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2142 VGND a_8500_4917# clknet_4_2_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2143 a_3091_14191# a_2309_14197# a_3007_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2144 tdc0.o_result\[107\] a_15595_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2145 a_1757_4405# a_1591_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2146 a_1646_9407# a_1478_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2147 VPWR tdc0.w_dly_sig\[86\] tdc0.w_dly_sig\[88\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2148 net11 a_14195_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X2149 a_17134_10383# a_16819_10535# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2150 VPWR tdc0.w_dly_sig_n\[48\] tdc0.w_dly_sig_n\[50\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2151 a_6798_10901# a_6630_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2152 VPWR tdc0.w_dly_sig\[54\] tdc0.w_dly_sig\[56\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2153 a_2455_17277# a_1757_16911# a_2198_17023# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2154 a_6664_4777# a_6265_4405# a_6538_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2156 a_1646_9407# a_1478_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2157 VPWR tdc0.w_dly_sig_n\[0\] tdc0.w_dly_sig_n\[2\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2158 a_6035_4221# a_5253_3855# a_5951_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2159 a_17801_14191# a_17463_14423# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2161 VPWR tdc0.w_dly_sig\[125\] a_17477_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2162 a_6998_2223# a_6725_2229# a_6913_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2163 tdc0.w_dly_sig_n\[116\] tdc0.w_dly_sig_n\[114\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2164 a_13695_14709# a_13979_14709# a_13914_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2165 tdc0.w_dly_sig_n\[125\] tdc0.w_dly_sig_n\[123\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2166 a_6630_10927# a_6357_10933# a_6545_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2167 VPWR a_17314_12559# clknet_4_14_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2168 tdc0.o_result\[17\] a_9339_17429# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2169 VGND _023_ a_8745_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2170 VGND net28 a_11321_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2171 VGND a_1554_11989# a_1512_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2172 a_17661_17999# a_17114_18273# a_17314_17973# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2173 clknet_4_5_0_clk a_3348_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X2174 tdc0.o_result\[17\] a_9339_17429# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2175 VGND net4 _006_ VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X2176 a_8010_8751# a_7737_8757# a_7925_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2177 VGND tdc0.w_dly_sig\[26\] tdc0.w_dly_sig_n\[26\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2178 a_9374_3967# a_9206_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2179 a_6572_8207# a_6173_8207# a_6446_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2180 VGND tdc0.w_dly_sig\[40\] tdc0.w_dly_sig_n\[40\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2181 tdc0.o_result\[35\] a_8051_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2182 a_5326_18111# a_5158_18365# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2183 tdc0.w_dly_sig\[129\] tdc0.w_dly_sig_n\[128\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2184 VPWR tdc0.w_dly_sig\[91\] tdc0.w_dly_sig\[93\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2185 VGND a_10515_7671# _000_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2186 a_15297_5193# _082_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X2187 tdc0.w_dly_sig_n\[16\] tdc0.w_dly_sig_n\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2188 a_10044_10383# tdc0.o_result\[53\] a_9741_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X2189 VPWR a_13606_5461# a_13533_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2190 VPWR a_13947_6183# _083_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X2191 tdc0.w_dly_sig\[77\] tdc0.w_dly_sig\[75\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2192 tdc0.w_dly_sig\[23\] tdc0.w_dly_sig\[21\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2193 a_11338_12381# a_11023_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2194 a_1577_14735# tdc0.w_dly_sig\[49\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2195 VGND tdc0.w_dly_sig\[118\] tdc0.w_dly_sig\[120\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2196 a_9975_4777# a_9839_4617# a_9555_4631# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2197 VPWR tdc0.w_dly_sig\[121\] tdc0.w_dly_sig\[123\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2198 VGND a_12548_14165# clknet_4_12_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2199 VPWR a_3283_17455# a_3451_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2200 VGND tdc0.w_dly_sig_n\[111\] tdc0.w_dly_sig\[112\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2201 VPWR tdc0.w_dly_sig\[70\] tdc0.w_dly_sig\[72\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2202 VPWR tdc0.w_dly_sig_n\[116\] tdc0.w_dly_sig_n\[118\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2203 a_13353_8207# a_13176_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2204 VGND a_3283_17455# a_3451_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2206 a_17210_2045# a_16771_1679# a_17125_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2207 VGND a_2198_4373# a_2156_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2208 tdc0.w_dly_sig_n\[25\] tdc0.w_dly_sig_n\[23\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2210 clknet_4_13_0_clk a_14388_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2211 _009_ net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X2212 VGND a_13415_10071# tdc0.o_result\[6\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2213 clknet_4_11_0_clk a_16762_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2214 tdc0.w_dly_sig_n\[95\] tdc0.w_dly_sig\[95\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2215 tdc0.w_dly_sig\[90\] tdc0.w_dly_sig_n\[89\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2216 tdc0.w_dly_sig_n\[59\] tdc0.w_dly_sig_n\[57\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2217 VGND tdc0.w_dly_sig\[47\] tdc0.w_dly_sig\[49\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2218 a_13979_3829# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2219 VPWR _012_ a_13817_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2220 VPWR a_10011_14887# tdc0.o_result\[15\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2221 a_4111_18365# a_3247_17999# a_3854_18111# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2222 a_6725_2229# a_6559_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2223 a_17199_4917# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2224 tdc0.w_dly_sig_n\[72\] tdc0.w_dly_sig_n\[70\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2225 a_16741_12559# a_16194_12833# a_16394_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2226 VPWR tdc0.w_dly_sig_n\[13\] tdc0.w_dly_sig\[14\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2227 tdc0.w_dly_sig_n\[66\] tdc0.w_dly_sig_n\[64\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2228 VPWR clknet_4_4_0_clk a_3247_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2229 a_6909_3317# a_6743_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2230 a_3785_1135# tdc0.w_dly_sig\[85\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2231 VPWR a_4498_4373# a_4425_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2232 VGND a_16451_7271# tdc0.o_result\[115\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2233 a_9255_17455# a_8473_17461# a_9171_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2234 VPWR tdc0.o_result\[21\] a_9953_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X2236 tdc0.w_dly_sig\[76\] tdc0.w_dly_sig_n\[75\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2237 VGND a_14370_17973# a_14299_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2238 tdc0.w_dly_sig\[125\] tdc0.w_dly_sig\[123\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2239 _016_ _001_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2240 VPWR a_6395_1947# a_6311_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2241 VGND clknet_4_2_0_clk a_6099_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2242 VPWR a_15427_17455# a_15595_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2243 tdc0.w_dly_sig\[122\] tdc0.w_dly_sig_n\[121\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2245 VPWR tdc0.w_dly_sig\[113\] a_18581_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2246 VPWR _022_ a_2685_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2247 VGND a_15427_17455# a_15595_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2248 a_1205_9295# a_1039_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2249 a_3854_18111# a_3686_18365# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2250 VGND tdc0.w_dly_sig\[125\] tdc0.w_dly_sig_n\[125\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2251 _026_ a_11490_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2252 _019_ a_11642_5461# a_11422_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2253 clknet_4_9_0_clk a_14664_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2254 a_16166_10159# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2256 clknet_4_15_0_clk a_16578_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2257 a_2030_17277# a_1757_16911# a_1945_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2258 VGND tdc0.w_dly_sig\[114\] a_17753_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2259 VGND clknet_4_0_0_clk a_5363_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2260 tdc0.w_dly_sig_n\[101\] tdc0.w_dly_sig_n\[99\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2263 a_3283_17455# a_2419_17461# a_3026_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2264 VPWR a_13358_11204# a_13287_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2265 tdc0.w_dly_sig\[65\] tdc0.w_dly_sig_n\[64\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2266 VGND a_16187_12533# a_16194_12833# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2267 VGND a_7286_7119# clknet_4_3_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2269 tdc0.w_dly_sig_n\[40\] tdc0.w_dly_sig_n\[38\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2270 a_6633_15823# a_6467_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2271 a_11987_10633# _045_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2272 a_13533_5487# a_12999_5493# a_13438_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2273 tdc0.w_dly_sig\[88\] tdc0.w_dly_sig\[86\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2274 tdc0.w_dly_sig\[84\] tdc0.w_dly_sig\[82\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2276 VPWR tdc0.w_dly_sig_n\[35\] tdc0.w_dly_sig\[36\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2277 VGND tdc0.w_dly_sig\[12\] tdc0.w_dly_sig_n\[12\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2278 VGND a_6614_8319# a_6572_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2279 VPWR tdc0.w_dly_sig_n\[95\] tdc0.w_dly_sig\[96\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2280 a_9043_8457# _030_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2281 VGND a_14583_8475# a_14541_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2283 VPWR clknet_4_7_0_clk a_8767_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2284 tdc0.w_dly_sig_n\[19\] tdc0.w_dly_sig_n\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2285 VGND a_9807_17687# _032_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2286 VGND a_7350_3285# a_7308_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2287 VGND tdc0.w_dly_sig_n\[41\] tdc0.w_dly_sig_n\[43\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2288 VPWR a_17746_9407# a_17673_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2289 a_11957_13481# a_11410_13225# a_11610_13380# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2290 VPWR a_7442_6143# a_7369_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2291 a_3686_10749# a_3247_10383# a_3601_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2292 VGND a_9650_7637# _025_ VGND sky130_fd_pr__nfet_01v8 ad=0.213 pd=1.3 as=0.0878 ps=0.92 w=0.65 l=0.15
X2293 VPWR tdc0.w_dly_sig_n\[87\] tdc0.w_dly_sig_n\[89\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2294 VGND tdc0.w_dly_sig_n\[121\] tdc0.w_dly_sig_n\[123\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2295 VPWR a_13795_10057# a_13802_9961# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2296 a_10239_8751# _028_ a_10321_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2297 tdc0.w_dly_sig_n\[116\] tdc0.w_dly_sig\[116\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2298 a_12226_3967# a_12058_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2299 a_17336_1679# a_16937_1679# a_17210_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2300 a_1788_10217# a_1389_9845# a_1662_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2301 VPWR tdc0.w_dly_sig_n\[123\] tdc0.w_dly_sig\[124\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2302 VPWR tdc0.w_dly_sig\[119\] tdc0.w_dly_sig\[121\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2303 VPWR a_11610_13380# a_11539_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2304 a_7856_14165# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2305 tdc0.o_result\[19\] a_5751_18267# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2307 a_4425_4399# a_3891_4405# a_4330_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2308 VPWR a_12548_4917# clknet_4_8_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2309 a_12548_14165# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2310 a_17950_3133# a_17703_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2311 a_8481_8207# tdc0.o_result\[44\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2312 VGND a_11610_14468# a_11539_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2313 a_11527_4399# _026_ a_11609_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2314 tdc0.w_dly_sig_n\[43\] tdc0.w_dly_sig\[43\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2315 a_17283_17687# a_17567_17673# a_17502_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2316 VGND a_12518_7119# _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2317 VGND a_16578_13103# clknet_4_15_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2318 a_15741_18365# a_15207_17999# a_15646_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2319 VGND _023_ a_8837_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2320 a_16035_8457# _020_ a_16117_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2321 a_4145_5865# a_3155_5493# a_4019_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2322 VGND net3 a_12171_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2323 VPWR a_17567_13621# a_17574_13921# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2324 VGND _010_ a_9757_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2325 VPWR net5 a_12318_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X2326 a_11067_9545# _013_ a_11149_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2328 a_3785_10927# tdc0.w_dly_sig\[56\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2329 VPWR tdc0.o_result\[110\] a_15565_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X2330 a_4479_3311# a_3615_3317# a_4222_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2331 a_2290_2879# a_2122_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2332 tdc0.w_dly_sig_n\[81\] tdc0.w_dly_sig\[81\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2333 a_1757_9839# a_1223_9845# a_1662_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2334 VPWR a_11403_14409# a_11410_14313# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2335 VPWR clknet_4_4_0_clk a_1499_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2336 VGND tdc0.w_dly_sig_n\[103\] tdc0.w_dly_sig_n\[105\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2337 a_6687_12015# a_5823_12021# a_6430_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2338 VPWR _007_ a_10873_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2339 clknet_4_0_0_clk a_4176_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2340 tdc0.w_dly_sig_n\[82\] tdc0.w_dly_sig_n\[80\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2341 tdc0.w_dly_sig\[87\] tdc0.w_dly_sig_n\[86\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2342 tdc0.w_dly_sig_n\[102\] tdc0.w_dly_sig_n\[100\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2344 VGND tdc0.w_dly_sig\[123\] a_18397_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2345 tdc0.w_dly_sig\[123\] tdc0.w_dly_sig_n\[122\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2346 a_3601_14735# tdc0.w_dly_sig\[47\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2347 a_8859_6281# _020_ a_8941_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2348 VPWR tdc0.w_dly_sig\[48\] tdc0.w_dly_sig\[50\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2349 clknet_4_6_0_clk a_6550_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2351 VPWR a_3026_17429# a_2953_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2352 a_6357_12015# a_5823_12021# a_6262_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2353 tdc0.o_result\[84\] a_4463_1109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2354 a_17923_13647# a_17703_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2355 a_2290_1109# a_2122_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2356 VPWR tdc0.w_dly_sig_n\[71\] tdc0.w_dly_sig_n\[73\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2358 a_17673_9661# a_17139_9295# a_17578_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2359 VPWR clknet_4_10_0_clk a_16771_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2361 VGND _022_ a_2857_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2363 VGND net5 a_11642_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2364 VPWR net7 a_5169_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2365 a_6357_10933# a_6191_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2366 a_12886_2223# a_12447_2229# a_12801_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2368 _041_ a_11435_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X2369 tdc0.w_dly_sig\[29\] tdc0.w_dly_sig\[27\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2370 tdc0.w_dly_sig_n\[0\] net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2372 VGND a_7959_1109# a_7917_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2373 a_17870_10205# a_17555_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2374 clknet_4_1_0_clk a_3790_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2375 a_2313_3311# tdc0.w_dly_sig\[81\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2376 VPWR _006_ a_12574_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X2377 VPWR tdc0.w_dly_sig\[60\] tdc0.w_dly_sig_n\[60\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2378 a_9125_6575# tdc0.o_result\[116\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2379 VPWR net4 a_12263_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=2.12 as=0.109 ps=1.36 w=0.42 l=0.15
X2380 tdc0.w_dly_sig\[33\] tdc0.w_dly_sig_n\[32\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2381 a_2497_14191# tdc0.w_dly_sig\[50\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2382 a_16301_17455# _007_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2383 a_11141_1679# a_10975_1679# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2384 a_11943_17687# a_12039_17687# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2385 tdc0.w_dly_sig_n\[17\] tdc0.w_dly_sig_n\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2386 a_4111_10749# a_3247_10383# a_3854_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2387 VGND a_17378_1791# a_17336_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2388 clknet_4_15_0_clk a_16578_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2389 VGND tdc0.w_dly_sig\[2\] tdc0.w_dly_sig\[4\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2390 VPWR tdc0.w_dly_sig\[3\] a_15545_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2391 VPWR _067_ a_8005_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2392 a_13054_2197# a_12886_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2394 tdc0.w_dly_sig_n\[126\] tdc0.w_dly_sig_n\[124\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2395 VGND a_13358_11204# a_13287_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2396 a_17525_14013# a_17187_13799# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2397 a_3417_8751# tdc0.w_dly_sig\[71\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2398 VGND a_7607_9839# a_7775_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2399 tdc0.o_result\[77\] a_2255_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2400 _005_ a_10759_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2401 VGND tdc0.w_dly_sig\[57\] tdc0.w_dly_sig\[59\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2402 a_9206_14191# a_8933_14197# a_9121_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2403 tdc0.o_result\[90\] a_7775_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2404 VPWR clknet_0_clk a_3348_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2405 VPWR a_15814_18111# a_15741_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2406 a_16248_12015# tdc0.o_result\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X2407 a_5123_13103# a_4425_13109# a_4866_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2408 VGND tdc0.w_dly_sig\[98\] tdc0.w_dly_sig_n\[98\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2409 a_12552_9545# _081_ a_12284_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2410 VGND tdc0.w_dly_sig_n\[76\] tdc0.w_dly_sig_n\[78\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2411 a_7286_7119# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2412 a_2029_11471# a_1039_11471# a_1903_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2413 VPWR a_6227_12925# a_6395_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2414 a_9298_18365# a_8859_17999# a_9213_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2415 a_15630_14847# a_15462_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2416 a_5901_16911# tdc0.w_dly_sig\[41\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2417 a_11600_7983# net4 a_11504_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.107 ps=0.98 w=0.65 l=0.15
X2420 tdc0.w_dly_sig\[60\] tdc0.w_dly_sig\[58\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2422 a_18153_8207# _025_ a_17719_8359# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2423 VGND a_10091_3311# a_10259_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2424 a_16247_2045# a_15465_1679# a_16163_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2425 a_2030_8751# a_1757_8757# a_1945_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2426 tdc0.w_dly_sig\[33\] tdc0.w_dly_sig\[31\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2427 a_14415_8573# a_13551_8207# a_14158_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2428 VPWR tdc0.w_dly_sig\[27\] tdc0.w_dly_sig_n\[27\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2429 tdc0.w_dly_sig\[106\] tdc0.w_dly_sig_n\[105\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2430 VGND clknet_4_0_0_clk a_1591_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2431 a_7373_5487# tdc0.w_dly_sig\[35\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2432 VGND tdc0.w_dly_sig\[83\] tdc0.w_dly_sig_n\[83\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2434 VPWR tdc0.w_dly_sig_n\[99\] tdc0.w_dly_sig\[100\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2435 a_8005_12809# _068_ a_7933_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2436 a_5694_3967# a_5526_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2437 a_16543_14887# a_16639_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2438 tdc0.w_dly_sig\[42\] tdc0.w_dly_sig\[40\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2439 VPWR tdc0.w_dly_sig_n\[47\] tdc0.w_dly_sig\[48\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2440 VGND tdc0.w_dly_sig\[4\] tdc0.w_dly_sig\[6\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2441 VGND tdc0.w_dly_sig_n\[2\] tdc0.w_dly_sig_n\[4\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2443 VGND tdc0.w_dly_sig_n\[40\] tdc0.w_dly_sig\[41\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2444 tdc0.w_dly_sig\[110\] tdc0.w_dly_sig\[108\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2445 a_9503_11043# _033_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2446 VPWR tdc0.w_dly_sig\[80\] tdc0.w_dly_sig\[82\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2447 VPWR _066_ a_16600_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2448 VGND a_10446_6549# _023_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2450 VPWR clknet_4_5_0_clk a_2143_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2451 VGND tdc0.o_result\[22\] a_16589_17775# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2452 a_1788_14735# a_1389_14735# a_1662_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2453 a_17555_4943# a_17335_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2454 VGND tdc0.w_dly_sig\[64\] tdc0.w_dly_sig\[66\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2455 a_10175_3311# a_9393_3317# a_10091_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2456 tdc0.o_result\[79\] a_2715_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2457 a_13012_2601# a_12613_2229# a_12886_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2458 VGND tdc0.w_dly_sig\[35\] tdc0.w_dly_sig\[37\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2459 VGND tdc0.w_dly_sig\[15\] tdc0.w_dly_sig_n\[15\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2460 VGND a_2715_5211# a_2673_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2461 a_10137_2543# tdc0.o_result\[95\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2462 a_16733_5461# net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X2463 VPWR tdc0.w_dly_sig\[77\] tdc0.w_dly_sig_n\[77\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2464 VGND _005_ a_12118_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2465 VGND tdc0.o_result\[118\] a_15853_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2466 VPWR a_3007_14191# a_3175_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2467 VGND tdc0.w_dly_sig\[21\] a_12877_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2468 tdc0.w_dly_sig\[82\] tdc0.w_dly_sig_n\[81\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2470 tdc0.w_dly_sig\[5\] tdc0.w_dly_sig\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2471 a_5805_13647# a_5639_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2472 VGND a_14526_2197# a_14484_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2473 VGND tdc0.w_dly_sig\[99\] tdc0.w_dly_sig_n\[99\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2474 a_14952_8751# _031_ a_14786_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2475 a_15545_13481# a_14991_13321# a_15198_13380# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2476 VGND tdc0.w_dly_sig\[52\] tdc0.w_dly_sig_n\[52\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2477 a_17118_8751# a_16845_8757# a_17033_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2478 a_13165_5493# a_12999_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2479 tdc0.w_dly_sig\[18\] tdc0.w_dly_sig_n\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2480 a_6361_8207# tdc0.w_dly_sig\[66\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2481 VPWR tdc0.w_dly_sig\[33\] tdc0.w_dly_sig_n\[33\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2482 tdc0.w_dly_sig_n\[83\] tdc0.w_dly_sig_n\[81\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2483 VPWR a_3698_12559# clknet_4_4_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2484 VGND tdc0.w_dly_sig\[89\] tdc0.w_dly_sig_n\[89\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2487 VPWR net2 a_12518_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.165 ps=1.33 w=1 l=0.15
X2488 a_1811_12015# a_1113_12021# a_1554_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2489 VPWR _036_ a_11724_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2490 a_7097_3311# tdc0.w_dly_sig\[91\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2491 VPWR a_2547_1135# a_2715_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2492 VGND a_16332_12015# uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2493 a_7331_16189# a_6467_15823# a_7074_15935# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2494 VGND a_7074_15935# a_7032_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2495 VPWR tdc0.w_dly_sig_n\[106\] tdc0.w_dly_sig_n\[108\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2496 a_2547_1135# a_1849_1141# a_2290_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2497 VGND a_15419_7895# _045_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2498 a_5717_12559# tdc0.w_dly_sig\[57\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2499 a_17283_2741# a_17574_3041# a_17525_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2500 a_4146_14013# a_3873_13647# a_4061_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2501 VGND a_4176_6005# clknet_4_0_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2502 VPWR _022_ a_3329_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2503 tdc0.w_dly_sig_n\[22\] tdc0.w_dly_sig_n\[20\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2504 VGND tdc0.w_dly_sig\[56\] tdc0.w_dly_sig_n\[56\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2506 tdc0.o_result\[61\] a_8695_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2507 VPWR tdc0.w_dly_sig_n\[73\] tdc0.w_dly_sig\[74\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2508 a_8711_12015# a_7847_12021# a_8454_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2509 VGND tdc0.w_dly_sig\[53\] tdc0.w_dly_sig\[55\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2510 tdc0.w_dly_sig\[114\] tdc0.w_dly_sig\[112\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2511 VGND tdc0.w_dly_sig_n\[41\] tdc0.w_dly_sig\[42\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2512 a_8574_4676# a_8367_4617# a_8750_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2513 a_4535_8751# _022_ a_4617_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2514 a_5602_7231# a_5434_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2516 VGND tdc0.w_dly_sig\[31\] tdc0.w_dly_sig_n\[31\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2517 a_8381_12015# a_7847_12021# a_8286_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2518 a_7185_5493# a_7019_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2519 a_14611_13335# a_14707_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2520 VGND clknet_4_2_0_clk a_6743_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2521 clknet_4_8_0_clk a_12548_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2522 VPWR a_4647_3285# a_4563_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2523 tdc0.w_dly_sig\[96\] tdc0.w_dly_sig\[94\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2524 tdc0.w_dly_sig_n\[103\] tdc0.w_dly_sig_n\[101\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2525 VPWR a_13311_2223# a_13479_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2526 a_11359_4943# net4 a_11241_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.143 ps=1.09 w=0.65 l=0.15
X2527 VPWR net3 a_10515_7671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2529 tdc0.w_dly_sig_n\[8\] tdc0.w_dly_sig\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2530 a_11447_2767# a_11318_3041# a_11027_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2531 a_5709_17999# a_4719_17999# a_5583_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2532 VGND tdc0.w_dly_sig\[34\] tdc0.w_dly_sig_n\[34\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2533 a_12210_9071# tdc0.o_result\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2534 VGND tdc0.w_dly_sig\[5\] a_15453_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2535 a_7817_17833# a_7270_17577# a_7470_17732# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2536 VPWR tdc0.w_dly_sig\[13\] tdc0.w_dly_sig\[15\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2537 a_11119_14423# a_11403_14409# a_11338_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2538 a_5721_6281# tdc0.o_result\[66\] a_5639_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2539 VGND a_16055_15003# a_16013_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2540 VPWR a_7131_4373# a_7047_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2541 a_9397_9295# tdc0.w_dly_sig\[31\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2542 tdc0.w_dly_sig_n\[3\] tdc0.w_dly_sig\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2543 a_6077_3855# a_5087_3855# a_5951_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2544 VGND a_10931_2919# tdc0.o_result\[102\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2545 VGND tdc0.w_dly_sig\[19\] a_7173_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2546 tdc0.o_result\[92\] a_7867_4123# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2548 tdc0.w_dly_sig\[69\] tdc0.w_dly_sig\[67\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2550 a_9485_7485# a_9319_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X2551 VPWR clknet_0_clk a_17314_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2552 VGND clknet_4_9_0_clk a_14563_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2553 a_10147_7369# _001_ a_10401_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2554 tdc0.o_result\[26\] a_15595_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2555 VPWR a_16163_10749# a_16331_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2556 tdc0.w_dly_sig_n\[88\] tdc0.w_dly_sig\[88\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2558 uo_out[7] a_11504_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2559 tdc0.w_dly_sig_n\[101\] tdc0.w_dly_sig\[101\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2560 a_2455_4399# a_1591_4405# a_2198_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2561 tdc0.o_result\[79\] a_2715_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2562 VPWR clknet_4_2_0_clk a_6559_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2563 tdc0.w_dly_sig_n\[11\] tdc0.w_dly_sig_n\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2564 VPWR a_9171_17455# a_9339_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2565 tdc0.o_result\[67\] a_4923_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2566 a_17406_4917# a_17206_5217# a_17555_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2567 a_2547_3133# a_1683_2767# a_2290_2879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2568 VGND tdc0.w_dly_sig_n\[68\] tdc0.w_dly_sig\[69\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2569 tdc0.w_dly_sig\[74\] tdc0.w_dly_sig_n\[73\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2570 tdc0.w_dly_sig\[68\] tdc0.w_dly_sig_n\[67\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2571 tdc0.w_dly_sig\[115\] tdc0.w_dly_sig_n\[114\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2572 VPWR a_2198_8725# a_2125_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2573 a_7626_7637# a_7458_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2575 VPWR tdc0.w_dly_sig_n\[119\] tdc0.w_dly_sig_n\[121\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2577 tdc0.w_dly_sig_n\[40\] tdc0.w_dly_sig\[40\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2578 VPWR a_11159_4943# _013_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2579 VPWR a_8500_4917# clknet_4_2_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2581 tdc0.w_dly_sig_n\[128\] tdc0.w_dly_sig\[128\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2582 a_11435_10633# _040_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2584 VGND a_8500_4917# clknet_4_2_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2586 VGND tdc0.w_dly_sig_n\[48\] tdc0.w_dly_sig\[49\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2587 a_13606_3285# a_13438_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2588 VPWR tdc0.w_dly_sig_n\[35\] tdc0.w_dly_sig_n\[37\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2589 a_17647_3543# a_17743_3543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2590 tdc0.w_dly_sig\[123\] tdc0.w_dly_sig\[121\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2591 a_9121_3855# tdc0.w_dly_sig\[110\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2592 a_17651_10071# a_17935_10057# a_17870_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2593 VPWR tdc0.w_dly_sig_n\[9\] tdc0.w_dly_sig\[10\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2594 a_8750_4399# a_8503_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2595 a_13311_2223# a_12613_2229# a_13054_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2597 VGND a_11504_11445# uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2598 a_13813_1135# tdc0.w_dly_sig\[100\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2599 a_17406_10357# a_17206_10657# a_17555_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2601 VGND tdc0.w_dly_sig_n\[115\] tdc0.w_dly_sig\[116\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2602 _026_ a_11490_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X2603 VGND a_17567_13621# a_17574_13921# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2604 a_14676_12809# _091_ a_14510_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2606 tdc0.w_dly_sig\[47\] tdc0.w_dly_sig_n\[46\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2607 VGND tdc0.w_dly_sig\[100\] tdc0.w_dly_sig\[102\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2608 a_4698_13103# a_4259_13109# a_4613_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2609 VGND tdc0.w_dly_sig\[43\] tdc0.w_dly_sig\[45\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2611 a_7691_9839# a_6909_9845# a_7607_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2612 tdc0.o_result\[96\] a_14951_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2613 VGND _049_ a_13091_7779# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X2614 VPWR a_8454_11989# a_8381_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2615 a_14208_14569# a_13809_14197# a_14082_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2616 a_11057_8751# tdc0.o_result\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2617 VPWR a_10931_2919# tdc0.o_result\[102\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2618 VGND a_9531_5095# _035_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2619 VPWR a_9839_4617# a_9846_4521# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2620 tdc0.w_dly_sig_n\[127\] tdc0.w_dly_sig\[127\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2621 a_15511_15279# a_14729_15285# a_15427_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2622 VGND a_16412_6549# clknet_4_10_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2623 tdc0.w_dly_sig\[49\] tdc0.w_dly_sig\[47\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2624 VGND a_16071_18365# a_16239_18267# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2625 VGND tdc0.w_dly_sig\[55\] tdc0.w_dly_sig\[57\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2626 a_13863_3311# a_13165_3317# a_13606_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2627 a_7124_2601# a_6725_2229# a_6998_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2628 VGND tdc0.w_dly_sig_n\[97\] tdc0.w_dly_sig\[98\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2629 uo_out[2] a_14676_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2630 a_3594_5487# a_3321_5493# a_3509_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2631 a_14952_8751# _031_ a_15220_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2632 VGND tdc0.w_dly_sig_n\[58\] tdc0.w_dly_sig\[59\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2633 VPWR tdc0.w_dly_sig_n\[54\] tdc0.w_dly_sig\[55\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2634 a_3812_14735# a_3413_14735# a_3686_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2635 tdc0.o_result\[21\] a_9891_18267# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2636 a_7755_12809# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2637 VGND tdc0.o_result\[124\] a_15761_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2638 VPWR tdc0.w_dly_sig_n\[42\] tdc0.w_dly_sig\[43\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2639 _068_ a_7571_17161# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2640 VPWR _025_ a_9125_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2641 a_8399_8457# _029_ a_8481_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2642 tdc0.o_result\[82\] a_2715_1109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2643 VGND tdc0.w_dly_sig\[19\] tdc0.w_dly_sig_n\[19\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2644 tdc0.w_dly_sig_n\[15\] tdc0.w_dly_sig_n\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2645 VPWR a_14583_8475# a_14499_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2646 VGND tdc0.w_dly_sig\[90\] tdc0.w_dly_sig\[92\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2647 VGND tdc0.w_dly_sig\[101\] tdc0.w_dly_sig\[103\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2648 VGND a_3854_18111# a_3812_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2649 VPWR tdc0.w_dly_sig_n\[19\] tdc0.w_dly_sig_n\[21\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2650 _012_ a_12518_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2651 tdc0.o_result\[33\] a_8603_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2652 VGND clknet_4_10_0_clk a_16771_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2653 a_11518_2741# a_11311_2741# a_11694_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2654 VPWR a_7039_8475# a_6955_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2655 VGND a_7286_7119# clknet_4_3_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2657 a_12134_6549# a_12792_6549# a_12726_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2658 a_2125_8751# a_1591_8757# a_2030_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2659 a_11119_13335# a_11403_13321# a_11338_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2660 VGND tdc0.o_result\[3\] a_16166_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2661 tdc0.w_dly_sig\[105\] tdc0.w_dly_sig\[103\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2662 tdc0.o_result\[87\] a_6395_1947# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2663 VPWR tdc0.w_dly_sig_n\[20\] tdc0.w_dly_sig\[21\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2664 VGND a_2623_8725# a_2581_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2665 tdc0.w_dly_sig_n\[117\] tdc0.w_dly_sig\[117\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2666 VGND tdc0.w_dly_sig\[33\] tdc0.w_dly_sig\[35\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2667 a_17753_4943# a_17199_4917# a_17406_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2668 VGND clknet_4_7_0_clk a_6467_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2669 _040_ a_10147_16073# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2670 VGND tdc0.w_dly_sig_n\[113\] tdc0.w_dly_sig_n\[115\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2671 VGND tdc0.w_dly_sig\[71\] tdc0.w_dly_sig_n\[71\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2672 VGND a_5199_6549# a_5157_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2673 a_12810_12381# a_12495_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2674 a_9779_6575# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2675 VGND a_11582_1791# a_11540_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2676 a_13625_1141# a_13459_1141# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2677 a_13311_2223# a_12447_2229# a_13054_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2678 a_15377_14735# tdc0.w_dly_sig\[28\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2679 VPWR a_17187_13799# tdc0.o_result\[123\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2680 _021_ a_8859_6281# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2681 VGND clknet_4_11_0_clk a_17139_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2682 VPWR a_1830_14847# a_1757_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2683 a_12292_8751# _005_ a_12376_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2684 VPWR a_17286_8725# a_17213_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2685 tdc0.w_dly_sig\[95\] tdc0.w_dly_sig_n\[94\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2686 VGND a_17107_17973# a_17114_18273# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2688 VPWR net10 a_9227_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2689 a_10873_16073# tdc0.o_result\[127\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2690 _051_ a_13091_7779# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X2691 a_12516_6895# net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.114 ps=1 w=0.65 l=0.15
X2692 VGND tdc0.w_dly_sig_n\[32\] tdc0.w_dly_sig_n\[34\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2693 tdc0.w_dly_sig\[77\] tdc0.w_dly_sig_n\[76\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2694 tdc0.w_dly_sig_n\[123\] tdc0.w_dly_sig_n\[121\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2695 clknet_4_7_0_clk a_7856_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2696 a_11490_6005# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.175 ps=1.35 w=1 l=0.15
X2697 a_11565_6575# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X2698 tdc0.w_dly_sig_n\[60\] tdc0.w_dly_sig\[60\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2699 VGND a_3698_12559# clknet_4_4_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2700 tdc0.o_result\[38\] a_6119_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2701 VGND a_17719_8359# _052_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2702 a_14273_2223# tdc0.w_dly_sig\[97\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2703 tdc0.w_dly_sig\[124\] tdc0.w_dly_sig_n\[123\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2704 tdc0.w_dly_sig\[121\] tdc0.w_dly_sig\[119\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2705 VPWR tdc0.w_dly_sig_n\[14\] tdc0.w_dly_sig\[15\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2706 clknet_4_12_0_clk a_12548_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2707 a_16166_10159# _096_ a_16332_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2709 _000_ a_10515_7671# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2710 a_18087_9661# a_17305_9295# a_18003_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2711 VGND tdc0.w_dly_sig_n\[51\] tdc0.w_dly_sig_n\[53\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2713 VPWR tdc0.w_dly_sig\[109\] tdc0.w_dly_sig_n\[109\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2714 VPWR tdc0.w_dly_sig\[83\] tdc0.w_dly_sig\[85\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2715 a_13690_7895# _000_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X2716 tdc0.w_dly_sig_n\[114\] tdc0.w_dly_sig\[114\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2718 a_16209_7779# _095_ a_16127_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2719 a_13931_10217# a_13802_9961# a_13511_10071# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2720 VGND clknet_0_clk a_16578_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2721 a_9581_3311# tdc0.w_dly_sig\[95\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2722 a_17567_17673# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2724 clknet_4_9_0_clk a_14664_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2725 VPWR tdc0.w_dly_sig\[7\] tdc0.w_dly_sig\[9\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2726 tdc0.w_dly_sig_n\[9\] tdc0.w_dly_sig\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2727 tdc0.w_dly_sig\[51\] tdc0.w_dly_sig_n\[50\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2728 tdc0.w_dly_sig\[120\] tdc0.w_dly_sig\[118\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2729 VPWR a_6579_17179# a_6495_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2730 _022_ a_11214_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2731 _011_ a_13459_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2732 VPWR tdc0.w_dly_sig_n\[60\] tdc0.w_dly_sig_n\[62\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2733 a_17042_17999# a_16727_18151# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2734 a_12039_17687# a_12330_17577# a_12281_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2735 a_11694_3133# a_11447_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2736 VGND _000_ a_11473_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.213 pd=1.3 as=0.0878 ps=0.92 w=0.65 l=0.15
X2737 VGND tdc0.w_dly_sig\[58\] tdc0.w_dly_sig_n\[58\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2738 tdc0.w_dly_sig_n\[118\] tdc0.w_dly_sig_n\[116\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2739 a_1757_8757# a_1591_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2740 tdc0.o_result\[44\] a_4555_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2741 VGND clknet_4_8_0_clk a_13919_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2742 VPWR tdc0.w_dly_sig\[95\] tdc0.w_dly_sig\[97\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2744 a_4176_6005# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2745 tdc0.o_result\[47\] a_2623_17179# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2746 tdc0.o_result\[58\] a_6947_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2747 a_3247_12015# _026_ a_3329_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2748 clknet_4_2_0_clk a_8500_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2749 VGND tdc0.w_dly_sig\[17\] a_7817_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2750 tdc0.w_dly_sig\[79\] tdc0.w_dly_sig\[77\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2751 a_13541_8751# tdc0.o_result\[84\] a_13459_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2752 a_9125_9071# tdc0.o_result\[89\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2753 a_18027_3529# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2754 VGND a_7699_6397# a_7867_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2755 a_6388_12393# a_5989_12021# a_6262_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2757 a_6411_17277# a_5713_16911# a_6154_17023# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2758 VPWR a_5751_18267# a_5667_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2759 VGND a_1979_11989# a_1937_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2760 tdc0.w_dly_sig\[94\] tdc0.w_dly_sig\[92\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2761 VPWR tdc0.w_dly_sig\[20\] tdc0.w_dly_sig\[22\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2762 VGND tdc0.w_dly_sig\[109\] tdc0.w_dly_sig\[111\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2763 a_15255_9295# a_15035_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2764 a_17199_10357# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2765 VPWR a_2623_4373# a_2539_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2766 a_7005_9295# tdc0.w_dly_sig\[61\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2767 a_11251_8457# _026_ a_11333_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2768 tdc0.w_dly_sig_n\[75\] tdc0.w_dly_sig\[75\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2769 VPWR _056_ a_11974_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X2770 a_5805_13647# a_5639_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2771 tdc0.w_dly_sig\[34\] tdc0.w_dly_sig\[32\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2773 a_17213_8751# a_16679_8757# a_17118_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2774 VPWR a_2715_3035# a_2631_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2776 tdc0.w_dly_sig_n\[7\] tdc0.w_dly_sig_n\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2777 a_4053_9129# a_3063_8757# a_3927_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2778 a_14116_8207# a_13717_8207# a_13990_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2779 VGND a_17711_8725# a_17669_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2780 tdc0.w_dly_sig\[31\] tdc0.w_dly_sig_n\[30\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2781 a_7507_2223# a_6725_2229# a_7423_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2782 _049_ a_10239_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2783 VPWR net5 a_14287_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2784 a_7534_1109# a_7366_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2785 VPWR net1 tdc0.w_dly_sig_n\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2786 VGND a_8543_7093# _020_ VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=1 as=0.0991 ps=0.955 w=0.65 l=0.15
X2787 a_9206_14191# a_8767_14197# a_9121_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2788 a_14335_15975# a_14431_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2789 VPWR tdc0.w_dly_sig\[108\] tdc0.w_dly_sig_n\[108\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2790 _067_ a_6467_7369# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2791 tdc0.w_dly_sig\[84\] tdc0.w_dly_sig_n\[83\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2792 a_8083_4631# a_8374_4521# a_8325_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2794 _079_ a_9043_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2795 _014_ a_13735_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2796 a_9585_11043# _035_ a_9503_11043# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2797 a_4471_15279# a_3689_15285# a_4387_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2798 VPWR tdc0.w_dly_sig\[93\] tdc0.w_dly_sig\[95\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2799 a_14615_9269# a_14906_9569# a_14857_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2800 VGND tdc0.w_dly_sig\[60\] tdc0.w_dly_sig\[62\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2801 VPWR a_2623_17179# a_2539_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2802 tdc0.o_result\[92\] a_7867_4123# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2803 tdc0.w_dly_sig_n\[63\] tdc0.w_dly_sig\[63\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2804 tdc0.w_dly_sig\[97\] tdc0.w_dly_sig\[95\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2805 VPWR tdc0.w_dly_sig\[123\] tdc0.w_dly_sig_n\[123\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2806 VGND net4 a_13183_6583# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2807 a_6522_6549# a_6354_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2808 VGND a_9723_18365# a_9891_18267# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2809 uo_out[3] a_16332_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2811 VPWR tdc0.w_dly_sig_n\[38\] tdc0.w_dly_sig\[39\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2812 VGND a_2087_9839# a_2255_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2813 VGND tdc0.w_dly_sig\[89\] tdc0.w_dly_sig\[91\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2815 VGND tdc0.w_dly_sig\[107\] a_14533_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2816 a_2593_10633# tdc0.o_result\[75\] a_2511_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2817 VPWR tdc0.w_dly_sig_n\[104\] tdc0.w_dly_sig\[105\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2818 VGND a_16762_8207# clknet_4_11_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2819 VPWR tdc0.w_dly_sig_n\[100\] tdc0.w_dly_sig_n\[102\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2820 VPWR a_12999_591# net2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2821 a_6227_12925# a_5529_12559# a_5970_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2822 tdc0.w_dly_sig\[20\] tdc0.w_dly_sig_n\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2823 tdc0.w_dly_sig_n\[94\] tdc0.w_dly_sig\[94\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2824 VPWR tdc0.w_dly_sig_n\[22\] tdc0.w_dly_sig\[23\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2825 tdc0.w_dly_sig\[106\] tdc0.w_dly_sig\[104\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2826 VPWR a_3762_5461# a_3689_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2827 VPWR _072_ a_11869_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2828 VPWR a_9155_16341# a_9071_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2829 VGND tdc0.w_dly_sig_n\[106\] tdc0.w_dly_sig\[107\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2830 a_11023_12247# a_11119_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2831 VPWR tdc0.w_dly_sig\[128\] a_18121_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2832 VGND a_6119_4123# a_6077_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
R11 uio_out[3] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2833 tdc0.w_dly_sig\[8\] tdc0.w_dly_sig\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2834 a_8661_17455# tdc0.w_dly_sig\[18\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2835 a_7002_18365# a_6755_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2836 a_13947_6183# tdc0.o_result\[106\] a_14093_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2837 a_4421_1513# a_3431_1141# a_4295_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2838 a_11225_5487# _002_ a_11422_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2839 VPWR tdc0.w_dly_sig_n\[61\] tdc0.w_dly_sig_n\[63\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2840 a_16289_1679# a_15299_1679# a_16163_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2841 VGND a_17314_12559# clknet_4_14_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2842 a_16845_8757# a_16679_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2843 VGND _099_ a_6467_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X2844 a_5526_15101# a_5253_14735# a_5441_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2845 tdc0.w_dly_sig_n\[27\] tdc0.w_dly_sig\[27\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2846 tdc0.o_result\[35\] a_8051_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2847 VPWR tdc0.w_dly_sig\[99\] tdc0.w_dly_sig\[101\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2848 net1 a_18187_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2850 VGND clknet_4_7_0_clk a_8123_16373# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2851 tdc0.w_dly_sig_n\[86\] tdc0.w_dly_sig_n\[84\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2852 a_7883_7663# a_7019_7669# a_7626_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2854 _012_ a_12518_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X2855 VPWR clknet_4_1_0_clk a_6007_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2856 a_15106_9269# a_14906_9569# a_15255_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2857 VPWR a_16543_14887# tdc0.o_result\[124\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2858 VGND tdc0.w_dly_sig\[21\] tdc0.w_dly_sig_n\[21\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2859 tdc0.w_dly_sig\[48\] tdc0.w_dly_sig_n\[47\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2860 VPWR tdc0.w_dly_sig\[35\] tdc0.w_dly_sig_n\[35\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2861 a_8837_12393# a_7847_12021# a_8711_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2862 tdc0.w_dly_sig\[12\] tdc0.w_dly_sig\[10\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2863 a_5713_16911# a_5547_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2864 a_16600_12015# _071_ a_16332_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2865 a_13921_7779# _001_ a_13825_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2866 a_3348_13077# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2867 tdc0.w_dly_sig\[98\] tdc0.w_dly_sig\[96\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2868 clknet_4_3_0_clk a_7286_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2869 VGND a_14158_8319# a_14116_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2870 tdc0.w_dly_sig\[57\] tdc0.w_dly_sig_n\[56\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2871 tdc0.w_dly_sig\[114\] tdc0.w_dly_sig_n\[113\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2872 a_14449_1513# a_13459_1141# a_14323_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2873 VPWR tdc0.w_dly_sig\[67\] tdc0.w_dly_sig\[69\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2874 VGND a_9650_7637# _025_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2876 VGND a_1738_13077# a_1696_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2877 a_7277_9839# a_6743_9845# a_7182_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2878 a_10011_14887# a_10107_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2879 VGND a_4498_4373# a_4456_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2880 VGND _007_ a_8745_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2881 a_8933_14197# a_8767_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2882 VPWR clknet_0_clk a_3698_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2885 a_9263_16189# a_8565_15823# a_9006_15935# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2886 a_12591_12247# a_12875_12233# a_12810_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2887 tdc0.w_dly_sig_n\[52\] tdc0.w_dly_sig\[52\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2888 a_13599_14887# a_13695_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2890 a_13823_5193# net8 a_13605_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2891 clknet_4_7_0_clk a_7856_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X2892 a_13690_7895# _003_ a_13993_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X2893 a_1995_13103# a_1297_13109# a_1738_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2894 VGND clknet_4_0_0_clk a_3707_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2895 VGND tdc0.w_dly_sig_n\[121\] tdc0.w_dly_sig\[122\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2896 VPWR tdc0.w_dly_sig\[47\] tdc0.w_dly_sig_n\[47\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2897 VPWR a_15595_17429# a_15511_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2898 a_7755_12809# _070_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2899 a_13459_8751# _010_ a_13541_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2900 VGND a_15327_13799# _008_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2901 clknet_4_12_0_clk a_12548_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X2903 VGND a_2071_9563# a_2029_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2904 a_5169_9295# tdc0.o_result\[46\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2905 VPWR tdc0.o_result\[112\] a_16951_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2906 VGND net10 a_9227_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2907 a_18027_12233# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2908 a_14431_15797# a_14715_15797# a_14650_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2909 tdc0.w_dly_sig\[117\] tdc0.w_dly_sig\[115\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2910 _356_.X a_16732_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2911 a_14388_13621# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2912 VPWR a_14899_9269# a_14906_9569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2913 a_8412_12393# a_8013_12021# a_8286_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2914 VGND clknet_4_4_0_clk a_947_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2915 VGND a_14991_13321# a_14998_13225# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2916 a_7479_13103# net6 a_7561_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2917 tdc0.w_dly_sig\[14\] tdc0.w_dly_sig_n\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2918 VGND tdc0.w_dly_sig_n\[22\] tdc0.w_dly_sig_n\[24\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2919 a_11865_2767# a_11318_3041# a_11518_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2920 tdc0.w_dly_sig_n\[69\] tdc0.w_dly_sig\[69\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2921 tdc0.w_dly_sig_n\[47\] tdc0.w_dly_sig_n\[45\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2922 VPWR a_9631_14191# a_9799_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2923 tdc0.w_dly_sig\[8\] tdc0.w_dly_sig_n\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2924 a_17477_14735# a_16930_15009# a_17130_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2925 VPWR a_7987_4631# tdc0.o_result\[108\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2927 a_16849_1135# tdc0.w_dly_sig\[102\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2928 tdc0.w_dly_sig_n\[20\] tdc0.w_dly_sig_n\[18\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2929 a_5123_13103# a_4259_13109# a_4866_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2931 VGND tdc0.w_dly_sig\[23\] tdc0.w_dly_sig\[25\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2932 tdc0.o_result\[57\] a_6855_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2933 a_6755_17999# a_6619_17973# a_6335_17973# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2935 VGND tdc0.w_dly_sig_n\[1\] tdc0.w_dly_sig\[2\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2937 tdc0.w_dly_sig_n\[98\] tdc0.w_dly_sig\[98\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2938 a_11403_14409# clknet_4_12_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2939 VGND _015_ a_11873_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2941 VPWR tdc0.o_result\[1\] a_12200_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X2942 tdc0.w_dly_sig\[53\] tdc0.w_dly_sig\[51\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2943 a_18054_4765# a_17739_4631# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2944 a_5986_17277# a_5547_16911# a_5901_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2945 a_8859_6281# _020_ a_8941_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2946 a_5905_5487# tdc0.o_result\[83\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2947 VPWR a_7883_5487# a_8051_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2948 a_11023_14423# a_11119_14423# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2949 a_2122_1135# a_1683_1141# a_2037_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2950 VGND _012_ a_16381_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2951 VPWR a_9799_14165# a_9715_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2952 tdc0.o_result\[76\] a_2439_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2953 VGND tdc0.w_dly_sig\[59\] tdc0.w_dly_sig_n\[59\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2954 _078_ a_9319_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2955 tdc0.w_dly_sig\[43\] tdc0.w_dly_sig_n\[42\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2956 a_15453_9295# a_14899_9269# a_15106_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2957 _031_ a_9043_8457# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X2958 a_13165_3317# a_12999_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2959 VPWR a_18142_10116# a_18071_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2960 a_1393_11471# tdc0.w_dly_sig\[73\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2961 a_15588_14735# a_15189_14735# a_15462_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2962 VGND tdc0.w_dly_sig_n\[18\] tdc0.w_dly_sig\[19\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2963 tdc0.w_dly_sig_n\[79\] tdc0.w_dly_sig\[79\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2964 a_17102_1109# a_16934_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2965 a_4617_9071# tdc0.o_result\[49\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2966 VPWR a_11058_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2967 a_16155_18365# a_15373_17999# a_16071_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2968 a_16163_10749# a_15465_10383# a_15906_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2969 a_2750_14165# a_2582_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2970 a_1389_14735# a_1223_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2971 VGND net4 a_10446_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2972 _001_ a_13919_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2973 a_2398_3311# a_2125_3317# a_2313_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2974 tdc0.w_dly_sig_n\[92\] tdc0.w_dly_sig\[92\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2975 a_4237_10383# a_3247_10383# a_4111_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2976 a_9298_18365# a_9025_17999# a_9213_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2977 a_5951_15101# a_5253_14735# a_5694_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2978 VPWR tdc0.w_dly_sig\[43\] tdc0.w_dly_sig_n\[43\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2979 a_5345_4943# a_5179_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2980 tdc0.w_dly_sig\[36\] tdc0.w_dly_sig_n\[35\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2981 VPWR tdc0.w_dly_sig_n\[36\] tdc0.w_dly_sig_n\[38\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2982 VPWR tdc0.w_dly_sig\[30\] tdc0.w_dly_sig_n\[30\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2983 VGND tdc0.w_dly_sig\[112\] a_10393_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2984 clknet_4_11_0_clk a_16762_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2985 VPWR a_8178_8725# a_8105_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2986 a_6077_14735# a_5087_14735# a_5951_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2987 tdc0.w_dly_sig\[73\] tdc0.w_dly_sig\[71\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2988 tdc0.w_dly_sig_n\[121\] tdc0.w_dly_sig_n\[119\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2989 VGND tdc0.w_dly_sig_n\[82\] tdc0.w_dly_sig\[83\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2990 a_14786_9071# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2991 VGND tdc0.w_dly_sig_n\[63\] tdc0.w_dly_sig_n\[65\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2992 a_12692_8029# a_12649_7814# a_12620_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X2993 a_17935_10057# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2994 VGND a_12548_4917# clknet_4_8_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2995 VGND _007_ a_8745_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2996 tdc0.w_dly_sig\[49\] tdc0.w_dly_sig_n\[48\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2997 tdc0.w_dly_sig_n\[122\] tdc0.w_dly_sig\[122\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2998 a_6545_10927# tdc0.w_dly_sig\[60\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2999 VPWR tdc0.w_dly_sig_n\[46\] tdc0.w_dly_sig_n\[48\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3000 a_4011_8751# a_3229_8757# a_3927_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3001 VGND a_6246_13759# a_6204_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3002 VGND a_11711_591# net5 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3003 VGND net1 tdc0.w_dly_sig\[2\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3004 VGND tdc0.w_dly_sig_n\[0\] tdc0.w_dly_sig\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3005 tdc0.w_dly_sig\[10\] tdc0.w_dly_sig_n\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3006 VGND a_2547_5309# a_2715_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3007 tdc0.w_dly_sig_n\[57\] tdc0.w_dly_sig_n\[55\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3008 a_17746_9407# a_17578_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3009 a_4655_5309# a_3873_4943# a_4571_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3010 a_1205_11471# a_1039_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3011 tdc0.w_dly_sig_n\[126\] tdc0.w_dly_sig\[126\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3012 VPWR a_14195_7663# net11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3013 a_14526_2197# a_14358_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3014 tdc0.w_dly_sig\[45\] tdc0.w_dly_sig\[43\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3015 a_17746_9407# a_17578_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3016 VPWR a_7856_14165# clknet_4_7_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3017 VGND tdc0.o_result\[2\] a_14510_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3018 a_7274_4221# a_6835_3855# a_7189_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3019 a_1811_12015# a_947_12021# a_1554_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3020 tdc0.w_dly_sig_n\[60\] tdc0.w_dly_sig_n\[58\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3021 a_5802_12925# a_5363_12559# a_5717_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3022 tdc0.w_dly_sig_n\[110\] tdc0.w_dly_sig\[110\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3023 a_15427_15279# a_14563_15285# a_15170_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3024 a_4314_13759# a_4146_14013# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3025 tdc0.o_result\[117\] a_17711_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3026 VGND a_6963_4399# a_7131_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3027 a_2125_3317# a_1959_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3028 a_10217_3689# a_9227_3317# a_10091_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3029 VPWR tdc0.w_dly_sig_n\[81\] tdc0.w_dly_sig\[82\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3030 VPWR tdc0.w_dly_sig\[86\] tdc0.w_dly_sig_n\[86\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3031 VGND clknet_0_clk a_7286_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3033 a_1481_12015# a_947_12021# a_1386_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3034 a_7458_5487# a_7185_5493# a_7373_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3035 VGND a_14676_12809# uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3036 a_7561_13103# tdc0.o_result\[52\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3037 VPWR tdc0.w_dly_sig\[38\] tdc0.w_dly_sig_n\[38\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3038 a_14335_3855# a_14115_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3040 VPWR tdc0.w_dly_sig\[32\] tdc0.w_dly_sig_n\[32\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3041 a_15097_15279# a_14563_15285# a_15002_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3042 VGND tdc0.w_dly_sig\[5\] tdc0.w_dly_sig\[7\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3043 tdc0.o_result\[41\] a_7499_16091# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3044 tdc0.w_dly_sig_n\[91\] tdc0.w_dly_sig\[91\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3045 tdc0.w_dly_sig_n\[67\] tdc0.w_dly_sig_n\[65\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3046 a_10326_14735# a_10011_14887# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3047 VPWR a_4739_13915# a_4655_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3048 tdc0.w_dly_sig_n\[21\] tdc0.w_dly_sig_n\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3049 a_2248_1513# a_1849_1141# a_2122_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3050 a_5986_17277# a_5713_16911# a_5901_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3051 VGND _003_ _023_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3052 tdc0.w_dly_sig_n\[115\] tdc0.w_dly_sig_n\[113\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3053 VPWR a_14922_15797# a_14851_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3054 VPWR tdc0.w_dly_sig_n\[69\] tdc0.w_dly_sig_n\[71\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3055 VGND tdc0.w_dly_sig\[78\] tdc0.w_dly_sig_n\[78\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3056 a_14375_5193# _015_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3057 a_17719_8359# tdc0.o_result\[119\] a_17865_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3058 a_13735_9545# _013_ a_13817_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3059 VGND tdc0.w_dly_sig\[41\] tdc0.w_dly_sig_n\[41\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3060 a_8105_8751# a_7571_8757# a_8010_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3061 VGND tdc0.w_dly_sig\[100\] tdc0.w_dly_sig_n\[100\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3062 _069_ a_8399_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3063 a_2857_10383# tdc0.o_result\[51\] a_2511_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3064 _053_ a_10975_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3065 VGND a_8603_8725# a_8561_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3066 tdc0.w_dly_sig\[27\] tdc0.w_dly_sig_n\[26\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3067 _009_ _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3068 a_1389_14735# a_1223_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3069 tdc0.w_dly_sig_n\[112\] tdc0.w_dly_sig_n\[110\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3070 a_7001_6031# a_6835_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3071 a_12696_7119# a_12642_7271# a_12600_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.107 ps=0.98 w=0.65 l=0.15
X3072 a_13438_3311# a_12999_3317# a_13353_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3073 VGND _044_ a_11987_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X3074 a_5073_17999# tdc0.w_dly_sig\[20\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3075 tdc0.w_dly_sig_n\[22\] tdc0.w_dly_sig\[22\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3076 tdc0.w_dly_sig\[65\] tdc0.w_dly_sig\[63\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3077 _095_ a_14747_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3078 VPWR tdc0.w_dly_sig_n\[33\] tdc0.w_dly_sig\[34\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3079 a_1849_1141# a_1683_1141# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3080 a_18077_7663# a_17739_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3081 a_7607_3311# a_6743_3317# a_7350_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3082 tdc0.w_dly_sig_n\[86\] tdc0.w_dly_sig\[86\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3083 a_15906_10495# a_15738_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3084 a_18050_14468# a_17850_14313# a_18199_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3085 a_9217_5487# tdc0.o_result\[90\] a_9135_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3086 a_9723_18365# a_9025_17999# a_9466_18111# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3087 VGND a_7683_9563# a_7641_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3088 a_3781_18365# a_3247_17999# a_3686_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3089 VPWR tdc0.w_dly_sig\[96\] tdc0.w_dly_sig_n\[96\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3091 VPWR a_14519_9447# tdc0.o_result\[4\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3093 a_4245_4399# tdc0.w_dly_sig\[68\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3094 tdc0.o_result\[63\] a_8879_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3095 VGND tdc0.w_dly_sig\[37\] tdc0.w_dly_sig_n\[37\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3096 a_9397_1679# tdc0.w_dly_sig\[96\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3098 VGND tdc0.w_dly_sig_n\[87\] tdc0.w_dly_sig\[88\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3099 tdc0.o_result\[63\] a_8879_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3100 VPWR a_12631_591# net4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3101 a_11786_14191# a_11539_14569# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3102 tdc0.w_dly_sig\[15\] tdc0.w_dly_sig_n\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3103 a_17305_9295# a_17139_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3104 a_16332_9839# _101_ a_16166_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3105 VGND tdc0.w_dly_sig_n\[34\] tdc0.w_dly_sig_n\[36\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3106 a_11759_14557# a_11539_14569# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3107 VGND tdc0.w_dly_sig\[14\] tdc0.w_dly_sig\[16\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3108 tdc0.w_dly_sig_n\[53\] tdc0.w_dly_sig_n\[51\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3109 VPWR tdc0.w_dly_sig\[84\] tdc0.w_dly_sig\[86\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3110 VGND a_13599_14887# tdc0.o_result\[28\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3111 VPWR a_4755_2045# a_4923_1947# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3112 VGND a_8879_11989# a_8837_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3113 a_7400_3855# a_7001_3855# a_7274_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3114 VGND a_16331_1947# a_16289_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3115 a_17335_4943# a_17206_5217# a_16915_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3116 VPWR clknet_4_1_0_clk a_1407_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3117 VPWR a_1554_11989# a_1481_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3118 VPWR tdc0.w_dly_sig\[42\] tdc0.w_dly_sig_n\[42\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3119 a_18121_2767# a_17574_3041# a_17774_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3120 clknet_0_clk a_11058_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3121 tdc0.w_dly_sig\[7\] tdc0.w_dly_sig_n\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3122 VGND a_9374_14165# a_9332_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3123 a_9807_17687# tdc0.o_result\[45\] a_9953_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3124 a_4333_6581# a_4167_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3125 VGND a_14163_17973# a_14170_18273# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3126 VPWR _001_ a_9503_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X3127 a_3413_14735# a_3247_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3128 a_8500_4917# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3129 a_12210_9071# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3130 VGND a_16819_5095# tdc0.o_result\[113\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3131 a_6467_7369# net7 a_6549_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3132 VGND clknet_4_0_0_clk a_3891_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3133 _082_ a_9135_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3134 VGND tdc0.w_dly_sig_n\[72\] tdc0.w_dly_sig_n\[74\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3135 a_14186_3829# a_13986_4129# a_14335_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3136 VGND a_17406_10357# a_17335_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3137 VPWR a_4387_15279# a_4555_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3138 a_3321_5493# a_3155_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3139 VGND clknet_4_1_0_clk a_6007_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3140 a_15106_9269# a_14899_9269# a_15282_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3141 a_7737_8757# a_7571_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3142 a_2953_17455# a_2419_17461# a_2858_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3143 a_8730_16341# a_8562_16367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3144 tdc0.w_dly_sig\[27\] tdc0.w_dly_sig\[25\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3145 VGND a_4387_15279# a_4555_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3146 a_18383_12381# a_18163_12393# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3147 a_9043_8457# _024_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3148 a_9991_9661# a_9209_9295# a_9907_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3149 a_6522_6549# a_6354_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3150 a_10147_7369# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3151 a_3790_7119# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3152 a_10033_9295# a_9043_9295# a_9907_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3153 a_17567_2741# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3154 tdc0.w_dly_sig_n\[44\] tdc0.w_dly_sig\[44\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3155 clknet_4_8_0_clk a_12548_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X3156 a_8562_16367# a_8289_16373# a_8477_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3157 tdc0.o_result\[105\] a_12651_4123# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3158 VPWR a_6550_13103# clknet_4_6_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3159 tdc0.w_dly_sig_n\[23\] tdc0.w_dly_sig_n\[21\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3160 a_14868_8751# _005_ a_14952_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3161 clknet_4_14_0_clk a_17314_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3162 a_10945_14735# a_10398_15009# a_10598_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3163 _010_ a_12134_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3164 VPWR tdc0.w_dly_sig_n\[15\] tdc0.w_dly_sig\[16\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3165 a_9282_13077# a_9114_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3166 VGND tdc0.w_dly_sig_n\[79\] tdc0.w_dly_sig\[80\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3167 VPWR a_2566_3285# a_2493_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3168 tdc0.w_dly_sig\[46\] tdc0.w_dly_sig\[44\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3170 a_11119_12247# a_11410_12137# a_11361_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3171 a_14098_17999# a_13783_18151# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3172 VGND tdc0.w_dly_sig\[102\] tdc0.w_dly_sig_n\[102\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3173 VPWR a_11159_4943# _013_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3174 a_13564_3689# a_13165_3317# a_13438_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3175 VGND a_2547_1135# a_2715_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3176 VPWR _000_ a_9747_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0746 ps=0.775 w=0.42 l=0.15
X3177 a_15545_13481# a_14998_13225# a_15198_13380# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3178 tdc0.w_dly_sig\[102\] tdc0.w_dly_sig\[100\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3180 VPWR a_15630_14847# a_15557_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3181 _099_ a_8399_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3182 a_12326_11721# _005_ a_11504_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3183 a_9206_4221# a_8933_3855# a_9121_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3184 VGND tdc0.w_dly_sig\[19\] tdc0.w_dly_sig\[21\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3186 a_13898_1135# a_13625_1141# a_13813_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3187 a_9121_14191# tdc0.w_dly_sig\[30\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3188 VPWR tdc0.w_dly_sig\[37\] tdc0.w_dly_sig\[39\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3189 a_17314_17973# a_17114_18273# a_17463_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
D0 VGND _092_ sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X3190 VPWR a_3854_18111# a_3781_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3191 VPWR a_15198_13380# a_15127_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3192 VPWR tdc0.w_dly_sig_n\[73\] tdc0.w_dly_sig_n\[75\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3193 tdc0.w_dly_sig_n\[94\] tdc0.w_dly_sig_n\[92\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3194 VGND a_14335_15975# tdc0.o_result\[25\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3195 VPWR tdc0.w_dly_sig_n\[57\] tdc0.w_dly_sig\[58\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3196 tdc0.w_dly_sig\[35\] tdc0.w_dly_sig\[33\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3197 VGND _003_ _016_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3198 a_10195_4765# a_9975_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3199 a_11610_14468# a_11403_14409# a_11786_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3200 a_4387_15279# a_3523_15285# a_4130_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3201 VPWR tdc0.w_dly_sig_n\[116\] tdc0.w_dly_sig\[117\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3202 _087_ a_5639_6281# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3203 tdc0.w_dly_sig_n\[58\] tdc0.w_dly_sig_n\[56\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3204 VGND tdc0.w_dly_sig\[1\] tdc0.w_dly_sig\[3\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3205 a_18179_8983# tdc0.o_result\[117\] a_18325_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3206 VPWR _010_ a_5905_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3207 a_16915_4917# a_17206_5217# a_17157_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3208 VPWR tdc0.w_dly_sig\[46\] tdc0.w_dly_sig_n\[46\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3209 tdc0.w_dly_sig_n\[123\] tdc0.w_dly_sig\[123\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3210 a_8987_16367# a_8289_16373# a_8730_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3211 a_11539_14569# a_11403_14409# a_11119_14423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3212 a_4057_15279# a_3523_15285# a_3962_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3213 a_15282_9661# a_15035_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3214 _054_ a_10226_11247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3215 VGND tdc0.w_dly_sig_n\[120\] tdc0.w_dly_sig_n\[122\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3216 a_12530_17732# a_12330_17577# a_12679_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3217 tdc0.w_dly_sig_n\[47\] tdc0.w_dly_sig\[47\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3218 VGND a_12134_6549# _010_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3219 VPWR tdc0.w_dly_sig_n\[43\] tdc0.w_dly_sig_n\[45\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3220 net1 a_18187_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3221 a_15002_17455# a_14729_17461# a_14917_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3222 a_9401_12335# tdc0.o_result\[57\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3223 VGND net1 tdc0.w_dly_sig_n\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3224 VPWR a_18179_8983# _039_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X3225 a_2363_10927# a_1665_10933# a_2106_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3226 VGND a_9707_13077# a_9665_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3227 a_8399_8457# _029_ a_8481_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3228 VPWR a_7626_5461# a_7553_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3229 VGND tdc0.w_dly_sig\[16\] tdc0.w_dly_sig_n\[16\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3230 a_16412_6549# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3231 tdc0.w_dly_sig\[23\] tdc0.w_dly_sig_n\[22\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3232 a_14533_3855# a_13979_3829# a_14186_3829# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3233 a_18142_6852# a_17942_6697# a_18291_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3234 VPWR a_11023_12247# tdc0.o_result\[9\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3235 a_3413_14735# a_3247_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3236 VGND a_4279_18267# a_4237_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3237 VGND tdc0.w_dly_sig_n\[31\] tdc0.w_dly_sig\[32\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3238 a_2171_15101# a_1389_14735# a_2087_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3239 VGND a_2455_4399# a_2623_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3240 a_17774_16644# a_17574_16489# a_17923_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3241 tdc0.w_dly_sig\[83\] tdc0.w_dly_sig\[81\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3243 a_7699_6397# a_6835_6031# a_7442_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3244 a_2493_3311# a_1959_3317# a_2398_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3245 a_4755_4399# a_3891_4405# a_4498_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3246 a_4103_5487# a_3321_5493# a_4019_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3247 VPWR net28 a_11149_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3248 a_17525_17455# a_17187_17687# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3249 a_7791_1135# a_7093_1141# a_7534_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3250 a_16881_15101# a_16543_14887# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3251 VPWR tdc0.w_dly_sig_n\[83\] tdc0.w_dly_sig\[84\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3252 VGND a_4755_2045# a_4923_1947# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
D1 VGND _060_ sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X3253 VPWR tdc0.w_dly_sig_n\[30\] tdc0.w_dly_sig_n\[32\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3254 VGND tdc0.w_dly_sig\[24\] tdc0.w_dly_sig\[26\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3255 a_17567_2741# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3256 VGND clknet_4_9_0_clk a_12999_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3257 clknet_4_3_0_clk a_7286_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3258 a_13231_12381# a_13011_12393# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3259 tdc0.w_dly_sig_n\[10\] tdc0.w_dly_sig\[10\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3260 tdc0.w_dly_sig_n\[35\] tdc0.w_dly_sig\[35\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3261 tdc0.w_dly_sig_n\[51\] tdc0.w_dly_sig\[51\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3262 VPWR clknet_4_5_0_clk a_5547_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3263 a_3597_8751# a_3063_8757# a_3502_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3264 tdc0.w_dly_sig\[52\] tdc0.w_dly_sig_n\[51\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3265 VGND net2 a_11386_6652# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X3266 VPWR tdc0.w_dly_sig\[29\] a_14533_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3267 a_3781_10749# a_3247_10383# a_3686_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3268 VPWR a_12148_6005# a_11490_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=2.12 as=0.165 ps=1.33 w=1 l=0.15
X3269 a_16934_1135# a_16495_1141# a_16849_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3271 a_12292_8751# tdc0.o_result\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X3272 VGND tdc0.w_dly_sig_n\[107\] tdc0.w_dly_sig_n\[109\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3273 tdc0.w_dly_sig_n\[124\] tdc0.w_dly_sig_n\[122\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3274 a_6779_6575# a_6081_6581# a_6522_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3275 a_11061_11721# _054_ a_10965_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3276 a_7189_3855# tdc0.w_dly_sig\[93\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3277 a_4061_13647# tdc0.w_dly_sig\[53\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3279 tdc0.o_result\[10\] a_14031_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3280 VGND a_6027_7387# a_5985_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3281 a_14717_17999# a_14170_18273# a_14370_17973# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3283 VPWR tdc0.w_dly_sig_n\[79\] tdc0.w_dly_sig_n\[81\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3284 VPWR tdc0.w_dly_sig_n\[81\] tdc0.w_dly_sig_n\[83\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3285 VGND tdc0.w_dly_sig_n\[16\] tdc0.w_dly_sig\[17\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3286 VGND a_11058_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3287 VGND tdc0.w_dly_sig_n\[80\] tdc0.w_dly_sig_n\[82\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3288 tdc0.o_result\[96\] a_14951_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3289 a_18255_8041# a_18119_7881# a_17835_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3291 VPWR a_7775_3285# a_7691_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3292 tdc0.w_dly_sig_n\[39\] tdc0.w_dly_sig_n\[37\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3293 VPWR a_2014_6549# a_1941_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3294 tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3295 a_5249_13481# a_4259_13109# a_5123_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3296 a_12875_12233# clknet_4_12_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3297 a_18142_6852# a_17935_6793# a_18318_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3298 a_14783_2223# a_13919_2229# a_14526_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3299 VGND tdc0.w_dly_sig_n\[62\] tdc0.w_dly_sig_n\[64\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3300 VGND clknet_4_7_0_clk a_8767_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3301 VPWR a_1903_9661# a_2071_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3302 _019_ _000_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3303 VPWR clknet_4_5_0_clk a_4719_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3305 a_17102_1109# a_16934_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3306 a_9666_3311# a_9393_3317# a_9581_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3307 tdc0.w_dly_sig\[81\] tdc0.w_dly_sig_n\[80\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3308 tdc0.w_dly_sig\[87\] tdc0.w_dly_sig\[85\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3309 tdc0.w_dly_sig\[25\] tdc0.w_dly_sig_n\[24\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3310 tdc0.w_dly_sig\[45\] tdc0.w_dly_sig_n\[44\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3311 a_7553_5487# a_7019_5493# a_7458_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3312 a_8853_7119# _002_ a_8764_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0619 ps=0.715 w=0.42 l=0.15
X3314 tdc0.w_dly_sig\[99\] tdc0.w_dly_sig_n\[98\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3315 tdc0.o_result\[65\] a_7039_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3316 a_12642_7271# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3317 a_10033_1679# a_9043_1679# a_9907_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3318 tdc0.w_dly_sig_n\[83\] tdc0.w_dly_sig\[83\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3320 VGND a_7131_4373# a_7089_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3321 VPWR tdc0.w_dly_sig_n\[84\] tdc0.w_dly_sig_n\[86\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3322 VGND a_18142_6852# a_18071_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3323 tdc0.w_dly_sig\[61\] tdc0.w_dly_sig_n\[60\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3324 tdc0.w_dly_sig_n\[125\] tdc0.w_dly_sig\[125\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3325 VPWR a_14664_6005# clknet_4_9_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3326 a_6997_8207# a_6007_8207# a_6871_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3327 VPWR tdc0.w_dly_sig_n\[124\] tdc0.w_dly_sig\[125\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3328 VPWR a_2531_10901# a_2447_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3329 tdc0.w_dly_sig_n\[29\] tdc0.w_dly_sig\[29\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3330 a_11146_4719# net8 a_10977_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X3331 a_17835_7895# a_18119_7881# a_18054_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3332 a_10965_11721# _055_ a_10883_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X3333 VPWR clknet_4_1_0_clk a_3155_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3334 VPWR tdc0.w_dly_sig\[73\] tdc0.w_dly_sig_n\[73\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3335 VGND tdc0.w_dly_sig\[20\] tdc0.w_dly_sig_n\[20\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3336 a_8481_12809# tdc0.o_result\[56\] a_8399_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3337 tdc0.w_dly_sig\[55\] tdc0.w_dly_sig_n\[54\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3338 VGND net5 a_11067_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3339 VPWR clknet_4_5_0_clk a_1591_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3340 VPWR _010_ a_10137_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3342 VGND a_6395_1947# a_6353_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3343 tdc0.w_dly_sig_n\[69\] tdc0.w_dly_sig_n\[67\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3344 VGND a_18142_10116# a_18071_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3345 a_2122_3133# a_1849_2767# a_2037_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3346 a_17107_17973# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3347 VGND a_15427_4399# a_15595_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3348 VGND a_11403_14409# a_11410_14313# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3349 VGND clknet_0_clk a_4176_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3350 a_18121_16745# a_17574_16489# a_17774_16644# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3351 a_11251_8457# _026_ a_11333_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3352 VPWR tdc0.w_dly_sig_n\[37\] tdc0.w_dly_sig_n\[39\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3353 VGND tdc0.w_dly_sig_n\[11\] tdc0.w_dly_sig_n\[13\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3354 VPWR a_17555_10071# tdc0.o_result\[121\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3355 VPWR a_3854_10495# a_3781_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3356 VGND a_5951_4221# a_6119_4123# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3357 a_8289_16373# a_8123_16373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3358 a_9393_3317# a_9227_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
D2 VGND _038_ sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X3360 VGND a_10075_9563# a_10033_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3362 a_12644_8751# _046_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X3363 a_1937_12393# a_947_12021# a_1811_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3364 VPWR a_11872_7093# a_11214_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=2.12 as=0.165 ps=1.33 w=1 l=0.15
X3365 VPWR clknet_4_0_0_clk a_1959_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3366 a_5087_9545# _029_ a_5169_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3367 tdc0.w_dly_sig_n\[9\] tdc0.w_dly_sig_n\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3368 tdc0.w_dly_sig_n\[106\] tdc0.w_dly_sig\[106\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3369 VPWR a_9374_3967# a_9301_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3370 VGND tdc0.w_dly_sig\[127\] tdc0.w_dly_sig_n\[127\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3371 VGND tdc0.w_dly_sig_n\[3\] tdc0.w_dly_sig_n\[5\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3372 tdc0.w_dly_sig_n\[38\] tdc0.w_dly_sig_n\[36\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3373 VGND tdc0.w_dly_sig_n\[84\] tdc0.w_dly_sig\[85\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3376 a_5717_1679# tdc0.w_dly_sig\[88\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3379 a_17985_3311# a_17647_3543# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3380 tdc0.w_dly_sig\[28\] tdc0.w_dly_sig\[26\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3381 VPWR tdc0.w_dly_sig_n\[88\] tdc0.w_dly_sig_n\[90\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3382 tdc0.o_result\[105\] a_12651_4123# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3383 VPWR a_4571_14013# a_4739_13915# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3384 VGND a_17935_10057# a_17942_9961# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3385 VGND _039_ a_11435_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X3386 VGND a_4111_18365# a_4279_18267# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3387 a_17923_2767# a_17703_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3388 VPWR clknet_4_1_0_clk a_3063_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3389 VGND tdc0.w_dly_sig_n\[29\] tdc0.w_dly_sig_n\[31\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3391 a_9006_15935# a_8838_16189# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3392 tdc0.w_dly_sig_n\[48\] tdc0.w_dly_sig_n\[46\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3393 tdc0.w_dly_sig\[30\] tdc0.w_dly_sig_n\[29\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3395 VPWR tdc0.w_dly_sig\[72\] tdc0.w_dly_sig\[74\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3396 VGND tdc0.w_dly_sig\[66\] tdc0.w_dly_sig\[68\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3397 tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3398 _025_ a_9650_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X3400 a_15035_9295# a_14906_9569# a_14615_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3401 a_3007_14191# a_2143_14197# a_2750_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3402 a_11214_7093# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.175 ps=1.35 w=1 l=0.15
X3403 tdc0.w_dly_sig_n\[106\] tdc0.w_dly_sig_n\[104\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3404 a_15453_9295# a_14906_9569# a_15106_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3406 a_9577_9661# a_9043_9295# a_9482_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3407 tdc0.o_result\[58\] a_6947_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3408 a_9171_17455# a_8473_17461# a_8914_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3409 VGND tdc0.w_dly_sig\[12\] tdc0.w_dly_sig\[14\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3410 a_11797_8867# _074_ a_11701_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3411 VGND net9 a_11321_17775# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3412 a_4330_2045# a_4057_1679# a_4245_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3413 VGND a_14287_7119# _003_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3414 VGND a_14519_9447# tdc0.o_result\[4\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3415 VGND a_16578_13103# clknet_4_15_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X3416 a_11539_14569# a_11410_14313# a_11119_14423# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3417 VGND a_3762_5461# a_3720_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3418 VGND a_7286_7119# clknet_4_3_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3419 a_2677_14191# a_2143_14197# a_2582_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3420 a_1512_12393# a_1113_12021# a_1386_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3421 VGND tdc0.w_dly_sig\[114\] tdc0.w_dly_sig\[116\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3422 VGND clknet_4_4_0_clk a_3431_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3423 VPWR tdc0.w_dly_sig\[79\] tdc0.w_dly_sig\[81\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3424 a_17286_8725# a_17118_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3425 clknet_4_11_0_clk a_16762_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3426 _029_ a_11122_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3427 a_14729_17461# a_14563_17461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3428 VPWR a_17359_1135# a_17527_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3429 a_17359_1135# a_16661_1141# a_17102_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3430 tdc0.w_dly_sig\[50\] tdc0.w_dly_sig\[48\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3431 VGND a_1903_9661# a_2071_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3432 tdc0.w_dly_sig_n\[64\] tdc0.w_dly_sig_n\[62\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3433 tdc0.w_dly_sig_n\[78\] tdc0.w_dly_sig\[78\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3435 VGND clknet_4_3_0_clk a_7019_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3436 a_6503_14013# a_5639_13647# a_6246_13759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3437 VPWR a_7867_6299# a_7783_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3438 a_16547_7093# a_16838_7393# a_16789_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3439 a_5434_7485# a_5161_7119# a_5349_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3440 VPWR a_4923_4373# a_4839_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3441 a_8481_11721# tdc0.o_result\[59\] a_8399_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3442 tdc0.w_dly_sig\[46\] tdc0.w_dly_sig_n\[45\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3443 VGND _008_ a_14195_8867# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3444 tdc0.w_dly_sig_n\[70\] tdc0.w_dly_sig\[70\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3445 a_18163_12393# a_18034_12137# a_17743_12247# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3446 VGND tdc0.w_dly_sig_n\[96\] tdc0.w_dly_sig_n\[98\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3447 a_7442_6143# a_7274_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3448 tdc0.w_dly_sig\[38\] tdc0.w_dly_sig\[36\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3449 a_10122_8207# _002_ a_10026_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
R12 VPWR tt_um_hpretl_tt06_tdc_24.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3451 VPWR a_8367_4617# a_8374_4521# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3452 a_2685_12015# tdc0.o_result\[48\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3453 a_6173_14013# a_5639_13647# a_6078_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3454 a_15189_14735# a_15023_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3455 a_9301_4221# a_8767_3855# a_9206_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3456 VPWR tdc0.w_dly_sig_n\[85\] tdc0.w_dly_sig_n\[87\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3457 a_5526_4221# a_5253_3855# a_5441_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3458 VGND tdc0.w_dly_sig_n\[8\] tdc0.w_dly_sig_n\[10\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3459 VGND tdc0.w_dly_sig_n\[27\] tdc0.w_dly_sig_n\[29\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3460 a_3781_3317# a_3615_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3461 a_13993_1135# a_13459_1141# a_13898_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3462 VGND tdc0.w_dly_sig_n\[89\] tdc0.w_dly_sig_n\[91\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3463 uo_out[3] a_16332_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X3464 VGND tdc0.w_dly_sig_n\[101\] tdc0.w_dly_sig_n\[103\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3465 tdc0.w_dly_sig\[74\] tdc0.w_dly_sig\[72\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3466 tdc0.w_dly_sig_n\[41\] tdc0.w_dly_sig_n\[39\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3467 VGND a_9155_16341# a_9113_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3468 VPWR _002_ a_11987_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X3469 VPWR a_12318_7637# _015_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.331 pd=1.71 as=0.135 ps=1.27 w=1 l=0.15
X3470 a_9221_8457# _027_ a_9125_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3471 VPWR tdc0.w_dly_sig_n\[24\] tdc0.w_dly_sig_n\[26\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3472 VGND tdc0.w_dly_sig\[66\] tdc0.w_dly_sig_n\[66\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3473 a_1478_11837# a_1039_11471# a_1393_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3474 VGND clknet_4_5_0_clk a_2143_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3475 VPWR tdc0.o_result\[105\] a_13823_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3476 tdc0.w_dly_sig\[107\] tdc0.w_dly_sig\[105\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3477 tdc0.w_dly_sig\[113\] tdc0.w_dly_sig\[111\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R13 VGND uio_out[0] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3478 VGND a_10423_591# net3 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3479 tdc0.o_result\[37\] a_9431_16091# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3480 a_5694_14847# a_5526_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3481 a_1761_6575# tdc0.w_dly_sig\[77\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3482 clknet_4_9_0_clk a_14664_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3483 a_7470_17732# a_7270_17577# a_7619_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3484 VPWR a_14951_2197# a_14867_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3485 tdc0.w_dly_sig\[34\] tdc0.w_dly_sig_n\[33\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3486 tdc0.w_dly_sig\[112\] tdc0.w_dly_sig\[110\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3487 a_18129_9295# a_17139_9295# a_18003_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3488 tdc0.w_dly_sig\[53\] tdc0.w_dly_sig_n\[52\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3489 VGND tdc0.w_dly_sig\[115\] tdc0.w_dly_sig_n\[115\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3490 VGND a_13603_7093# net10 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3491 a_7090_9661# a_6651_9295# a_7005_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3492 VPWR a_16155_14423# _089_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X3493 a_17774_2741# a_17574_3041# a_17923_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3494 VPWR clknet_4_2_0_clk a_8399_1141# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3495 tdc0.o_result\[40\] a_6579_17179# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3496 VPWR a_9834_3285# a_9761_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3497 clknet_4_10_0_clk a_16412_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3498 VGND tdc0.w_dly_sig\[119\] tdc0.w_dly_sig_n\[119\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3499 VGND tdc0.w_dly_sig_n\[62\] tdc0.w_dly_sig\[63\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3500 VGND net11 a_15093_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3501 a_6835_12809# _090_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X3502 VGND tdc0.w_dly_sig_n\[18\] tdc0.w_dly_sig_n\[20\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3504 VPWR a_16163_2045# a_16331_1947# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3505 clknet_4_0_0_clk a_4176_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3506 VPWR a_8711_12015# a_8879_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3507 tdc0.w_dly_sig_n\[37\] tdc0.w_dly_sig\[37\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3508 a_17502_13647# a_17187_13799# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3510 a_11146_4719# tdc0.o_result\[86\] a_11060_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X3511 VGND a_18119_7881# a_18126_7785# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3512 VPWR tdc0.w_dly_sig\[103\] a_11865_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3513 a_14093_6031# _013_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X3514 tdc0.w_dly_sig_n\[36\] tdc0.w_dly_sig_n\[34\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3515 tdc0.w_dly_sig\[83\] tdc0.w_dly_sig_n\[82\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3516 tdc0.w_dly_sig_n\[77\] tdc0.w_dly_sig_n\[75\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3517 tdc0.w_dly_sig\[16\] tdc0.w_dly_sig\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3518 VGND tdc0.w_dly_sig\[10\] tdc0.w_dly_sig\[12\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3519 VGND tdc0.w_dly_sig_n\[97\] tdc0.w_dly_sig_n\[99\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3520 tdc0.w_dly_sig_n\[28\] tdc0.w_dly_sig_n\[26\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3521 tdc0.o_result\[103\] a_17803_1947# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3522 a_16543_14887# a_16639_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3523 VPWR tdc0.w_dly_sig\[17\] tdc0.w_dly_sig\[19\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3524 VPWR a_5859_7485# a_6027_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3525 tdc0.w_dly_sig_n\[42\] tdc0.w_dly_sig\[42\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3526 a_6883_17687# a_6979_17687# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3527 VGND tdc0.w_dly_sig_n\[8\] tdc0.w_dly_sig\[9\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3528 a_11539_13481# a_11410_13225# a_11119_13335# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3529 _015_ a_12318_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3530 VGND _009_ a_13805_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3531 VGND clknet_4_5_0_clk a_3247_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3532 VGND a_2623_4373# a_2581_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3533 a_12284_9545# _005_ a_12200_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3534 VGND tdc0.w_dly_sig\[117\] tdc0.w_dly_sig\[119\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3535 VGND a_10075_1947# a_10033_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3536 tdc0.w_dly_sig_n\[4\] tdc0.w_dly_sig_n\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3537 tdc0.w_dly_sig_n\[17\] tdc0.w_dly_sig\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3538 a_7185_5493# a_7019_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3539 VPWR a_9431_16091# a_9347_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3540 VPWR tdc0.w_dly_sig_n\[108\] tdc0.w_dly_sig\[109\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3541 a_2455_8751# a_1757_8757# a_2198_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3542 tdc0.w_dly_sig\[54\] tdc0.w_dly_sig_n\[53\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3543 a_15071_15823# a_14851_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3544 VPWR a_2290_2879# a_2217_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3545 VPWR a_6246_13759# a_6173_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3547 VGND tdc0.w_dly_sig_n\[125\] tdc0.w_dly_sig_n\[127\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3548 tdc0.w_dly_sig_n\[120\] tdc0.w_dly_sig\[120\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3549 tdc0.w_dly_sig_n\[50\] tdc0.w_dly_sig\[50\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3551 tdc0.w_dly_sig\[61\] tdc0.w_dly_sig\[59\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3552 a_16071_18365# a_15373_17999# a_15814_18111# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3554 a_14082_6575# a_13809_6581# a_13997_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3555 a_5031_6575# a_4333_6581# a_4774_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3556 a_13730_10205# a_13415_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3557 clknet_4_14_0_clk a_17314_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3558 VPWR tdc0.w_dly_sig\[124\] tdc0.w_dly_sig_n\[124\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3559 VPWR a_4498_1791# a_4425_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3560 a_12148_6005# _000_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.176 ps=1.68 w=0.42 l=0.15
X3561 tdc0.o_result\[3\] a_16331_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3562 a_4272_13647# a_3873_13647# a_4146_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3563 a_11745_6575# _003_ a_11649_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3564 a_13507_11293# a_13287_11305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3565 a_15189_14735# a_15023_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3567 VPWR tdc0.w_dly_sig\[39\] tdc0.w_dly_sig\[41\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3568 VPWR a_18326_7940# a_18255_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3569 VPWR a_16831_7093# a_16838_7393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3570 tdc0.w_dly_sig\[4\] tdc0.w_dly_sig\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3571 a_10505_5193# tdc0.o_result\[111\] a_10423_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3572 a_10147_16073# net6 a_10229_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3573 a_9481_5807# tdc0.o_result\[34\] a_9135_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3574 clknet_0_clk a_11058_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3575 VGND _012_ a_9941_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3576 VPWR ui_in[4] a_10423_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3577 VPWR clknet_4_9_0_clk a_13643_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3578 a_9761_3311# a_9227_3317# a_9666_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3579 uo_out[0] a_16332_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3580 a_11333_15599# tdc0.o_result\[41\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3581 VGND tdc0.w_dly_sig\[104\] tdc0.w_dly_sig_n\[104\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3582 a_11133_11721# _053_ a_11061_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3583 VPWR a_12007_1947# a_11923_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3584 a_8745_12559# tdc0.o_result\[120\] a_8399_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3585 VGND tdc0.w_dly_sig\[31\] tdc0.w_dly_sig\[33\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3586 VGND tdc0.w_dly_sig_n\[7\] tdc0.w_dly_sig\[8\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3587 VGND a_16762_8207# clknet_4_11_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3588 VGND net28 a_10585_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3589 tdc0.w_dly_sig\[39\] tdc0.w_dly_sig\[37\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3590 VPWR a_8527_10927# a_8695_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3591 a_11974_11721# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X3592 VPWR a_3698_12559# clknet_4_4_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3593 VPWR _003_ a_9485_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X3594 a_7216_9295# a_6817_9295# a_7090_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3595 tdc0.w_dly_sig\[42\] tdc0.w_dly_sig_n\[41\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3596 a_2455_8751# a_1591_8757# a_2198_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3597 a_5158_18365# a_4719_17999# a_5073_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3598 tdc0.w_dly_sig\[82\] tdc0.w_dly_sig\[80\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3601 a_7856_14165# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3602 clknet_0_clk a_11058_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3603 VPWR a_3790_7119# clknet_4_1_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3604 tdc0.w_dly_sig\[3\] tdc0.w_dly_sig\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3605 a_9681_11043# _034_ a_9585_11043# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3606 a_6273_17455# tdc0.o_result\[42\] a_6191_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3607 VPWR tdc0.w_dly_sig_n\[107\] tdc0.w_dly_sig\[108\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3608 clknet_0_clk a_11058_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3610 tdc0.o_result\[74\] a_1979_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3611 a_12548_14165# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3612 tdc0.w_dly_sig_n\[87\] tdc0.w_dly_sig\[87\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3613 tdc0.w_dly_sig_n\[46\] tdc0.w_dly_sig\[46\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3614 _055_ a_10423_5193# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3615 VGND tdc0.w_dly_sig_n\[118\] tdc0.w_dly_sig\[119\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3616 _022_ a_11214_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3617 tdc0.o_result\[74\] a_1979_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3618 VGND a_16332_12015# uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3619 clknet_4_6_0_clk a_6550_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3620 VGND a_7775_3285# a_7733_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3621 VGND a_16181_5461# _084_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3622 tdc0.w_dly_sig\[64\] tdc0.w_dly_sig_n\[63\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3623 VPWR a_10046_4676# a_9975_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3624 tdc0.w_dly_sig_n\[122\] tdc0.w_dly_sig_n\[120\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3625 VPWR clknet_4_2_0_clk a_9043_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3626 a_16394_12533# a_16194_12833# a_16543_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3627 a_14370_17973# a_14170_18273# a_14519_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3628 tdc0.w_dly_sig\[15\] tdc0.w_dly_sig\[13\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3629 tdc0.w_dly_sig\[24\] tdc0.w_dly_sig\[22\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3630 tdc0.w_dly_sig_n\[45\] tdc0.w_dly_sig_n\[43\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3631 tdc0.o_result\[76\] a_2439_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3632 a_13109_10927# a_12771_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3634 a_6537_16911# a_5547_16911# a_6411_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3635 a_12284_9545# _081_ a_12552_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3636 VGND a_10759_8181# _005_ VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X3637 VPWR a_6239_18151# tdc0.o_result\[18\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3638 tdc0.w_dly_sig\[108\] tdc0.w_dly_sig\[106\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3639 a_4425_2045# a_3891_1679# a_4330_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3640 a_9941_11471# tdc0.o_result\[29\] a_9595_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3641 tdc0.w_dly_sig\[112\] tdc0.w_dly_sig_n\[111\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3642 tdc0.w_dly_sig\[88\] tdc0.w_dly_sig_n\[87\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3643 a_15738_10749# a_15465_10383# a_15653_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3644 tdc0.w_dly_sig_n\[108\] tdc0.w_dly_sig_n\[106\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3645 a_3509_5487# tdc0.w_dly_sig\[72\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3646 a_9043_6575# _026_ a_9125_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3647 VPWR clknet_4_5_0_clk a_3247_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3648 VPWR a_5602_7231# a_5529_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3649 a_2087_15101# a_1223_14735# a_1830_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3650 VPWR a_15170_4373# a_15097_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3651 VGND a_15595_4373# a_15553_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3652 VPWR clknet_4_2_0_clk a_9227_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3653 VPWR clknet_4_3_0_clk a_6835_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3654 tdc0.w_dly_sig_n\[71\] tdc0.w_dly_sig\[71\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3655 a_9025_17999# a_8859_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3656 VGND a_16163_2045# a_16331_1947# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3657 tdc0.w_dly_sig\[125\] tdc0.w_dly_sig_n\[124\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3658 a_17543_8751# a_16845_8757# a_17286_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3659 VGND tdc0.w_dly_sig\[122\] tdc0.w_dly_sig_n\[122\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3660 a_17555_6807# a_17651_6807# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3661 tdc0.w_dly_sig_n\[14\] tdc0.w_dly_sig\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3662 tdc0.w_dly_sig_n\[76\] tdc0.w_dly_sig_n\[74\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3663 VPWR a_5694_3967# a_5621_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3664 a_5529_7485# a_4995_7119# a_5434_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3665 tdc0.w_dly_sig_n\[52\] tdc0.w_dly_sig_n\[50\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3666 a_3026_17429# a_2858_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3667 a_10391_14709# clknet_4_12_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3668 VPWR a_11943_17687# tdc0.o_result\[20\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3669 tdc0.w_dly_sig\[109\] tdc0.w_dly_sig\[107\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3670 tdc0.o_result\[103\] a_17803_1947# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R14 uio_oe[6] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3672 VGND tdc0.w_dly_sig\[8\] tdc0.w_dly_sig\[10\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3673 VPWR a_3348_13077# clknet_4_5_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3675 tdc0.w_dly_sig_n\[37\] tdc0.w_dly_sig_n\[35\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3676 VGND tdc0.w_dly_sig_n\[89\] tdc0.w_dly_sig\[90\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3677 a_6043_5309# a_5179_4943# a_5786_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3678 VPWR tdc0.w_dly_sig_n\[27\] tdc0.w_dly_sig\[28\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3679 a_15269_15823# a_14722_16097# a_14922_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3681 a_3969_3311# tdc0.w_dly_sig\[84\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3682 a_6112_16911# a_5713_16911# a_5986_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3683 tdc0.w_dly_sig_n\[30\] tdc0.w_dly_sig\[30\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3684 VPWR tdc0.w_dly_sig_n\[123\] tdc0.w_dly_sig_n\[125\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3685 _090_ a_3247_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X3686 VGND tdc0.w_dly_sig_n\[70\] tdc0.w_dly_sig_n\[72\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3688 VGND net10 a_6537_17775# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3689 VGND tdc0.w_dly_sig\[92\] tdc0.w_dly_sig\[94\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3690 a_13625_1141# a_13459_1141# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3691 clknet_4_8_0_clk a_12548_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3692 VGND a_7258_9407# a_7216_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3693 a_8745_11471# tdc0.o_result\[123\] a_8399_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3694 a_8481_6575# tdc0.o_result\[91\] a_8399_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3695 VGND a_12875_12233# a_12882_12137# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3696 tdc0.w_dly_sig_n\[8\] tdc0.w_dly_sig_n\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3697 tdc0.w_dly_sig_n\[45\] tdc0.w_dly_sig\[45\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3698 VPWR tdc0.w_dly_sig\[25\] tdc0.w_dly_sig_n\[25\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3699 VGND a_13599_4007# tdc0.o_result\[106\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3700 tdc0.w_dly_sig\[97\] tdc0.w_dly_sig_n\[96\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3701 a_9991_2045# a_9209_1679# a_9907_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3702 net2 a_12999_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X3703 tdc0.w_dly_sig_n\[102\] tdc0.w_dly_sig\[102\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3704 a_6453_4399# tdc0.w_dly_sig\[89\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3705 a_13511_10071# a_13802_9961# a_13753_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3706 a_1485_13103# tdc0.w_dly_sig\[51\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3707 a_2217_5309# a_1683_4943# a_2122_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3708 tdc0.o_result\[33\] a_8603_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3709 VGND tdc0.w_dly_sig_n\[128\] tdc0.w_dly_sig\[129\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3710 a_14157_4917# net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X3711 a_8941_6281# tdc0.o_result\[68\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3712 a_15170_17429# a_15002_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3713 VPWR a_18119_4617# a_18126_4521# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3714 tdc0.w_dly_sig_n\[89\] tdc0.w_dly_sig\[89\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3715 a_7366_1135# a_6927_1141# a_7281_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3716 a_17543_8751# a_16679_8757# a_17286_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3717 a_4222_3285# a_4054_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3718 VPWR tdc0.w_dly_sig\[21\] tdc0.w_dly_sig\[23\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3719 a_8102_10927# a_7829_10933# a_8017_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3720 VPWR a_9723_18365# a_9891_18267# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3721 tdc0.o_result\[45\] a_3451_17429# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3722 VPWR tdc0.w_dly_sig_n\[90\] tdc0.w_dly_sig\[91\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3723 VGND _069_ a_7755_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X3724 a_15381_5487# _015_ a_15235_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X3725 VGND a_17314_17973# a_17243_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3726 VPWR _052_ a_11133_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3727 tdc0.o_result\[45\] a_3451_17429# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3728 a_15162_5095# _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X3730 a_7097_9839# tdc0.w_dly_sig\[63\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3731 VPWR tdc0.w_dly_sig\[102\] tdc0.w_dly_sig\[104\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3732 VPWR a_6227_2045# a_6395_1947# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3733 VGND clknet_4_3_0_clk a_9043_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3734 VGND a_17803_1947# a_17761_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3736 a_10177_7983# _003_ a_10093_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.0878 ps=0.92 w=0.65 l=0.15
X3737 VPWR a_11058_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3738 _046_ a_11987_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X3739 VPWR tdc0.w_dly_sig\[65\] tdc0.w_dly_sig\[67\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3740 VPWR a_5031_17455# a_5199_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3741 VGND tdc0.w_dly_sig\[125\] tdc0.w_dly_sig\[127\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3742 tdc0.w_dly_sig_n\[32\] tdc0.w_dly_sig\[32\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3743 a_5621_4221# a_5087_3855# a_5526_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3744 a_4479_3311# a_3781_3317# a_4222_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3745 VPWR clknet_0_clk a_8500_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3746 a_10011_14887# a_10107_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3747 tdc0.w_dly_sig_n\[20\] tdc0.w_dly_sig\[20\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3748 a_4195_18365# a_3413_17999# a_4111_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3750 a_9213_17999# tdc0.w_dly_sig\[22\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3751 _010_ a_12134_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X3752 VPWR a_14250_6549# a_14177_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3753 a_6430_11989# a_6262_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3754 _091_ a_6835_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X3755 VPWR a_16451_7271# tdc0.o_result\[115\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3756 VPWR tdc0.w_dly_sig\[6\] tdc0.w_dly_sig_n\[6\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3757 VGND tdc0.w_dly_sig\[123\] tdc0.w_dly_sig\[125\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3758 VPWR a_9907_9661# a_10075_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3760 _033_ a_9595_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3761 a_13817_9545# tdc0.o_result\[60\] a_13735_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3762 tdc0.w_dly_sig_n\[48\] tdc0.w_dly_sig\[48\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3763 VPWR a_13599_4007# tdc0.o_result\[106\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3764 VGND a_12548_4917# clknet_4_8_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3766 a_9389_15823# a_8399_15823# a_9263_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3767 VPWR tdc0.w_dly_sig\[4\] tdc0.w_dly_sig_n\[4\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3768 a_10391_14709# clknet_4_12_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3769 a_13947_3311# a_13165_3317# a_13863_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3770 VGND a_18171_9563# a_18129_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3771 _037_ a_10239_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3772 VPWR clknet_4_14_0_clk a_15299_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3773 a_13603_7093# _009_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X3774 a_5851_13335# tdc0.o_result\[54\] a_5997_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X3775 tdc0.w_dly_sig\[38\] tdc0.w_dly_sig_n\[37\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3776 tdc0.w_dly_sig_n\[44\] tdc0.w_dly_sig_n\[42\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3777 tdc0.w_dly_sig\[91\] tdc0.w_dly_sig_n\[90\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3778 tdc0.w_dly_sig\[94\] tdc0.w_dly_sig_n\[93\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3779 a_3367_17455# a_2585_17461# a_3283_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3780 VGND clknet_0_clk a_16412_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3781 a_18071_6953# a_17942_6697# a_17651_6807# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3782 VGND _002_ _016_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3783 VPWR tdc0.w_dly_sig\[98\] tdc0.w_dly_sig\[100\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3784 a_17038_7093# a_16831_7093# a_17214_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3785 tdc0.w_dly_sig_n\[61\] tdc0.w_dly_sig_n\[59\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3786 VPWR tdc0.w_dly_sig_n\[38\] tdc0.w_dly_sig_n\[40\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3787 a_4019_5487# a_3155_5493# a_3762_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3788 VPWR tdc0.w_dly_sig_n\[95\] tdc0.w_dly_sig_n\[97\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3789 VPWR tdc0.w_dly_sig_n\[98\] tdc0.w_dly_sig\[99\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3790 a_13905_8207# tdc0.w_dly_sig\[12\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3791 VGND tdc0.w_dly_sig\[14\] a_11957_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3792 _072_ a_11251_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3793 VPWR a_2623_8725# a_2539_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3794 a_14186_3829# a_13979_3829# a_14362_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3795 tdc0.w_dly_sig_n\[26\] tdc0.w_dly_sig_n\[24\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3796 VPWR a_17935_10057# a_17942_9961# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3798 a_14407_1135# a_13625_1141# a_14323_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3800 a_7492_1513# a_7093_1141# a_7366_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3801 VGND a_11027_6005# net7 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3802 VGND tdc0.o_result\[109\] a_9965_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3803 a_4111_15101# a_3247_14735# a_3854_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3804 VPWR a_17774_17732# a_17703_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3805 clknet_4_2_0_clk a_8500_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3806 VPWR tdc0.w_dly_sig\[79\] tdc0.w_dly_sig_n\[79\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3807 VGND a_16578_13103# clknet_4_15_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3808 a_2547_3133# a_1849_2767# a_2290_2879# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3809 a_4793_13103# a_4259_13109# a_4698_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3810 VPWR tdc0.w_dly_sig\[44\] tdc0.w_dly_sig\[46\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3811 VGND a_14951_2197# a_14909_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3812 _043_ a_11067_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X3813 a_5901_16911# tdc0.w_dly_sig\[41\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3814 VGND tdc0.w_dly_sig_n\[15\] tdc0.w_dly_sig_n\[17\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3815 VPWR tdc0.w_dly_sig\[120\] tdc0.w_dly_sig\[122\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3816 a_3007_14191# a_2309_14197# a_2750_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3817 a_16732_11445# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3819 a_3854_14847# a_3686_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3820 a_16289_10383# a_15299_10383# a_16163_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3821 VPWR tdc0.w_dly_sig_n\[75\] tdc0.w_dly_sig_n\[77\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3822 a_15761_13647# _007_ a_15327_13799# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3823 a_5721_6281# tdc0.o_result\[82\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3824 VGND a_16831_7093# a_16838_7393# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3825 a_11974_11721# _061_ a_11504_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3826 tdc0.w_dly_sig\[19\] tdc0.w_dly_sig\[17\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3827 VPWR tdc0.w_dly_sig_n\[118\] tdc0.w_dly_sig_n\[120\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3828 a_17567_13621# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3830 VPWR clknet_4_0_0_clk a_3431_1141# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3831 tdc0.w_dly_sig\[118\] tdc0.w_dly_sig_n\[117\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3833 uo_out[1] a_12284_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3834 VGND a_13690_7895# _004_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X3835 a_9493_2223# tdc0.o_result\[93\] a_9411_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3836 VGND tdc0.w_dly_sig\[111\] a_18121_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3837 a_10241_17775# _029_ a_9807_17687# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3838 VGND _028_ a_8745_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3839 VPWR a_16578_13103# clknet_4_15_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3840 VGND tdc0.w_dly_sig\[106\] tdc0.w_dly_sig_n\[106\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3841 tdc0.o_result\[97\] a_12007_1947# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3842 a_17214_7485# a_16967_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3843 a_3870_10927# a_3431_10933# a_3785_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3844 _096_ a_16127_7779# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X3845 VPWR a_7791_1135# a_7959_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3846 a_1665_10933# a_1499_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3847 tdc0.w_dly_sig_n\[10\] tdc0.w_dly_sig_n\[8\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3848 a_6550_13103# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3849 tdc0.w_dly_sig_n\[29\] tdc0.w_dly_sig_n\[27\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3850 VPWR _047_ a_13341_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3851 a_6717_10633# _098_ a_6645_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3853 VGND a_6227_2045# a_6395_1947# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3854 VGND a_3670_8725# a_3628_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3855 a_7783_4221# a_7001_3855# a_7699_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3856 net8 a_12171_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X3857 net5 a_11711_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X3858 VPWR a_6211_5211# a_6127_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3859 VPWR tdc0.w_dly_sig_n\[122\] tdc0.w_dly_sig\[123\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3860 a_14362_4221# a_14115_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3862 a_14510_12559# _091_ a_14676_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3863 VGND tdc0.w_dly_sig_n\[77\] tdc0.w_dly_sig_n\[79\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3864 clknet_4_10_0_clk a_16412_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3865 tdc0.w_dly_sig\[41\] tdc0.w_dly_sig\[39\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3866 uo_out[4] a_14952_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3867 a_3812_10383# a_3413_10383# a_3686_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3868 VPWR tdc0.w_dly_sig\[2\] a_17753_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3869 VPWR a_12548_14165# clknet_4_12_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3870 tdc0.w_dly_sig\[113\] tdc0.w_dly_sig_n\[112\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3871 VGND a_9907_9661# a_10075_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3872 VGND tdc0.w_dly_sig\[10\] a_11957_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3873 tdc0.w_dly_sig_n\[35\] tdc0.w_dly_sig_n\[33\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3875 VGND tdc0.w_dly_sig\[27\] tdc0.w_dly_sig\[29\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3876 VPWR tdc0.w_dly_sig\[91\] tdc0.w_dly_sig_n\[91\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3878 VGND clknet_4_2_0_clk a_9043_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3880 a_10226_11247# _016_ a_10057_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X3881 VPWR a_4866_13077# a_4793_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3882 VPWR a_6411_17277# a_6579_17179# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3883 tdc0.w_dly_sig_n\[65\] tdc0.w_dly_sig_n\[63\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3884 VPWR a_17711_8725# a_17627_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3885 a_9366_10071# _080_ a_9669_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X3886 a_1945_4399# tdc0.w_dly_sig\[79\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3887 a_14645_5807# tdc0.o_result\[96\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3888 a_9753_11043# _033_ a_9681_11043# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3889 a_4057_1679# a_3891_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3890 a_10226_11247# tdc0.o_result\[55\] a_10140_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X3891 a_4195_10749# a_3413_10383# a_4111_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3892 VPWR tdc0.w_dly_sig\[68\] tdc0.w_dly_sig\[70\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3893 tdc0.w_dly_sig_n\[6\] tdc0.w_dly_sig_n\[4\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3894 tdc0.w_dly_sig\[85\] tdc0.w_dly_sig\[83\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R15 uio_out[7] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3896 VGND tdc0.w_dly_sig_n\[124\] tdc0.w_dly_sig_n\[126\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3897 tdc0.o_result\[71\] a_4187_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3898 VPWR a_9907_2045# a_10075_1947# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3899 VGND tdc0.w_dly_sig\[57\] tdc0.w_dly_sig_n\[57\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3900 VGND a_11058_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3901 tdc0.w_dly_sig\[68\] tdc0.w_dly_sig\[66\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3902 a_10975_8751# net7 a_11057_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3903 VGND _012_ a_9757_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3904 VPWR a_6883_17687# tdc0.o_result\[16\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3905 a_16732_11445# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3906 tdc0.w_dly_sig\[9\] tdc0.w_dly_sig_n\[8\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3907 VGND clknet_0_clk a_6550_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3908 a_1849_4943# a_1683_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3909 a_7837_12809# _070_ a_7755_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X3910 tdc0.w_dly_sig_n\[100\] tdc0.w_dly_sig\[100\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3911 tdc0.w_dly_sig_n\[115\] tdc0.w_dly_sig\[115\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3912 VPWR tdc0.o_result\[114\] a_16399_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3913 tdc0.w_dly_sig_n\[62\] tdc0.w_dly_sig_n\[60\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3914 VGND a_12376_8751# uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3916 a_8435_8751# a_7737_8757# a_8178_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3917 a_17314_12559# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3918 VPWR _001_ a_9485_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.143 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3919 a_11692_7119# net4 a_11596_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.107 ps=0.98 w=0.65 l=0.15
X3921 a_9677_5193# _020_ a_9531_5095# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X3922 VPWR _019_ a_8941_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3923 a_4498_1791# a_4330_2045# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3924 VGND tdc0.w_dly_sig\[74\] tdc0.w_dly_sig\[76\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3925 a_5717_12559# tdc0.w_dly_sig\[57\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3926 a_7875_1135# a_7093_1141# a_7791_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3928 VPWR tdc0.w_dly_sig\[58\] tdc0.w_dly_sig\[60\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3929 tdc0.w_dly_sig_n\[124\] tdc0.w_dly_sig\[124\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3930 a_15553_17833# a_14563_17461# a_15427_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3931 tdc0.w_dly_sig_n\[32\] tdc0.w_dly_sig_n\[30\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3932 a_17774_13621# a_17574_13921# a_17923_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3933 VPWR a_17739_7895# tdc0.o_result\[118\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3934 a_7599_9661# a_6817_9295# a_7515_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3935 clknet_4_12_0_clk a_12548_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3936 a_9577_2045# a_9043_1679# a_9482_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3937 tdc0.w_dly_sig\[80\] tdc0.w_dly_sig\[78\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3938 a_13993_7779# _002_ a_13921_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3940 a_9849_17999# a_8859_17999# a_9723_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3941 VPWR a_13599_14887# tdc0.o_result\[28\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3942 VPWR a_2455_17277# a_2623_17179# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3943 a_18121_16745# a_17567_16585# a_17774_16644# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3944 VGND tdc0.w_dly_sig_n\[111\] tdc0.w_dly_sig_n\[113\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3945 VPWR tdc0.w_dly_sig_n\[5\] tdc0.w_dly_sig\[6\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3947 tdc0.o_result\[69\] a_4739_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3948 tdc0.w_dly_sig_n\[98\] tdc0.w_dly_sig_n\[96\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3950 VGND _032_ a_9503_11043# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3951 VPWR tdc0.w_dly_sig_n\[74\] tdc0.w_dly_sig_n\[76\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3952 VGND a_8527_10927# a_8695_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3953 net4 a_12631_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X3954 VGND _007_ a_11597_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3955 a_14715_15797# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3956 a_10026_8207# _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.175 ps=1.26 w=0.42 l=0.15
X3957 VGND tdc0.w_dly_sig_n\[78\] tdc0.w_dly_sig_n\[80\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3958 VPWR a_3698_12559# clknet_4_4_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3959 a_2309_14197# a_2143_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3960 a_4571_5309# a_3873_4943# a_4314_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3961 tdc0.w_dly_sig_n\[91\] tdc0.w_dly_sig_n\[89\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3962 a_2030_8751# a_1591_8757# a_1945_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3963 clknet_4_7_0_clk a_7856_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3964 VGND tdc0.w_dly_sig_n\[101\] tdc0.w_dly_sig\[102\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3965 a_14541_8207# a_13551_8207# a_14415_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3966 VGND clknet_0_clk a_3790_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3967 _059_ a_10791_16073# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3968 clknet_0_clk a_11058_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3969 VPWR tdc0.w_dly_sig\[5\] a_15453_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3970 tdc0.o_result\[49\] a_3175_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3971 a_8435_8751# a_7571_8757# a_8178_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3973 uo_out[5] a_11456_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3975 VPWR tdc0.w_dly_sig\[3\] tdc0.w_dly_sig\[5\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3976 a_14673_16189# a_14335_15975# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3977 clknet_4_12_0_clk a_12548_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3978 tdc0.o_result\[97\] a_12007_1947# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3979 VGND net5 a_12783_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X3981 _056_ a_10883_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X3982 clknet_4_6_0_clk a_6550_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3983 VPWR tdc0.w_dly_sig_n\[17\] tdc0.w_dly_sig\[18\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3984 VPWR a_1811_12015# a_1979_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3985 VGND a_4739_13915# a_4697_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3986 a_17870_6941# a_17555_6807# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3987 VPWR a_14031_3285# a_13947_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3988 VPWR tdc0.w_dly_sig\[120\] tdc0.w_dly_sig_n\[120\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3989 tdc0.w_dly_sig_n\[12\] tdc0.w_dly_sig_n\[10\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3990 uo_out[0] a_16332_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3991 a_9424_17999# a_9025_17999# a_9298_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3992 a_16301_17455# net9 a_16155_17687# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X3993 a_12801_2223# tdc0.w_dly_sig\[99\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3994 a_16022_7119# tdc0.o_result\[115\] a_15936_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X3996 VGND tdc0.w_dly_sig_n\[65\] tdc0.w_dly_sig\[66\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3997 a_14335_15975# a_14431_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3998 a_8745_6895# tdc0.o_result\[35\] a_8399_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3999 a_11321_9071# tdc0.o_result\[9\] a_10975_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4000 tdc0.o_result\[12\] a_14675_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4001 VPWR tdc0.w_dly_sig_n\[20\] tdc0.w_dly_sig_n\[22\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4002 a_11973_3855# tdc0.w_dly_sig\[106\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4003 clknet_4_3_0_clk a_7286_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4004 a_8795_12015# a_8013_12021# a_8711_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4005 VPWR a_9485_7485# _028_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X4006 a_18119_4617# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4007 tdc0.w_dly_sig_n\[54\] tdc0.w_dly_sig_n\[52\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4008 VGND a_10598_14709# a_10527_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4009 VGND _014_ a_14195_8867# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X4010 VGND a_11456_10927# uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4011 VGND a_4463_10901# a_4421_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4012 a_10321_10633# tdc0.o_result\[77\] a_10239_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4013 tdc0.o_result\[81\] a_2715_3035# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4014 tdc0.w_dly_sig_n\[74\] tdc0.w_dly_sig_n\[72\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4015 a_14533_14735# a_13986_15009# a_14186_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4016 a_4222_3285# a_4054_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4017 a_17703_2767# a_17574_3041# a_17283_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4018 tdc0.w_dly_sig_n\[63\] tdc0.w_dly_sig_n\[61\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4019 a_1662_9839# a_1389_9845# a_1577_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4020 VGND clknet_4_4_0_clk a_1039_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4021 net3 a_10423_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4024 VPWR _010_ a_6549_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4025 VGND tdc0.o_result\[26\] a_16589_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4027 VPWR clknet_0_clk a_16762_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4028 VGND tdc0.w_dly_sig\[112\] tdc0.w_dly_sig\[114\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4030 a_9650_9407# a_9482_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4032 a_17385_7119# a_16838_7393# a_17038_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4033 tdc0.w_dly_sig_n\[33\] tdc0.w_dly_sig\[33\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4034 VPWR tdc0.w_dly_sig\[82\] tdc0.w_dly_sig_n\[82\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4035 tdc0.w_dly_sig\[62\] tdc0.w_dly_sig\[60\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4036 VGND tdc0.w_dly_sig\[115\] a_18673_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4037 VGND a_9907_2045# a_10075_1947# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4038 VGND tdc0.w_dly_sig\[118\] tdc0.w_dly_sig_n\[118\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4039 tdc0.w_dly_sig\[55\] tdc0.w_dly_sig\[53\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4040 VGND a_1830_14847# a_1788_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4041 a_14533_3855# a_13986_4129# a_14186_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4042 VGND tdc0.w_dly_sig\[3\] tdc0.w_dly_sig_n\[3\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4043 _023_ _001_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4044 tdc0.w_dly_sig\[10\] tdc0.w_dly_sig\[8\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4045 a_2030_17277# a_1591_16911# a_1945_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4046 VPWR tdc0.w_dly_sig\[122\] tdc0.w_dly_sig\[124\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4047 VPWR tdc0.w_dly_sig_n\[82\] tdc0.w_dly_sig_n\[84\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4048 VPWR tdc0.w_dly_sig\[87\] tdc0.w_dly_sig_n\[87\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4049 a_11122_7637# a_11780_7637# a_11714_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4051 VPWR clknet_4_7_0_clk a_8399_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4052 tdc0.w_dly_sig\[5\] tdc0.w_dly_sig_n\[4\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4054 VPWR net5 a_12134_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4055 tdc0.o_result\[117\] a_17711_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4056 tdc0.o_result\[3\] a_16331_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4057 tdc0.w_dly_sig\[28\] tdc0.w_dly_sig_n\[27\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4058 a_16600_9839# _096_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X4059 tdc0.w_dly_sig_n\[55\] tdc0.w_dly_sig\[55\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4060 tdc0.o_result\[8\] a_14675_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4061 VGND tdc0.w_dly_sig\[122\] a_18489_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4062 uo_out[6] a_12376_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4063 a_3417_8751# tdc0.w_dly_sig\[71\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4064 VPWR tdc0.w_dly_sig_n\[9\] tdc0.w_dly_sig_n\[11\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4065 a_13823_5193# _020_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4066 a_2156_9129# a_1757_8757# a_2030_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4067 VGND clknet_4_4_0_clk a_6191_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4068 VPWR tdc0.w_dly_sig_n\[115\] tdc0.w_dly_sig_n\[117\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4069 a_17935_6793# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4070 VGND tdc0.w_dly_sig\[51\] tdc0.w_dly_sig\[53\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4071 VGND a_3175_14165# a_3133_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4072 tdc0.w_dly_sig\[72\] tdc0.w_dly_sig_n\[71\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4073 a_17835_4631# a_18119_4617# a_18054_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4074 VPWR a_14388_13621# clknet_4_13_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4075 VGND tdc0.w_dly_sig\[107\] tdc0.w_dly_sig_n\[107\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4076 _002_ a_13183_6583# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4077 VPWR a_14664_6005# clknet_4_9_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4078 VPWR a_6826_17973# a_6755_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4079 VPWR a_8819_7637# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4080 VGND tdc0.w_dly_sig_n\[21\] tdc0.w_dly_sig\[22\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4081 a_17118_8751# a_16679_8757# a_17033_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4082 a_9366_10071# _077_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X4083 a_2489_11305# a_1499_10933# a_2363_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4084 tdc0.w_dly_sig_n\[25\] tdc0.w_dly_sig\[25\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4085 VGND tdc0.w_dly_sig_n\[74\] tdc0.w_dly_sig\[75\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4086 VPWR tdc0.w_dly_sig_n\[61\] tdc0.w_dly_sig\[62\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4087 tdc0.w_dly_sig_n\[40\] tdc0.w_dly_sig_n\[38\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4088 _016_ _003_ a_10595_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4089 VGND a_17359_1135# a_17527_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4090 VGND tdc0.w_dly_sig\[81\] tdc0.w_dly_sig\[83\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4091 VPWR tdc0.w_dly_sig\[39\] tdc0.w_dly_sig_n\[39\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4093 VGND net3 a_10515_7671# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4094 tdc0.w_dly_sig\[2\] tdc0.w_dly_sig_n\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4095 _058_ a_9411_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4096 tdc0.w_dly_sig_n\[65\] tdc0.w_dly_sig\[65\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4097 a_11504_7983# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.114 ps=1 w=0.65 l=0.15
X4098 a_11321_17775# tdc0.o_result\[23\] a_10975_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4099 VGND a_17739_4631# tdc0.o_result\[114\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4100 VGND tdc0.w_dly_sig_n\[0\] tdc0.w_dly_sig\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4101 VGND tdc0.w_dly_sig_n\[25\] tdc0.w_dly_sig_n\[27\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4102 a_14178_9839# a_13931_10217# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4103 tdc0.w_dly_sig\[70\] tdc0.w_dly_sig\[68\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4104 VGND a_7331_16189# a_7499_16091# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4105 a_16181_5461# net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X4106 VPWR a_11058_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4107 a_17567_13621# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4108 tdc0.w_dly_sig_n\[82\] tdc0.w_dly_sig\[82\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4109 tdc0.w_dly_sig\[86\] tdc0.w_dly_sig_n\[85\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4110 a_14510_12559# _086_ a_14676_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4111 a_1757_8757# a_1591_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4112 VPWR a_6043_5309# a_6211_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4113 VGND clknet_4_1_0_clk a_1407_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4114 a_14158_8319# a_13990_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4115 a_18581_12393# a_18034_12137# a_18234_12292# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4116 VGND _005_ a_14510_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4117 a_7561_13423# tdc0.o_result\[36\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4119 clknet_4_5_0_clk a_3348_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4121 a_8841_13109# a_8675_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4122 VGND _012_ a_11597_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X4124 a_4333_6581# a_4167_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4125 tdc0.w_dly_sig\[4\] tdc0.w_dly_sig_n\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4126 VPWR tdc0.w_dly_sig\[54\] tdc0.w_dly_sig_n\[54\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4127 a_5158_18365# a_4885_17999# a_5073_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4128 a_7369_4221# a_6835_3855# a_7274_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4129 tdc0.o_result\[22\] a_16239_18267# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4130 a_4774_17429# a_4606_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4131 a_14381_6031# _020_ a_13947_6183# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4132 VPWR a_18234_12292# a_18163_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4133 VPWR tdc0.w_dly_sig\[85\] tdc0.w_dly_sig_n\[85\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4135 VGND a_14676_12809# uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4136 a_12706_17455# a_12459_17833# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4137 tdc0.w_dly_sig\[56\] tdc0.w_dly_sig_n\[55\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4138 VGND a_12548_4917# clknet_4_8_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4139 VPWR tdc0.w_dly_sig\[117\] a_18489_6953# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4140 a_3927_8751# a_3229_8757# a_3670_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4141 tdc0.w_dly_sig_n\[6\] tdc0.w_dly_sig\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4142 VPWR tdc0.w_dly_sig\[74\] tdc0.w_dly_sig_n\[74\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4143 a_9209_9295# a_9043_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4144 VPWR a_18003_9661# a_18171_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4145 VGND tdc0.w_dly_sig_n\[13\] tdc0.w_dly_sig_n\[15\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4146 VPWR a_5851_13335# _042_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X4147 tdc0.w_dly_sig_n\[67\] tdc0.w_dly_sig\[67\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4148 tdc0.w_dly_sig\[71\] tdc0.w_dly_sig\[69\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4149 a_13795_10057# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4150 VGND tdc0.w_dly_sig_n\[108\] tdc0.w_dly_sig_n\[110\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4151 tdc0.w_dly_sig_n\[64\] tdc0.w_dly_sig\[64\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4152 tdc0.w_dly_sig_n\[4\] tdc0.w_dly_sig\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4153 VPWR tdc0.w_dly_sig\[105\] tdc0.w_dly_sig_n\[105\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4154 VGND tdc0.w_dly_sig_n\[26\] tdc0.w_dly_sig_n\[28\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4155 a_14729_4405# a_14563_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4156 VPWR a_4479_3311# a_4647_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4157 VGND tdc0.w_dly_sig\[106\] tdc0.w_dly_sig\[108\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4158 a_2673_4943# a_1683_4943# a_2547_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4159 a_4057_1679# a_3891_1679# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4160 a_8837_5807# tdc0.o_result\[32\] a_8491_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4161 VGND _007_ a_11137_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X4162 VPWR tdc0.w_dly_sig_n\[102\] tdc0.w_dly_sig\[103\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4163 VGND tdc0.w_dly_sig_n\[119\] tdc0.w_dly_sig\[120\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4165 a_9757_2543# tdc0.o_result\[85\] a_9411_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4166 VGND _042_ a_11987_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X4168 VGND tdc0.w_dly_sig\[48\] tdc0.w_dly_sig\[50\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4169 VPWR a_8603_8725# a_8519_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4170 a_3785_10927# tdc0.w_dly_sig\[56\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4171 VGND tdc0.w_dly_sig\[78\] tdc0.w_dly_sig\[80\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4172 a_17753_10383# a_17199_10357# a_17406_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4173 VPWR a_6963_4399# a_7131_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4174 a_17244_9129# a_16845_8757# a_17118_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4175 tdc0.w_dly_sig\[111\] tdc0.w_dly_sig\[109\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4176 tdc0.w_dly_sig\[99\] tdc0.w_dly_sig\[97\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4178 tdc0.w_dly_sig\[129\] tdc0.w_dly_sig\[127\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4179 VPWR tdc0.w_dly_sig\[50\] tdc0.w_dly_sig_n\[50\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4180 a_9953_17455# _029_ a_9807_17687# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X4181 a_4824_13481# a_4425_13109# a_4698_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4184 clknet_4_1_0_clk a_3790_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4185 VGND a_4923_4373# a_4881_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4187 VGND a_5031_6575# a_5199_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4188 VPWR tdc0.w_dly_sig_n\[72\] tdc0.w_dly_sig\[73\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4189 tdc0.w_dly_sig\[31\] tdc0.w_dly_sig\[29\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4190 a_7626_7637# a_7458_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4192 VGND a_3854_14847# a_3812_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4193 a_18077_4399# a_17739_4631# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4194 a_9650_1791# a_9482_2045# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4195 tdc0.w_dly_sig\[67\] tdc0.w_dly_sig_n\[66\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4196 tdc0.w_dly_sig_n\[17\] tdc0.w_dly_sig_n\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4197 tdc0.w_dly_sig\[122\] tdc0.w_dly_sig\[120\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4199 VGND tdc0.w_dly_sig\[126\] a_18121_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4200 tdc0.w_dly_sig_n\[105\] tdc0.w_dly_sig\[105\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4201 VGND a_6239_18151# tdc0.o_result\[18\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4202 VGND a_15170_4373# a_15128_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4203 a_16845_8757# a_16679_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4204 a_12530_17732# a_12323_17673# a_12706_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4205 tdc0.w_dly_sig\[16\] tdc0.w_dly_sig_n\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4206 VGND a_18027_12233# a_18034_12137# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4207 VGND tdc0.w_dly_sig_n\[50\] tdc0.w_dly_sig\[51\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4209 VPWR a_1830_9813# a_1757_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4210 a_9741_10357# _016_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X4211 a_11504_11445# _061_ a_11974_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4212 tdc0.w_dly_sig_n\[95\] tdc0.w_dly_sig_n\[93\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4213 a_5897_2045# a_5363_1679# a_5802_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4215 VPWR a_8695_10901# a_8611_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4216 VPWR a_7286_7119# clknet_4_3_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4217 a_12459_17833# a_12323_17673# a_12039_17687# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4218 _076_ a_11619_8867# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X4219 a_11338_14557# a_11023_14423# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4220 VGND tdc0.w_dly_sig_n\[91\] tdc0.w_dly_sig\[92\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4222 a_13429_12393# a_12882_12137# a_13082_12292# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4223 a_9650_7637# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.327 ps=1.65 w=1 l=0.15
X4224 VGND a_9006_1109# a_8964_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4225 tdc0.w_dly_sig\[21\] tdc0.w_dly_sig\[19\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4226 VPWR tdc0.w_dly_sig\[9\] tdc0.w_dly_sig\[11\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4227 a_2122_3133# a_1683_2767# a_2037_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4228 clknet_4_10_0_clk a_16412_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4229 a_11872_7093# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.176 ps=1.68 w=0.42 l=0.15
X4230 a_7825_3855# a_6835_3855# a_7699_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4231 tdc0.w_dly_sig\[107\] tdc0.w_dly_sig_n\[106\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4232 tdc0.w_dly_sig\[58\] tdc0.w_dly_sig_n\[57\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4233 a_17703_16745# a_17567_16585# a_17283_16599# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4234 VGND tdc0.w_dly_sig\[96\] tdc0.w_dly_sig\[98\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4235 VPWR a_7856_14165# clknet_4_7_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4236 a_2198_4373# a_2030_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4237 a_17279_14735# a_17059_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X4239 a_3698_12559# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4240 a_18475_4765# a_18255_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X4241 a_6538_4399# a_6265_4405# a_6453_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4242 VPWR a_12548_14165# clknet_4_12_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4243 VPWR tdc0.w_dly_sig\[32\] tdc0.w_dly_sig\[34\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4245 a_10585_10383# tdc0.o_result\[13\] a_10239_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4246 VGND tdc0.w_dly_sig\[73\] tdc0.w_dly_sig\[75\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4247 a_9297_17833# a_8307_17461# a_9171_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4250 a_5253_3855# a_5087_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4251 tdc0.w_dly_sig_n\[68\] tdc0.w_dly_sig\[68\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4252 a_15002_4399# a_14563_4405# a_14917_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4253 VGND net6 a_9389_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X4255 VPWR tdc0.w_dly_sig_n\[30\] tdc0.w_dly_sig\[31\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4256 VGND a_18003_9661# a_18171_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4257 a_13437_2601# a_12447_2229# a_13311_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4258 VGND net2 a_13919_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4260 a_15465_1679# a_15299_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4261 tdc0.w_dly_sig_n\[28\] tdc0.w_dly_sig\[28\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4262 clknet_4_4_0_clk a_3698_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4264 a_15162_5095# _082_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X4265 VPWR tdc0.w_dly_sig\[11\] tdc0.w_dly_sig\[13\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4266 VGND a_7856_14165# clknet_4_7_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4267 VPWR tdc0.w_dly_sig_n\[50\] tdc0.w_dly_sig_n\[52\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4268 _020_ a_8543_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X4269 a_8819_7637# _023_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X4270 tdc0.o_result\[94\] a_10259_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4271 VGND _089_ a_6835_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X4272 a_14349_10217# a_13802_9961# a_14002_10116# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4273 tdc0.w_dly_sig\[44\] tdc0.w_dly_sig\[42\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4274 a_8838_1135# a_8399_1141# a_8753_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4276 VGND a_11058_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4277 a_2290_5055# a_2122_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4278 a_13989_3689# a_12999_3317# a_13863_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4279 tdc0.o_result\[34\] a_8051_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4280 a_11609_4399# tdc0.o_result\[78\] a_11527_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4281 tdc0.w_dly_sig\[96\] tdc0.w_dly_sig_n\[95\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4282 _057_ a_10239_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4284 tdc0.w_dly_sig_n\[87\] tdc0.w_dly_sig_n\[85\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4285 net1 a_18187_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4286 VPWR tdc0.w_dly_sig\[116\] tdc0.w_dly_sig\[118\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4287 a_14829_7663# tdc0.o_result\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X4288 _024_ a_7479_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4289 a_17187_16599# a_17283_16599# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4290 a_10055_2223# _028_ a_10137_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4291 tdc0.w_dly_sig_n\[89\] tdc0.w_dly_sig_n\[87\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4292 tdc0.w_dly_sig\[70\] tdc0.w_dly_sig_n\[69\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4293 a_12726_6895# a_11987_6575# a_12612_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.137 ps=1.07 w=0.65 l=0.15
X4294 a_2511_10633# _026_ a_2593_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4296 VGND a_14250_6549# a_14208_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4297 VPWR tdc0.w_dly_sig\[110\] tdc0.w_dly_sig\[112\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4298 clknet_0_clk a_11058_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4299 VGND clknet_4_1_0_clk a_3155_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4300 a_9006_1109# a_8838_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4302 VPWR a_12284_9545# uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4304 VGND a_14031_3285# a_13989_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4305 VGND tdc0.w_dly_sig\[45\] tdc0.w_dly_sig_n\[45\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4306 tdc0.w_dly_sig\[73\] tdc0.w_dly_sig_n\[72\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R16 VPWR tt_um_hpretl_tt06_tdc_15.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4310 VPWR tdc0.w_dly_sig_n\[125\] tdc0.w_dly_sig\[126\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4311 a_2248_2767# a_1849_2767# a_2122_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4312 a_6817_9295# a_6651_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4313 a_1205_9295# a_1039_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4314 a_1903_9661# a_1039_9295# a_1646_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4315 VGND a_18187_10901# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4316 clknet_4_8_0_clk a_12548_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4317 a_14645_5487# tdc0.o_result\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X4318 a_8289_16373# a_8123_16373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4319 a_11057_9071# tdc0.o_result\[65\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4320 a_2198_4373# a_2030_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4321 tdc0.w_dly_sig\[6\] tdc0.w_dly_sig_n\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4322 VPWR tdc0.w_dly_sig\[61\] tdc0.w_dly_sig\[63\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4323 a_9493_12809# tdc0.o_result\[63\] a_9411_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4324 a_4425_13109# a_4259_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4325 a_5859_7485# a_5161_7119# a_5602_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4326 a_3413_10383# a_3247_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4327 clknet_4_5_0_clk a_3348_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4328 a_9332_14569# a_8933_14197# a_9206_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4329 VPWR tdc0.w_dly_sig_n\[59\] tdc0.w_dly_sig_n\[61\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4330 a_5441_14735# tdc0.w_dly_sig\[39\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4331 a_8574_4676# a_8374_4521# a_8723_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4332 a_9319_7485# _002_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4333 a_2773_17455# tdc0.w_dly_sig\[46\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4334 a_6537_17775# tdc0.o_result\[18\] a_6191_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4335 a_15170_4373# a_15002_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4336 a_9217_5487# tdc0.o_result\[34\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X4337 tdc0.w_dly_sig_n\[113\] tdc0.w_dly_sig\[113\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4339 clknet_0_clk a_11058_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4340 VPWR a_14715_15797# a_14722_16097# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4341 a_6955_8573# a_6173_8207# a_6871_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4342 VPWR a_18187_10901# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4343 VPWR tdc0.w_dly_sig\[19\] a_7173_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4344 VGND a_14952_8751# uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4345 tdc0.o_result\[54\] a_5291_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4346 VGND tdc0.w_dly_sig_n\[109\] tdc0.w_dly_sig\[110\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4347 VGND a_6947_6549# a_6905_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4348 a_8543_7093# _003_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.143 ps=1.33 w=0.42 l=0.15
X4350 a_8010_8751# a_7571_8757# a_7925_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4351 tdc0.w_dly_sig\[40\] tdc0.w_dly_sig\[38\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4352 a_15753_6281# _064_ a_15657_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4353 VPWR tdc0.w_dly_sig_n\[56\] tdc0.w_dly_sig\[57\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4354 tdc0.o_result\[54\] a_5291_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4355 VPWR a_5199_17429# a_5115_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4356 a_9631_4221# a_8767_3855# a_9374_3967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4357 a_5253_3855# a_5087_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4358 a_12792_6549# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.312 ps=2.12 w=0.42 l=0.15
X4359 a_9282_13077# a_9114_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4361 a_7571_17161# _029_ a_7653_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4362 a_7442_3967# a_7274_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4364 a_4061_4943# tdc0.w_dly_sig\[70\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4366 VPWR a_2455_4399# a_2623_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4367 a_2455_4399# a_1757_4405# a_2198_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4368 VGND a_13947_6183# _083_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4369 tdc0.w_dly_sig\[77\] tdc0.w_dly_sig\[75\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4370 a_15653_10383# tdc0.w_dly_sig\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4371 VPWR tdc0.w_dly_sig\[11\] tdc0.w_dly_sig_n\[11\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4372 VPWR tdc0.w_dly_sig_n\[94\] tdc0.w_dly_sig_n\[96\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4373 _028_ a_9485_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.143 ps=1.33 w=1 l=0.15
X4374 tdc0.o_result\[48\] a_2255_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4375 a_8964_1513# a_8565_1141# a_8838_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4376 tdc0.w_dly_sig_n\[81\] tdc0.w_dly_sig_n\[79\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4377 tdc0.w_dly_sig\[30\] tdc0.w_dly_sig\[28\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4379 VGND tdc0.w_dly_sig_n\[116\] tdc0.w_dly_sig_n\[118\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4380 a_16332_12015# _066_ a_16166_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X4381 a_16197_17999# a_15207_17999# a_16071_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4382 VGND a_11159_4943# _013_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4383 VGND a_8500_4917# clknet_4_2_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4384 a_1945_16911# tdc0.w_dly_sig\[48\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4385 a_10975_5487# _001_ a_11225_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4386 VPWR a_16412_6549# clknet_4_10_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4387 VGND tdc0.w_dly_sig_n\[37\] tdc0.w_dly_sig\[38\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4388 a_18255_4777# a_18119_4617# a_17835_4631# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4389 VPWR a_14335_15975# tdc0.o_result\[25\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4390 VPWR tdc0.w_dly_sig_n\[109\] tdc0.w_dly_sig_n\[111\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4391 clknet_4_13_0_clk a_14388_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X4392 VPWR a_16732_11445# _356_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4393 VPWR tdc0.o_result\[100\] a_14375_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
R17 uio_oe[5] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4394 VGND a_14507_14191# a_14675_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4396 a_8473_17461# a_8307_17461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4398 a_4146_5309# a_3707_4943# a_4061_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4399 VPWR a_2439_6549# a_2355_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4400 VPWR tdc0.w_dly_sig_n\[58\] tdc0.w_dly_sig_n\[60\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4401 _060_ a_10055_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4402 clknet_4_14_0_clk a_17314_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4403 a_14729_17461# a_14563_17461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4404 a_1903_11837# a_1039_11471# a_1646_11583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4405 VGND tdc0.w_dly_sig_n\[13\] tdc0.w_dly_sig\[14\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4406 VPWR a_5970_12671# a_5897_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4407 VGND tdc0.w_dly_sig_n\[45\] tdc0.w_dly_sig_n\[47\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4408 tdc0.o_result\[10\] a_14031_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4409 _097_ a_5823_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4411 VGND a_3348_13077# clknet_4_5_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4412 VPWR a_7699_6397# a_7867_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4413 a_13269_7779# _049_ a_13173_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4414 a_9650_7637# _002_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.21 ps=1.42 w=1 l=0.15
X4415 a_17985_12015# a_17647_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4416 a_5207_13103# a_4425_13109# a_5123_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4417 tdc0.w_dly_sig_n\[114\] tdc0.w_dly_sig_n\[112\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4418 tdc0.w_dly_sig_n\[88\] tdc0.w_dly_sig_n\[86\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4419 tdc0.w_dly_sig_n\[127\] tdc0.w_dly_sig\[127\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4420 tdc0.w_dly_sig_n\[5\] tdc0.w_dly_sig_n\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4421 a_10147_16073# net6 a_10229_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4422 a_7350_3285# a_7182_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4423 a_1573_11837# a_1039_11471# a_1478_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4424 VPWR tdc0.w_dly_sig_n\[126\] tdc0.w_dly_sig_n\[128\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4425 tdc0.w_dly_sig\[118\] tdc0.w_dly_sig\[116\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4426 VGND a_2290_2879# a_2248_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4427 a_5161_7119# a_4995_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4428 VPWR tdc0.w_dly_sig_n\[88\] tdc0.w_dly_sig\[89\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4429 VPWR clknet_4_5_0_clk a_2419_17461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4430 a_16301_6281# _020_ a_16155_6183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X4431 net10 a_13603_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4432 tdc0.w_dly_sig\[78\] tdc0.w_dly_sig\[76\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4433 a_11414_2045# a_10975_1679# a_11329_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4434 a_8543_7093# a_8995_7093# a_8953_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4435 tdc0.w_dly_sig\[54\] tdc0.w_dly_sig\[52\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4436 VPWR tdc0.w_dly_sig_n\[77\] tdc0.w_dly_sig\[78\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4437 VGND tdc0.w_dly_sig_n\[42\] tdc0.w_dly_sig\[43\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4438 _068_ a_7571_17161# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4439 VPWR a_18234_3588# a_18163_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4440 VPWR a_6706_4373# a_6633_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4441 tdc0.o_result\[26\] a_15595_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4442 VGND a_9459_4631# tdc0.o_result\[111\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4443 VGND tdc0.w_dly_sig\[59\] tdc0.w_dly_sig\[61\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4444 tdc0.w_dly_sig_n\[24\] tdc0.w_dly_sig_n\[22\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4445 a_9121_14191# tdc0.w_dly_sig\[30\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4446 VPWR tdc0.w_dly_sig_n\[91\] tdc0.w_dly_sig_n\[93\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4447 a_8921_4777# a_8367_4617# a_8574_4676# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4448 tdc0.w_dly_sig\[65\] tdc0.w_dly_sig_n\[64\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4449 VGND a_17130_14709# a_17059_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4450 VPWR tdc0.w_dly_sig\[67\] tdc0.w_dly_sig_n\[67\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4451 a_15170_4373# a_15002_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4452 VPWR a_14388_13621# clknet_4_13_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4453 a_1853_10927# tdc0.w_dly_sig\[52\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4454 VPWR tdc0.w_dly_sig_n\[103\] tdc0.w_dly_sig\[104\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4455 tdc0.w_dly_sig\[6\] tdc0.w_dly_sig\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4456 tdc0.w_dly_sig\[18\] tdc0.w_dly_sig\[16\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4457 a_8136_9129# a_7737_8757# a_8010_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4458 a_7607_3311# a_6909_3317# a_7350_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4459 tdc0.w_dly_sig\[59\] tdc0.w_dly_sig\[57\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4460 a_9597_9955# _078_ a_9501_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4461 VGND tdc0.w_dly_sig_n\[35\] tdc0.w_dly_sig\[36\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4462 tdc0.w_dly_sig_n\[76\] tdc0.w_dly_sig\[76\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4463 VGND a_17774_13621# a_17703_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4464 a_17743_12247# a_18027_12233# a_17962_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4465 a_17555_6807# a_17651_6807# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4466 a_10747_14735# a_10527_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X4468 tdc0.w_dly_sig\[22\] tdc0.w_dly_sig_n\[21\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4469 VGND tdc0.w_dly_sig_n\[65\] tdc0.w_dly_sig_n\[67\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4470 tdc0.w_dly_sig\[62\] tdc0.w_dly_sig_n\[61\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4471 VGND clknet_4_2_0_clk a_8399_1141# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4472 VGND tdc0.w_dly_sig\[92\] tdc0.w_dly_sig_n\[92\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4473 tdc0.w_dly_sig\[119\] tdc0.w_dly_sig\[117\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4474 _040_ a_10147_16073# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4475 VGND a_14002_10116# a_13931_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4476 VPWR a_14250_14165# a_14177_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4477 a_11869_8867# _073_ a_11797_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4478 VPWR clknet_4_13_0_clk a_14563_17461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4479 tdc0.w_dly_sig_n\[80\] tdc0.w_dly_sig_n\[78\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4480 VGND _037_ a_11435_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X4481 a_3133_14569# a_2143_14197# a_3007_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4483 VPWR tdc0.w_dly_sig\[5\] tdc0.w_dly_sig_n\[5\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4485 a_15427_4399# a_14729_4405# a_15170_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4486 VPWR a_15427_4399# a_15595_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4487 VGND tdc0.o_result\[113\] a_12633_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4488 a_12201_8457# _002_ a_12117_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4489 tdc0.w_dly_sig_n\[116\] tdc0.w_dly_sig\[116\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4490 tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4491 a_7399_17833# a_7263_17673# a_6979_17687# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4492 a_1757_15101# a_1223_14735# a_1662_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4493 tdc0.w_dly_sig_n\[27\] tdc0.w_dly_sig_n\[25\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4494 a_12518_7119# a_12263_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.312 ps=2.12 w=1 l=0.15
X4495 a_12483_4221# a_11619_3855# a_12226_3967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4496 tdc0.o_result\[77\] a_2255_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4497 VGND a_8051_7637# a_8009_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4498 VPWR tdc0.w_dly_sig\[49\] tdc0.w_dly_sig_n\[49\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4499 a_2213_10217# a_1223_9845# a_2087_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4500 clknet_4_5_0_clk a_3348_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4501 tdc0.w_dly_sig\[115\] tdc0.w_dly_sig\[113\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4502 a_6630_10927# a_6191_10933# a_6545_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4503 VGND a_12376_8751# uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4504 a_7737_8757# a_7571_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4505 VPWR a_9799_4123# a_9715_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4507 VPWR tdc0.w_dly_sig\[126\] tdc0.w_dly_sig_n\[126\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4509 a_9650_7637# a_9503_7663# a_10291_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.143 ps=1.09 w=0.65 l=0.15
X4510 uo_out[4] a_14952_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X4511 VPWR tdc0.w_dly_sig\[90\] tdc0.w_dly_sig_n\[90\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4512 VPWR tdc0.w_dly_sig\[93\] tdc0.w_dly_sig_n\[93\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4513 VPWR tdc0.w_dly_sig_n\[102\] tdc0.w_dly_sig_n\[104\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4514 a_14510_12559# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4515 VGND tdc0.w_dly_sig_n\[110\] tdc0.w_dly_sig\[111\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4516 a_4272_4943# a_3873_4943# a_4146_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4517 a_1895_12015# a_1113_12021# a_1811_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4518 a_17125_1679# tdc0.w_dly_sig\[104\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4519 a_6917_12809# _090_ a_6835_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
R18 tt_um_hpretl_tt06_tdc_16.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4520 VGND a_9339_17429# a_9297_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4521 a_1646_11583# a_1478_11837# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4522 VGND clknet_4_7_0_clk a_8675_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4523 VPWR tdc0.w_dly_sig_n\[75\] tdc0.w_dly_sig\[76\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4524 a_10349_15101# a_10011_14887# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4525 VGND a_12199_4631# _080_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4526 tdc0.w_dly_sig_n\[54\] tdc0.w_dly_sig\[54\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4528 VGND a_7867_4123# a_7825_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4529 VGND clknet_4_2_0_clk a_8767_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4530 VGND a_17527_1109# a_17485_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4531 VGND _002_ a_11343_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4532 VPWR a_1646_11583# a_1573_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4533 VGND tdc0.w_dly_sig_n\[63\] tdc0.w_dly_sig\[64\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4534 a_16323_12559# a_16194_12833# a_15903_12533# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4535 a_16399_5487# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4536 tdc0.w_dly_sig\[24\] tdc0.w_dly_sig_n\[23\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4538 clknet_4_9_0_clk a_14664_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4539 a_2685_12335# tdc0.o_result\[72\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4540 VPWR tdc0.w_dly_sig_n\[66\] tdc0.w_dly_sig\[67\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4541 a_13825_7779# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X4542 VGND tdc0.w_dly_sig\[7\] tdc0.w_dly_sig_n\[7\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4543 VPWR clknet_4_6_0_clk a_5823_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4544 VGND a_12134_6549# _010_ VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4545 VGND tdc0.w_dly_sig_n\[0\] tdc0.w_dly_sig\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4546 VGND a_15630_14847# a_15588_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4547 a_6633_4399# a_6099_4405# a_6538_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4548 VPWR a_11490_6005# _026_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X4549 a_12210_9071# _046_ a_12376_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4550 tdc0.w_dly_sig_n\[85\] tdc0.w_dly_sig_n\[83\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4551 _070_ a_2603_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4552 VGND _087_ a_6835_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X4553 a_11540_1679# a_11141_1679# a_11414_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4554 a_12148_6005# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.312 ps=2.12 w=0.42 l=0.15
X4555 VGND a_13795_10057# a_13802_9961# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4556 a_9293_8457# _024_ a_9221_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4558 a_16578_13103# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4559 a_4755_2045# a_3891_1679# a_4498_1791# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4560 tdc0.w_dly_sig_n\[68\] tdc0.w_dly_sig_n\[66\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4562 tdc0.w_dly_sig\[123\] tdc0.w_dly_sig_n\[122\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4563 a_16915_10357# a_17199_10357# a_17134_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4564 a_15465_1679# a_15299_1679# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4565 tdc0.w_dly_sig_n\[119\] tdc0.w_dly_sig\[119\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4566 a_12833_12015# a_12495_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4567 VPWR tdc0.o_result\[12\] a_15473_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X4568 tdc0.w_dly_sig_n\[56\] tdc0.w_dly_sig_n\[54\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4569 a_5031_17455# a_4333_17461# a_4774_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4570 _098_ a_6099_16367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4571 VGND tdc0.w_dly_sig\[61\] tdc0.w_dly_sig_n\[61\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4572 a_11786_12015# a_11539_12393# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4573 VGND clknet_4_9_0_clk a_13643_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4574 tdc0.o_result\[68\] a_6211_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4575 VGND tdc0.w_dly_sig_n\[71\] tdc0.w_dly_sig_n\[73\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4576 VPWR tdc0.w_dly_sig_n\[26\] tdc0.w_dly_sig\[27\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4577 tdc0.w_dly_sig\[79\] tdc0.w_dly_sig\[77\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4578 a_7182_9839# a_6909_9845# a_7097_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4579 a_15971_15101# a_15189_14735# a_15887_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4580 a_7185_7669# a_7019_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4581 a_6725_10927# a_6191_10933# a_6630_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4582 tdc0.w_dly_sig_n\[56\] tdc0.w_dly_sig\[56\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4583 tdc0.w_dly_sig\[120\] tdc0.w_dly_sig_n\[119\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4584 a_5859_7485# a_4995_7119# a_5602_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4585 a_11987_10633# _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4586 a_10321_12015# tdc0.o_result\[79\] a_10239_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4587 tdc0.w_dly_sig_n\[93\] tdc0.w_dly_sig\[93\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4588 a_15427_4399# a_14563_4405# a_15170_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4589 tdc0.w_dly_sig\[104\] tdc0.w_dly_sig\[102\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4590 a_2037_1135# tdc0.w_dly_sig\[83\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4591 VPWR _022_ a_10057_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4592 VPWR tdc0.w_dly_sig_n\[46\] tdc0.w_dly_sig\[47\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4593 tdc0.w_dly_sig_n\[90\] tdc0.w_dly_sig_n\[88\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4594 clknet_4_1_0_clk a_3790_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4595 clknet_4_1_0_clk a_3790_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4596 a_12886_2223# a_12613_2229# a_12801_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4597 VPWR tdc0.w_dly_sig\[97\] tdc0.w_dly_sig\[99\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4599 VGND a_4038_1109# a_3996_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4600 a_16332_9839# _005_ a_16248_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4601 tdc0.w_dly_sig_n\[41\] tdc0.w_dly_sig\[41\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4602 _071_ a_7755_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4603 VGND tdc0.w_dly_sig_n\[43\] tdc0.w_dly_sig\[44\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4605 a_5928_12559# a_5529_12559# a_5802_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4606 VGND a_6503_14013# a_6671_13915# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4607 VPWR clknet_4_6_0_clk a_6743_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4608 a_4613_13103# tdc0.w_dly_sig\[55\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4609 tdc0.o_result\[89\] a_7591_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4610 a_9263_1135# a_8399_1141# a_9006_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4611 tdc0.w_dly_sig_n\[107\] tdc0.w_dly_sig\[107\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4612 VPWR net11 a_14645_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4613 a_9757_12559# tdc0.o_result\[31\] a_9411_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4614 _019_ _001_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4615 VPWR tdc0.w_dly_sig_n\[10\] tdc0.w_dly_sig\[11\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4616 VPWR tdc0.w_dly_sig_n\[78\] tdc0.w_dly_sig\[79\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4617 _036_ a_9503_11043# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X4618 VPWR tdc0.w_dly_sig\[50\] tdc0.w_dly_sig\[52\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R19 VGND uio_oe[4] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4619 VGND a_4314_5055# a_4272_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4620 a_2547_5309# a_1683_4943# a_2290_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4623 VGND a_11122_7637# _029_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4624 a_3873_13647# a_3707_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4626 VGND tdc0.w_dly_sig\[62\] tdc0.w_dly_sig\[64\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4627 VPWR tdc0.w_dly_sig_n\[6\] tdc0.w_dly_sig\[7\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4628 VPWR tdc0.w_dly_sig\[116\] a_17385_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4629 VPWR tdc0.w_dly_sig\[88\] tdc0.w_dly_sig\[90\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4630 VPWR clknet_4_2_0_clk a_8767_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4631 tdc0.o_result\[44\] a_4555_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4632 VPWR tdc0.w_dly_sig\[107\] a_14533_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4633 a_17865_8457# _015_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X4634 VPWR tdc0.w_dly_sig_n\[113\] tdc0.w_dly_sig\[114\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4635 a_13606_5461# a_13438_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4636 tdc0.w_dly_sig_n\[33\] tdc0.w_dly_sig_n\[31\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4637 a_5326_18111# a_5158_18365# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4638 VGND tdc0.w_dly_sig\[25\] tdc0.w_dly_sig\[27\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4639 tdc0.w_dly_sig_n\[104\] tdc0.w_dly_sig_n\[102\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4640 a_17753_10383# a_17206_10657# a_17406_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4641 VGND a_16155_17687# _047_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4642 VGND a_13151_11145# a_13158_11049# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4643 VGND a_2071_11739# a_2029_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4644 a_14526_2197# a_14358_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4645 VPWR tdc0.w_dly_sig_n\[69\] tdc0.w_dly_sig\[70\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4646 VPWR tdc0.w_dly_sig\[15\] a_11957_14569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4647 tdc0.w_dly_sig\[33\] tdc0.w_dly_sig\[31\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4648 clknet_4_11_0_clk a_16762_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4649 a_2171_9839# a_1389_9845# a_2087_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4650 a_12613_2229# a_12447_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4651 a_3870_1135# a_3431_1141# a_3785_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4652 a_18071_10217# a_17935_10057# a_17651_10071# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4653 VGND a_17187_2919# tdc0.o_result\[110\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4654 VGND tdc0.w_dly_sig\[44\] tdc0.w_dly_sig_n\[44\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4655 uo_out[6] a_12376_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X4656 tdc0.w_dly_sig_n\[1\] tdc0.w_dly_sig\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4657 a_11610_12292# a_11403_12233# a_11786_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4658 VPWR tdc0.w_dly_sig\[84\] tdc0.w_dly_sig_n\[84\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4659 VPWR tdc0.w_dly_sig_n\[21\] tdc0.w_dly_sig_n\[23\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4660 a_5951_4221# a_5087_3855# a_5694_3967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4661 a_2037_2767# tdc0.w_dly_sig\[82\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4662 VGND net28 a_10585_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X4663 tdc0.w_dly_sig_n\[72\] tdc0.w_dly_sig\[72\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4664 VPWR _097_ a_6717_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4665 VGND a_15170_17429# a_15128_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4666 a_18121_13647# a_17574_13921# a_17774_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4667 VPWR a_6798_10901# a_6725_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4668 VPWR tdc0.w_dly_sig\[126\] tdc0.w_dly_sig\[128\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4669 uo_out[7] a_11504_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4670 a_2125_17277# a_1591_16911# a_2030_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4672 a_8543_7093# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.128 ps=1.03 w=0.42 l=0.15
X4673 a_3781_15101# a_3247_14735# a_3686_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4674 VGND _022_ a_7825_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X4675 a_11539_12393# a_11403_12233# a_11119_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4676 VPWR tdc0.w_dly_sig_n\[52\] tdc0.w_dly_sig_n\[54\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4677 a_18397_14569# a_17843_14409# a_18050_14468# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4678 tdc0.w_dly_sig\[75\] tdc0.w_dly_sig\[73\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4679 VGND a_14195_7663# net11 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4680 tdc0.w_dly_sig\[56\] tdc0.w_dly_sig\[54\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4681 a_18121_13647# a_17567_13621# a_17774_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4682 a_2213_14735# a_1223_14735# a_2087_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4683 a_2106_10901# a_1938_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4684 VPWR tdc0.o_result\[7\] a_12326_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X4685 VGND a_7223_10901# a_7181_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4686 a_14507_6575# a_13643_6581# a_14250_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4687 a_13086_11293# a_12771_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4688 a_12644_8751# _051_ a_12376_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4689 VPWR a_18326_4676# a_18255_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4690 VGND clk a_11058_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4691 tdc0.w_dly_sig\[57\] tdc0.w_dly_sig\[55\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4692 VGND clknet_4_0_0_clk a_1683_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4693 VPWR a_9263_16189# a_9431_16091# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4694 a_6913_2223# tdc0.w_dly_sig\[90\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4695 tdc0.w_dly_sig\[13\] tdc0.w_dly_sig\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4696 net7 a_11027_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4697 tdc0.w_dly_sig\[59\] tdc0.w_dly_sig_n\[58\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4698 VGND tdc0.w_dly_sig\[33\] tdc0.w_dly_sig_n\[33\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4699 a_5823_5487# net7 a_5905_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4700 VGND tdc0.w_dly_sig\[2\] a_17753_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4701 a_17490_18365# a_17243_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4702 a_15381_5487# net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X4703 VPWR tdc0.w_dly_sig_n\[56\] tdc0.w_dly_sig_n\[58\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4704 tdc0.w_dly_sig\[72\] tdc0.w_dly_sig\[70\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4705 VGND net2 a_12810_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.107 ps=0.98 w=0.65 l=0.15
X4707 a_4606_17455# a_4333_17461# a_4521_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4709 VPWR a_12651_4123# a_12567_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4710 a_6821_15823# tdc0.w_dly_sig\[42\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4711 _023_ net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4712 a_10321_9071# tdc0.o_result\[94\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4713 VPWR clknet_4_7_0_clk a_8859_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4714 tdc0.w_dly_sig_n\[99\] tdc0.w_dly_sig_n\[97\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4715 clknet_0_clk a_11058_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4716 a_13605_4917# net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X4717 VGND a_14415_8573# a_14583_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4718 VPWR tdc0.w_dly_sig_n\[2\] tdc0.w_dly_sig\[3\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4719 VGND tdc0.w_dly_sig\[47\] tdc0.w_dly_sig_n\[47\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4720 tdc0.w_dly_sig_n\[80\] tdc0.w_dly_sig\[80\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4721 VPWR tdc0.w_dly_sig_n\[98\] tdc0.w_dly_sig_n\[100\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4722 VGND tdc0.w_dly_sig\[55\] tdc0.w_dly_sig_n\[55\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4723 VGND a_10391_14709# a_10398_15009# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4724 VGND a_18187_10901# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4725 a_5161_7119# a_4995_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4726 tdc0.w_dly_sig_n\[0\] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4727 VPWR tdc0.w_dly_sig_n\[112\] tdc0.w_dly_sig\[113\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4728 VPWR tdc0.w_dly_sig_n\[49\] tdc0.w_dly_sig\[50\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4729 a_7933_12809# _069_ a_7837_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4730 tdc0.w_dly_sig\[71\] tdc0.w_dly_sig_n\[70\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4731 VGND a_11023_12247# tdc0.o_result\[9\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4733 a_12548_4917# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4736 VPWR tdc0.w_dly_sig\[18\] tdc0.w_dly_sig_n\[18\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4738 a_3996_1513# a_3597_1141# a_3870_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4739 VGND a_13606_5461# a_13564_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4740 VGND tdc0.w_dly_sig\[13\] tdc0.w_dly_sig\[15\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4741 tdc0.w_dly_sig_n\[111\] tdc0.w_dly_sig\[111\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4742 VPWR a_4923_1947# a_4839_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4743 VPWR tdc0.w_dly_sig_n\[64\] tdc0.w_dly_sig_n\[66\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4744 a_5721_6031# tdc0.o_result\[66\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4745 a_18179_8983# tdc0.o_result\[101\] a_18325_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X4746 a_16570_12925# a_16323_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4747 VPWR a_2198_17023# a_2125_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4748 a_16451_7271# a_16547_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4749 VPWR a_3854_14847# a_3781_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4750 tdc0.w_dly_sig_n\[20\] tdc0.w_dly_sig_n\[18\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4751 tdc0.w_dly_sig\[89\] tdc0.w_dly_sig\[87\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4752 a_3329_12015# tdc0.o_result\[50\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X4753 a_17661_17999# a_17107_17973# a_17314_17973# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4754 VGND _001_ _016_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4755 a_7829_10933# a_7663_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4756 tdc0.w_dly_sig_n\[16\] tdc0.w_dly_sig\[16\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4757 a_6265_4405# a_6099_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4758 VGND clknet_4_4_0_clk a_3247_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4759 VPWR tdc0.w_dly_sig\[10\] tdc0.w_dly_sig_n\[10\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4760 VGND tdc0.w_dly_sig\[51\] tdc0.w_dly_sig_n\[51\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4761 a_11057_17775# tdc0.o_result\[47\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4762 VPWR a_7350_9813# a_7277_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4763 VGND tdc0.w_dly_sig\[56\] tdc0.w_dly_sig\[58\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4764 a_7085_12809# _088_ a_7013_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4765 tdc0.w_dly_sig_n\[78\] tdc0.w_dly_sig_n\[76\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4766 VPWR tdc0.w_dly_sig_n\[51\] tdc0.w_dly_sig\[52\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R20 uio_oe[7] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4767 VGND clknet_4_1_0_clk a_3063_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4768 net1 a_18187_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4769 VPWR a_15595_4373# a_15511_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4770 a_11422_5487# a_11642_5461# _019_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4771 VGND tdc0.w_dly_sig_n\[122\] tdc0.w_dly_sig_n\[124\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4772 VPWR a_17187_2919# tdc0.o_result\[110\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4773 a_13914_14735# a_13599_14887# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4774 a_7350_3285# a_7182_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4775 tdc0.w_dly_sig_n\[100\] tdc0.w_dly_sig_n\[98\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4776 VGND tdc0.w_dly_sig_n\[55\] tdc0.w_dly_sig\[56\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4778 a_17314_17973# a_17107_17973# a_17490_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4779 VGND _001_ a_9503_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4780 VGND tdc0.w_dly_sig_n\[0\] tdc0.w_dly_sig\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4781 a_11873_4719# tdc0.o_result\[102\] a_11527_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4782 a_7641_9295# a_6651_9295# a_7515_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4783 net28 a_12574_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X4785 a_15419_7895# tdc0.o_result\[110\] a_15565_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X4786 VPWR tdc0.w_dly_sig\[82\] tdc0.w_dly_sig\[84\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4787 VGND a_17739_7895# tdc0.o_result\[118\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4788 tdc0.w_dly_sig_n\[58\] tdc0.w_dly_sig\[58\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4789 tdc0.w_dly_sig_n\[11\] tdc0.w_dly_sig\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4790 a_12877_17833# a_12323_17673# a_12530_17732# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4791 VPWR clknet_4_0_0_clk a_1683_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4792 a_16381_8207# tdc0.o_result\[27\] a_16035_8457# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4793 VGND tdc0.w_dly_sig_n\[35\] tdc0.w_dly_sig_n\[37\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4794 a_4885_17999# a_4719_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4795 a_11329_1679# tdc0.w_dly_sig\[98\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4797 a_17243_17999# a_17107_17973# a_16823_17973# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4798 VPWR a_9431_1109# a_9347_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4799 VGND a_2087_15101# a_2255_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4800 VGND a_4279_15003# a_4237_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4801 VGND tdc0.w_dly_sig_n\[24\] tdc0.w_dly_sig\[25\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4802 a_1570_13103# a_1131_13109# a_1485_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4803 tdc0.w_dly_sig\[92\] tdc0.w_dly_sig_n\[91\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4804 a_18142_10116# a_17942_9961# a_18291_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4805 tdc0.w_dly_sig\[48\] tdc0.w_dly_sig\[46\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4806 _026_ a_11490_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4807 VPWR a_12171_5487# net8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4808 a_6755_17999# a_6626_18273# a_6335_17973# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4809 VPWR tdc0.w_dly_sig_n\[90\] tdc0.w_dly_sig_n\[92\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4810 a_17774_2741# a_17567_2741# a_17950_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4811 a_11597_15599# tdc0.o_result\[25\] a_11251_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4812 tdc0.w_dly_sig_n\[108\] tdc0.w_dly_sig\[108\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4813 VPWR a_2715_5211# a_2631_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4814 a_5529_12559# a_5363_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
R21 uio_oe[2] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4816 VPWR clknet_4_7_0_clk a_8307_17461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4817 a_11456_10927# _036_ a_11290_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X4818 a_13705_11305# a_13158_11049# a_13358_11204# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4819 VPWR tdc0.w_dly_sig\[116\] tdc0.w_dly_sig_n\[116\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4820 VGND a_3348_13077# clknet_4_5_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4821 VPWR a_10391_14709# a_10398_15009# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4822 tdc0.w_dly_sig_n\[112\] tdc0.w_dly_sig\[112\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4824 a_13606_5461# a_13438_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4825 VPWR tdc0.w_dly_sig\[29\] tdc0.w_dly_sig_n\[29\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4826 VGND a_4479_3311# a_4647_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4827 a_4061_4943# tdc0.w_dly_sig\[70\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4828 VGND a_4647_3285# a_4605_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4829 a_6181_16367# tdc0.o_result\[43\] a_6099_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4830 a_4513_15657# a_3523_15285# a_4387_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4831 VPWR net28 a_11057_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4832 a_8399_12809# _013_ a_8481_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4833 VGND tdc0.w_dly_sig_n\[54\] tdc0.w_dly_sig\[55\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4834 VGND clknet_4_0_0_clk a_3431_1141# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4835 a_1757_16911# a_1591_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4836 VPWR ui_in[3] a_12999_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4837 a_2030_4399# a_1591_4405# a_1945_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4838 VGND _022_ a_10044_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4839 a_16394_12533# a_16187_12533# a_16570_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4840 a_6545_10927# tdc0.w_dly_sig\[60\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4841 a_10229_16073# tdc0.o_result\[37\] a_10147_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4842 a_16117_8457# tdc0.o_result\[107\] a_16035_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4843 a_11154_5095# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X4844 tdc0.w_dly_sig_n\[128\] tdc0.w_dly_sig_n\[126\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4845 a_10505_5193# tdc0.o_result\[71\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X4847 _012_ a_12518_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4848 tdc0.w_dly_sig\[105\] tdc0.w_dly_sig_n\[104\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4849 _048_ a_5087_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4850 a_16323_12559# a_16187_12533# a_15903_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4851 VPWR a_16412_6549# clknet_4_10_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4852 VPWR a_14388_13621# clknet_4_13_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4853 a_13997_14191# tdc0.w_dly_sig\[13\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4854 a_12981_2223# a_12447_2229# a_12886_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4855 VPWR tdc0.w_dly_sig\[81\] tdc0.w_dly_sig_n\[81\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4856 tdc0.w_dly_sig_n\[103\] tdc0.w_dly_sig\[103\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4857 a_11137_15823# tdc0.o_result\[127\] a_10791_16073# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4858 a_9589_7119# a_9319_7485# a_9485_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4859 a_11060_4719# _010_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4860 VPWR _003_ a_10975_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4861 VGND tdc0.w_dly_sig_n\[44\] tdc0.w_dly_sig\[45\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4863 VGND _015_ a_14460_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4864 VPWR tdc0.w_dly_sig_n\[7\] tdc0.w_dly_sig_n\[9\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4866 VPWR tdc0.w_dly_sig\[23\] tdc0.w_dly_sig_n\[23\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4867 VPWR tdc0.w_dly_sig_n\[86\] tdc0.w_dly_sig\[87\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4868 VPWR a_16733_5461# _064_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4869 a_7047_4399# a_6265_4405# a_6963_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4870 VPWR a_14675_6549# a_14591_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4871 VGND tdc0.w_dly_sig_n\[53\] tdc0.w_dly_sig_n\[55\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4872 a_5526_15101# a_5087_14735# a_5441_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4873 _093_ a_16035_8457# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4874 a_9595_11721# _013_ a_9677_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4875 tdc0.o_result\[27\] a_16055_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4876 VPWR tdc0.o_result\[103\] a_17865_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X4877 VGND tdc0.w_dly_sig\[62\] tdc0.w_dly_sig_n\[62\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4878 a_11027_2741# a_11318_3041# a_11269_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X4879 VPWR tdc0.w_dly_sig\[26\] tdc0.w_dly_sig\[28\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4880 VPWR tdc0.w_dly_sig\[117\] tdc0.w_dly_sig_n\[117\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4881 a_5073_17999# tdc0.w_dly_sig\[20\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4882 tdc0.w_dly_sig_n\[116\] tdc0.w_dly_sig_n\[114\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4883 a_16937_1679# a_16771_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4884 VGND a_8574_4676# a_8503_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4885 a_11435_10633# _038_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4886 tdc0.o_result\[43\] a_4279_18267# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4887 tdc0.w_dly_sig_n\[5\] tdc0.w_dly_sig\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4888 a_3873_13647# a_3707_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4889 VGND a_14186_14709# a_14115_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4890 a_11872_6031# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.114 ps=1 w=0.65 l=0.15
X4891 tdc0.w_dly_sig\[22\] tdc0.w_dly_sig\[20\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4892 VGND tdc0.w_dly_sig_n\[29\] tdc0.w_dly_sig\[30\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4893 a_15473_13897# net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X4894 a_15814_18111# a_15646_18365# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4895 tdc0.w_dly_sig\[110\] tdc0.w_dly_sig_n\[109\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4896 a_9531_5095# tdc0.o_result\[69\] a_9677_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X4897 tdc0.w_dly_sig_n\[49\] tdc0.w_dly_sig\[49\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4898 a_8503_4777# a_8374_4521# a_8083_4631# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4899 VPWR a_7607_3311# a_7775_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4900 VGND a_9741_10357# _034_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X4901 VPWR a_12284_9545# uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4902 VGND net10 a_6445_16687# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X4903 VGND tdc0.w_dly_sig\[113\] tdc0.w_dly_sig_n\[113\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4904 tdc0.w_dly_sig\[66\] tdc0.w_dly_sig_n\[65\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4905 a_1945_8751# tdc0.w_dly_sig\[74\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4906 a_7182_3311# a_6743_3317# a_7097_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4907 a_15170_17429# a_15002_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4908 clknet_4_9_0_clk a_14664_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4909 a_3597_10933# a_3431_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4910 a_7258_9407# a_7090_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4911 VPWR clknet_4_8_0_clk a_12447_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4912 VGND tdc0.w_dly_sig\[70\] tdc0.w_dly_sig\[72\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4913 _022_ a_11214_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4914 a_9677_5193# _019_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X4915 tdc0.w_dly_sig_n\[92\] tdc0.w_dly_sig_n\[90\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4916 a_14676_12809# _086_ a_14510_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X4917 tdc0.w_dly_sig_n\[118\] tdc0.w_dly_sig_n\[116\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4918 VPWR a_7166_2197# a_7093_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4919 a_15906_1791# a_15738_2045# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4920 a_7917_1513# a_6927_1141# a_7791_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4921 a_2156_4777# a_1757_4405# a_2030_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4922 VGND a_11386_6652# _006_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4923 a_4498_4373# a_4330_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4924 VPWR a_9707_13077# a_9623_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
R22 VGND uio_out[5] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4926 tdc0.w_dly_sig_n\[7\] tdc0.w_dly_sig\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4927 a_6587_14013# a_5805_13647# a_6503_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4928 a_15906_1791# a_15738_2045# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4929 VPWR tdc0.w_dly_sig_n\[45\] tdc0.w_dly_sig\[46\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4930 a_8399_11721# _013_ a_8481_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4931 a_3283_17455# a_2585_17461# a_3026_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4932 VPWR _076_ a_12552_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X4933 _101_ a_6467_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4934 VPWR tdc0.o_result\[10\] a_15381_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X4935 VPWR tdc0.w_dly_sig_n\[83\] tdc0.w_dly_sig_n\[85\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4936 a_8500_4917# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4937 tdc0.w_dly_sig\[116\] tdc0.w_dly_sig_n\[115\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4938 a_6835_12809# _088_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4939 VGND tdc0.w_dly_sig\[36\] tdc0.w_dly_sig\[38\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4940 a_4295_1135# a_3431_1141# a_4038_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4941 VPWR tdc0.w_dly_sig\[42\] tdc0.w_dly_sig\[44\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4942 a_16923_14709# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4943 a_4521_6575# tdc0.w_dly_sig\[67\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4944 tdc0.w_dly_sig_n\[118\] tdc0.w_dly_sig\[118\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4945 a_14747_7663# _015_ a_14829_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4946 VPWR clknet_0_clk a_7856_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4947 a_17719_2045# a_16937_1679# a_17635_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4948 a_3502_8751# a_3229_8757# a_3417_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4949 clknet_4_4_0_clk a_3698_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4950 a_13353_5487# tdc0.w_dly_sig\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4951 a_16022_7119# net8 a_15853_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X4952 VGND a_4111_15101# a_4279_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4953 a_8481_6575# tdc0.o_result\[35\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X4954 a_6430_11989# a_6262_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4955 VPWR tdc0.w_dly_sig_n\[39\] tdc0.w_dly_sig_n\[41\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4956 tdc0.o_result\[94\] a_10259_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4957 tdc0.w_dly_sig\[34\] tdc0.w_dly_sig\[32\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4958 VPWR clknet_0_clk a_12548_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4959 a_14499_8573# a_13717_8207# a_14415_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4961 a_4146_5309# a_3873_4943# a_4061_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4962 tdc0.w_dly_sig_n\[61\] tdc0.w_dly_sig\[61\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4963 VPWR tdc0.w_dly_sig_n\[105\] tdc0.w_dly_sig\[106\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4964 a_1757_4405# a_1591_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4965 a_11058_9839# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4966 a_9374_14165# a_9206_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4967 a_2309_14197# a_2143_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4968 a_15887_15101# a_15023_14735# a_15630_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4969 a_16661_1141# a_16495_1141# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4970 a_1577_9839# tdc0.w_dly_sig\[78\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4971 VPWR tdc0.w_dly_sig_n\[55\] tdc0.w_dly_sig_n\[57\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4972 a_6262_12015# a_5989_12021# a_6177_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4973 tdc0.w_dly_sig\[51\] tdc0.w_dly_sig\[49\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4974 a_6311_12925# a_5529_12559# a_6227_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4975 VGND tdc0.w_dly_sig\[108\] tdc0.w_dly_sig\[110\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4976 _019_ a_11642_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4977 a_11023_13335# a_11119_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4978 VGND tdc0.w_dly_sig_n\[112\] tdc0.w_dly_sig_n\[114\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4980 tdc0.w_dly_sig\[100\] tdc0.w_dly_sig_n\[99\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4981 tdc0.w_dly_sig\[127\] tdc0.w_dly_sig\[125\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4982 tdc0.w_dly_sig_n\[99\] tdc0.w_dly_sig\[99\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4983 VGND tdc0.w_dly_sig_n\[57\] tdc0.w_dly_sig_n\[59\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4984 VPWR a_9282_13077# a_9209_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4985 VGND a_11159_4943# _013_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4986 VPWR tdc0.w_dly_sig_n\[52\] tdc0.w_dly_sig\[53\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4987 a_15557_15101# a_15023_14735# a_15462_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4988 a_15427_17455# a_14729_17461# a_15170_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4989 VPWR a_17406_10357# a_17335_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4990 a_17719_8359# tdc0.o_result\[103\] a_17865_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X4991 tdc0.w_dly_sig\[44\] tdc0.w_dly_sig_n\[43\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4992 a_5533_4943# tdc0.w_dly_sig\[69\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4993 VPWR a_7499_16091# a_7415_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4994 VPWR a_18027_3529# a_18034_3433# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4995 tdc0.w_dly_sig_n\[104\] tdc0.w_dly_sig\[104\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4997 a_14085_2229# a_13919_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4998 VGND a_5602_7231# a_5560_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5000 VGND clknet_4_5_0_clk a_4719_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5001 VGND ui_in[6] a_11711_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X5002 VGND a_6550_13103# clknet_4_6_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5003 _061_ a_10607_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X5004 VGND a_14899_9269# a_14906_9569# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5005 VPWR a_16819_5095# tdc0.o_result\[113\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5006 a_7093_2223# a_6559_2229# a_6998_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5007 clknet_4_10_0_clk a_16412_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5008 tdc0.w_dly_sig\[11\] tdc0.w_dly_sig_n\[10\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5009 a_14829_7983# tdc0.o_result\[99\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5010 tdc0.w_dly_sig\[52\] tdc0.w_dly_sig\[50\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5011 a_4130_15253# a_3962_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5012 a_7308_3689# a_6909_3317# a_7182_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5013 a_5713_16911# a_5547_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5014 VGND tdc0.w_dly_sig\[46\] tdc0.w_dly_sig_n\[46\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5015 VPWR clknet_4_5_0_clk a_3707_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5016 a_7331_16189# a_6633_15823# a_7074_15935# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5018 tdc0.w_dly_sig\[64\] tdc0.w_dly_sig\[62\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5019 tdc0.w_dly_sig_n\[97\] tdc0.w_dly_sig\[97\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5020 tdc0.o_result\[22\] a_16239_18267# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5021 VPWR tdc0.w_dly_sig\[38\] tdc0.w_dly_sig\[40\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5022 a_6353_1679# a_5363_1679# a_6227_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5023 VPWR tdc0.w_dly_sig\[61\] tdc0.w_dly_sig_n\[61\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5024 a_5618_5309# a_5179_4943# a_5533_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5026 VGND tdc0.o_result\[1\] a_12118_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5028 VPWR tdc0.w_dly_sig\[17\] tdc0.w_dly_sig_n\[17\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5029 tdc0.w_dly_sig\[104\] tdc0.w_dly_sig_n\[103\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5030 a_11214_7093# a_11067_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X5031 VGND tdc0.w_dly_sig\[107\] tdc0.w_dly_sig\[109\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5032 a_4498_4373# a_4330_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5033 VGND tdc0.o_result\[106\] a_14381_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5034 VGND tdc0.w_dly_sig_n\[53\] tdc0.w_dly_sig\[54\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5035 a_14952_8751# _018_ a_14786_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5036 tdc0.w_dly_sig\[101\] tdc0.w_dly_sig_n\[100\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5038 tdc0.o_result\[62\] a_7775_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5039 tdc0.o_result\[38\] a_6119_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5040 tdc0.o_result\[90\] a_7775_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5041 tdc0.w_dly_sig\[111\] tdc0.w_dly_sig_n\[110\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5042 VPWR tdc0.w_dly_sig\[28\] tdc0.w_dly_sig\[30\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5043 a_1604_11471# a_1205_11471# a_1478_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5044 VPWR tdc0.w_dly_sig\[22\] tdc0.w_dly_sig_n\[22\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5045 VGND tdc0.w_dly_sig\[113\] tdc0.w_dly_sig\[115\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5046 VPWR clknet_4_4_0_clk a_1131_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5047 a_10975_5487# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5048 VPWR a_17038_7093# a_16967_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5049 a_6909_3317# a_6743_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5050 VPWR tdc0.w_dly_sig\[94\] tdc0.w_dly_sig\[96\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5051 a_16923_14709# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5052 tdc0.w_dly_sig\[2\] net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5053 a_7883_7663# a_7185_7669# a_7626_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5054 VPWR a_1995_13103# a_2163_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5055 a_7817_17833# a_7263_17673# a_7470_17732# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X5056 a_3854_10495# a_3686_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5057 tdc0.w_dly_sig\[128\] tdc0.w_dly_sig\[126\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5058 VPWR a_11504_11445# uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5059 VPWR tdc0.w_dly_sig\[2\] tdc0.w_dly_sig\[4\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5060 VPWR a_2547_5309# a_2715_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5061 tdc0.w_dly_sig_n\[107\] tdc0.w_dly_sig_n\[105\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5062 a_4755_4399# a_4057_4405# a_4498_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5063 VGND a_1995_13103# a_2163_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5065 tdc0.o_result\[71\] a_4187_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5066 a_5639_6281# net7 a_5721_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5067 tdc0.w_dly_sig_n\[127\] tdc0.w_dly_sig_n\[125\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5068 VPWR tdc0.w_dly_sig\[88\] tdc0.w_dly_sig_n\[88\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5069 VGND tdc0.w_dly_sig\[67\] tdc0.w_dly_sig\[69\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5070 a_17935_6793# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5071 tdc0.w_dly_sig_n\[71\] tdc0.w_dly_sig_n\[69\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5072 tdc0.w_dly_sig_n\[19\] tdc0.w_dly_sig\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5074 tdc0.w_dly_sig\[12\] tdc0.w_dly_sig_n\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5075 VPWR a_17739_4631# tdc0.o_result\[114\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5076 VGND tdc0.w_dly_sig\[101\] tdc0.w_dly_sig_n\[101\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5077 a_2539_4399# a_1757_4405# a_2455_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5080 a_5529_12559# a_5363_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5081 uo_out[5] a_11456_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5082 uo_out[2] a_14676_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X5083 VPWR _019_ a_10505_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5084 a_16166_12335# tdc0.o_result\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X5085 VGND tdc0.w_dly_sig_n\[67\] tdc0.w_dly_sig\[68\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5087 VPWR a_6119_15003# a_6035_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5088 a_9482_9661# a_9209_9295# a_9397_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5089 tdc0.w_dly_sig\[7\] tdc0.w_dly_sig\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5090 VPWR tdc0.w_dly_sig_n\[66\] tdc0.w_dly_sig_n\[68\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5091 a_6191_17455# _029_ a_6273_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5092 a_13863_5487# a_12999_5493# a_13606_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5094 tdc0.w_dly_sig\[117\] tdc0.w_dly_sig\[115\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5095 a_14388_13621# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5096 a_8562_16367# a_8123_16373# a_8477_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5097 a_14783_2223# a_14085_2229# a_14526_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5098 a_14922_15797# a_14722_16097# a_15071_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5099 a_2198_17023# a_2030_17277# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5100 tdc0.w_dly_sig\[3\] tdc0.w_dly_sig_n\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5101 VPWR ui_in[5] a_12631_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5102 a_14857_9661# a_14519_9447# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5103 VGND tdc0.w_dly_sig_n\[28\] tdc0.w_dly_sig\[29\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5104 VGND tdc0.w_dly_sig\[22\] tdc0.w_dly_sig\[24\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5105 VPWR tdc0.w_dly_sig\[4\] tdc0.w_dly_sig\[6\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5106 a_12284_9545# _076_ a_12118_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5107 tdc0.w_dly_sig_n\[96\] tdc0.w_dly_sig\[96\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5108 VPWR a_11490_6005# _026_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5109 a_12210_9071# _051_ a_12376_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5110 a_17962_12381# a_17647_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5111 a_9493_2223# tdc0.o_result\[85\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5112 a_14917_15279# tdc0.w_dly_sig\[27\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5113 a_5744_4943# a_5345_4943# a_5618_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5114 tdc0.w_dly_sig\[50\] tdc0.w_dly_sig_n\[49\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5115 a_10228_8207# _001_ a_10122_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.0798 ps=0.8 w=0.42 l=0.15
X5116 a_6239_18151# a_6335_17973# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5117 VGND a_4314_13759# a_4272_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5118 VGND tdc0.w_dly_sig_n\[96\] tdc0.w_dly_sig\[97\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5119 a_9125_8457# _030_ a_9043_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X5120 VPWR tdc0.w_dly_sig\[64\] tdc0.w_dly_sig\[66\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5121 a_17651_6807# a_17935_6793# a_17870_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5122 tdc0.w_dly_sig_n\[18\] tdc0.w_dly_sig\[18\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5123 a_9839_4617# clknet_4_8_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5124 a_13353_3311# tdc0.w_dly_sig\[101\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5125 a_9779_6575# _001_ a_10029_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5126 a_7173_17999# a_6626_18273# a_6826_17973# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5127 a_8753_15823# tdc0.w_dly_sig\[38\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5129 VPWR a_17199_4917# a_17206_5217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5130 _029_ a_11122_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X5131 VPWR a_4463_1109# a_4379_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5132 VGND tdc0.w_dly_sig_n\[124\] tdc0.w_dly_sig\[125\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5133 tdc0.w_dly_sig\[53\] tdc0.w_dly_sig\[51\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5134 a_7607_9839# a_6909_9845# a_7350_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5135 VPWR tdc0.w_dly_sig\[14\] tdc0.w_dly_sig_n\[14\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5137 tdc0.w_dly_sig\[93\] tdc0.w_dly_sig_n\[92\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5138 a_15220_8751# _031_ a_14952_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5139 VPWR a_3670_8725# a_3597_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
R23 VGND uio_oe[1] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5140 VGND a_11943_17687# tdc0.o_result\[20\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5141 tdc0.w_dly_sig_n\[70\] tdc0.w_dly_sig_n\[68\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5142 VGND a_4038_10901# a_3996_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5143 _031_ a_9043_8457# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5145 VPWR a_17314_12559# clknet_4_14_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5146 VGND a_12548_14165# clknet_4_12_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5147 a_5970_1791# a_5802_2045# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5148 tdc0.w_dly_sig_n\[39\] tdc0.w_dly_sig\[39\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5149 VPWR a_4314_5055# a_4241_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5150 a_8995_7093# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5151 VGND tdc0.w_dly_sig_n\[60\] tdc0.w_dly_sig_n\[62\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5152 _001_ a_13919_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5153 a_2631_1135# a_1849_1141# a_2547_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5154 VPWR a_12518_7119# _012_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5155 a_16937_1679# a_16771_1679# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5156 a_5284_17999# a_4885_17999# a_5158_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5157 tdc0.w_dly_sig\[58\] tdc0.w_dly_sig\[56\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5158 VGND a_13311_2223# a_13479_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5159 tdc0.w_dly_sig_n\[57\] tdc0.w_dly_sig\[57\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5160 VGND a_12530_17732# a_12459_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
R24 VPWR tt_um_hpretl_tt06_tdc_17.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5161 a_1830_14847# a_1662_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5162 VGND tdc0.w_dly_sig\[30\] tdc0.w_dly_sig_n\[30\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5163 a_17651_10071# a_17942_9961# a_17893_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5164 a_15002_17455# a_14563_17461# a_14917_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5165 VGND tdc0.w_dly_sig\[103\] tdc0.w_dly_sig\[105\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5167 a_11159_4943# a_11154_5095# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=2.52 w=1 l=0.15
X5168 VPWR a_3790_7119# clknet_4_1_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5170 VGND tdc0.w_dly_sig_n\[6\] tdc0.w_dly_sig_n\[8\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5171 VPWR a_13070_8207# a_13176_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X5172 a_16741_12559# a_16187_12533# a_16394_12533# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X5173 a_14717_17999# a_14163_17973# a_14370_17973# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X5174 tdc0.w_dly_sig_n\[50\] tdc0.w_dly_sig_n\[48\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5175 a_13395_2223# a_12613_2229# a_13311_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5176 a_16823_17973# a_17114_18273# a_17065_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5177 tdc0.w_dly_sig_n\[2\] tdc0.w_dly_sig_n\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5178 a_17305_9295# a_17139_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5179 VGND tdc0.w_dly_sig\[77\] tdc0.w_dly_sig_n\[77\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5180 VPWR tdc0.o_result\[6\] a_12292_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X5181 a_18003_9661# a_17139_9295# a_17746_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5182 VPWR tdc0.w_dly_sig_n\[94\] tdc0.w_dly_sig\[95\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5184 VPWR tdc0.w_dly_sig\[41\] tdc0.w_dly_sig\[43\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5185 VPWR _023_ a_8481_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5186 VGND tdc0.w_dly_sig_n\[19\] tdc0.w_dly_sig\[20\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5187 a_15653_10383# tdc0.w_dly_sig\[4\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5188 a_12495_12247# a_12591_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5191 a_11649_6575# net4 a_11565_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5192 VGND tdc0.w_dly_sig_n\[12\] tdc0.w_dly_sig_n\[14\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5193 a_5349_7119# tdc0.w_dly_sig\[65\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5194 VPWR clknet_4_8_0_clk a_10975_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5195 a_11619_8867# _075_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X5196 VGND a_5786_5055# a_5744_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5197 VPWR tdc0.w_dly_sig\[40\] tdc0.w_dly_sig_n\[40\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5198 a_3873_4943# a_3707_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5199 a_5157_6953# a_4167_6581# a_5031_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5200 VPWR a_10515_7671# _000_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5201 VGND tdc0.w_dly_sig\[7\] a_14349_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5202 a_12323_17673# clknet_4_13_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5203 a_14299_17999# a_14163_17973# a_13879_17973# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5204 VGND tdc0.w_dly_sig\[32\] tdc0.w_dly_sig_n\[32\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5205 VGND _001_ a_13690_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5206 clknet_4_12_0_clk a_12548_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5207 a_9665_13481# a_8675_13109# a_9539_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5209 tdc0.w_dly_sig\[9\] tdc0.w_dly_sig\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5210 tdc0.w_dly_sig\[114\] tdc0.w_dly_sig\[112\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5211 a_4241_5309# a_3707_4943# a_4146_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5212 VPWR tdc0.w_dly_sig_n\[114\] tdc0.w_dly_sig\[115\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5213 a_8914_17429# a_8746_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5214 tdc0.w_dly_sig\[50\] tdc0.w_dly_sig\[48\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5215 VPWR a_11214_7093# _022_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X5216 VPWR tdc0.o_result\[54\] a_5997_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X5218 clknet_4_15_0_clk a_16578_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5219 VPWR tdc0.w_dly_sig\[48\] tdc0.w_dly_sig_n\[48\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5220 a_6411_17277# a_5547_16911# a_6154_17023# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5221 VGND a_6154_17023# a_6112_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5222 VGND tdc0.o_result\[119\] a_18153_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5223 a_15903_12533# a_16194_12833# a_16145_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5224 VPWR a_10759_8181# _005_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5225 tdc0.w_dly_sig_n\[95\] tdc0.w_dly_sig\[95\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5226 VGND tdc0.w_dly_sig\[15\] tdc0.w_dly_sig\[17\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5227 VPWR _008_ a_14445_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
R25 VPWR tt_um_hpretl_tt06_tdc_23.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5228 a_15465_10383# a_15299_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5229 VPWR tdc0.w_dly_sig\[47\] tdc0.w_dly_sig\[49\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5230 VPWR tdc0.w_dly_sig\[103\] tdc0.w_dly_sig_n\[103\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5231 a_6081_17277# a_5547_16911# a_5986_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5232 tdc0.o_result\[89\] a_7591_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5233 VPWR tdc0.w_dly_sig\[71\] tdc0.w_dly_sig\[73\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5234 VPWR tdc0.w_dly_sig_n\[42\] tdc0.w_dly_sig_n\[44\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5235 VPWR tdc0.w_dly_sig\[77\] tdc0.w_dly_sig\[79\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5236 tdc0.w_dly_sig\[60\] tdc0.w_dly_sig_n\[59\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5237 a_17893_6575# a_17555_6807# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5238 a_12867_11159# a_13158_11049# a_13109_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5239 VGND tdc0.w_dly_sig\[127\] a_17661_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5240 a_16766_7119# a_16451_7271# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5242 tdc0.w_dly_sig_n\[97\] tdc0.w_dly_sig_n\[95\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5243 tdc0.w_dly_sig\[65\] tdc0.w_dly_sig\[63\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5244 tdc0.w_dly_sig\[125\] tdc0.w_dly_sig\[123\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5245 VGND a_2566_3285# a_2524_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5246 a_2198_8725# a_2030_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5247 VPWR a_17774_2741# a_17703_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5248 VGND a_13979_3829# a_13986_4129# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5249 tdc0.w_dly_sig\[75\] tdc0.w_dly_sig_n\[74\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5250 a_9677_11721# tdc0.o_result\[61\] a_9595_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5251 VGND a_15887_15101# a_16055_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5252 a_11154_5095# net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5253 tdc0.w_dly_sig_n\[62\] tdc0.w_dly_sig\[62\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5254 a_7699_6397# a_7001_6031# a_7442_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5255 VGND tdc0.w_dly_sig_n\[24\] tdc0.w_dly_sig_n\[26\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5256 tdc0.w_dly_sig\[93\] tdc0.w_dly_sig\[91\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5257 a_13151_11145# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5258 a_13908_4943# tdc0.o_result\[105\] a_13605_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X5259 VPWR a_9650_9407# a_9577_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5260 VGND clknet_4_5_0_clk a_3707_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5261 a_3877_15279# tdc0.w_dly_sig\[45\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5262 a_4195_15101# a_3413_14735# a_4111_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5263 tdc0.w_dly_sig_n\[21\] tdc0.w_dly_sig\[21\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5264 VPWR tdc0.w_dly_sig_n\[34\] tdc0.w_dly_sig\[35\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5265 _088_ a_6191_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5267 a_5997_13423# _022_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X5268 VPWR tdc0.w_dly_sig\[63\] tdc0.w_dly_sig_n\[63\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5269 VPWR a_11058_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5270 tdc0.w_dly_sig\[88\] tdc0.w_dly_sig\[86\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5271 a_6906_16189# a_6633_15823# a_6821_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5273 a_11119_13335# a_11410_13225# a_11361_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5274 tdc0.w_dly_sig\[124\] tdc0.w_dly_sig\[122\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5275 a_2198_8725# a_2030_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5277 a_7013_12809# _089_ a_6917_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X5278 a_6549_10633# _100_ a_6467_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X5279 a_17669_9129# a_16679_8757# a_17543_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5280 a_7281_1135# tdc0.w_dly_sig\[92\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5281 VPWR a_9807_17687# _032_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X5282 VGND tdc0.w_dly_sig\[17\] tdc0.w_dly_sig\[19\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5283 VPWR a_9650_7637# _025_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.135 ps=1.27 w=1 l=0.15
X5284 VPWR clknet_0_clk a_12548_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5285 a_15093_7983# tdc0.o_result\[11\] a_14747_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5286 VGND _000_ _016_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5287 clknet_4_1_0_clk a_3790_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5288 a_3790_7119# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X5289 VPWR tdc0.w_dly_sig\[94\] tdc0.w_dly_sig_n\[94\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5291 a_10585_12335# tdc0.o_result\[15\] a_10239_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5292 tdc0.w_dly_sig_n\[110\] tdc0.w_dly_sig_n\[108\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5293 a_6269_6575# tdc0.w_dly_sig\[59\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5294 clknet_4_4_0_clk a_3698_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5295 VGND a_16923_14709# a_16930_15009# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5296 VPWR a_6154_17023# a_6081_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5297 a_9029_13103# tdc0.w_dly_sig\[32\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5298 VPWR a_12548_14165# clknet_4_12_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5300 _009_ a_11938_8253# a_12297_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.52 pd=3.04 as=0.135 ps=1.27 w=1 l=0.15
X5301 a_9025_17999# a_8859_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5302 VGND tdc0.w_dly_sig\[113\] a_18581_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5303 tdc0.w_dly_sig_n\[73\] tdc0.w_dly_sig\[73\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5304 a_7825_13423# tdc0.o_result\[52\] a_7479_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5305 a_11422_5487# _002_ a_11225_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5306 tdc0.w_dly_sig_n\[60\] tdc0.w_dly_sig\[60\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5308 a_14335_14735# a_14115_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X5309 a_13717_8207# a_13551_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5310 clknet_4_15_0_clk a_16578_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5311 VGND tdc0.w_dly_sig\[124\] tdc0.w_dly_sig_n\[124\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5312 a_13805_9071# tdc0.o_result\[20\] a_13459_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5314 VPWR _010_ a_9493_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5315 VGND tdc0.w_dly_sig\[39\] tdc0.w_dly_sig\[41\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5316 a_7967_7663# a_7185_7669# a_7883_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5317 VPWR clknet_4_5_0_clk a_3523_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5318 a_8017_10927# tdc0.w_dly_sig\[62\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5319 a_6227_12925# a_5363_12559# a_5970_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5320 VPWR a_11023_13335# tdc0.o_result\[13\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5321 VPWR tdc0.w_dly_sig\[114\] tdc0.w_dly_sig_n\[114\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5322 a_2122_5309# a_1849_4943# a_2037_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5323 a_17743_3543# a_18027_3529# a_17962_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5324 a_13979_14709# clknet_4_13_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5325 VGND tdc0.w_dly_sig_n\[73\] tdc0.w_dly_sig_n\[75\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5326 VPWR a_16819_10535# tdc0.o_result\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5327 tdc0.w_dly_sig_n\[113\] tdc0.w_dly_sig_n\[111\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5328 a_10505_4943# tdc0.o_result\[111\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5329 VPWR a_7515_9661# a_7683_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5330 a_17774_17732# a_17574_17577# a_17923_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5331 a_17463_14423# a_17559_14423# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5332 VPWR tdc0.w_dly_sig_n\[33\] tdc0.w_dly_sig_n\[35\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5333 VPWR a_17187_16599# tdc0.o_result\[125\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5334 VPWR a_13979_3829# a_13986_4129# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5335 VGND clknet_4_2_0_clk a_6559_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5336 VPWR tdc0.w_dly_sig_n\[103\] tdc0.w_dly_sig_n\[105\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5337 a_14949_13103# a_14611_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5338 VGND tdc0.w_dly_sig_n\[116\] tdc0.w_dly_sig\[117\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5339 _087_ a_5639_6281# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5340 _025_ a_9650_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5341 a_4057_4405# a_3891_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5342 tdc0.w_dly_sig\[19\] tdc0.w_dly_sig_n\[18\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5343 a_10759_8181# _004_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X5344 tdc0.o_result\[80\] a_2991_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5345 a_7093_1141# a_6927_1141# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5346 a_16762_8207# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5347 VGND tdc0.w_dly_sig_n\[4\] tdc0.w_dly_sig_n\[6\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5348 a_8270_10901# a_8102_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5349 VPWR a_2455_8751# a_2623_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5350 a_17761_1679# a_16771_1679# a_17635_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5351 a_16951_5487# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5352 a_9125_8751# tdc0.o_result\[89\] a_9043_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5353 a_8473_17461# a_8307_17461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5354 VGND clknet_4_5_0_clk a_5547_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5355 a_6614_8319# a_6446_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5356 VGND a_6883_17687# tdc0.o_result\[16\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5357 VPWR tdc0.w_dly_sig_n\[127\] tdc0.w_dly_sig\[128\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5358 tdc0.w_dly_sig\[29\] tdc0.w_dly_sig\[27\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5359 tdc0.w_dly_sig_n\[46\] tdc0.w_dly_sig\[46\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5360 a_6177_12015# tdc0.w_dly_sig\[58\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5361 VPWR a_3451_17429# a_3367_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5362 _055_ a_10423_5193# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5363 a_6614_8319# a_6446_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5364 tdc0.o_result\[70\] a_4095_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5365 VPWR a_16071_18365# a_16239_18267# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5366 a_5157_17833# a_4167_17461# a_5031_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5367 a_17286_8725# a_17118_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5368 VPWR clknet_4_4_0_clk a_4259_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5369 a_3996_11305# a_3597_10933# a_3870_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5370 tdc0.w_dly_sig\[41\] tdc0.w_dly_sig_n\[40\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5371 a_14899_9269# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5372 a_11149_9545# tdc0.o_result\[62\] a_11067_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5373 VGND tdc0.w_dly_sig_n\[28\] tdc0.w_dly_sig_n\[30\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5374 a_5533_4943# tdc0.w_dly_sig\[69\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5375 VGND a_7470_17732# a_7399_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X5376 _049_ a_10239_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5377 a_16301_6281# _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X5378 VGND a_9839_4617# a_9846_4521# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5379 VPWR a_9459_4631# tdc0.o_result\[111\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5380 VPWR a_5123_13103# a_5291_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5381 tdc0.w_dly_sig\[69\] tdc0.w_dly_sig_n\[68\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5382 tdc0.w_dly_sig\[11\] tdc0.w_dly_sig\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5383 VPWR tdc0.o_result\[122\] a_16301_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X5384 VPWR a_5951_15101# a_6119_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5385 VPWR a_6550_13103# clknet_4_6_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5386 VGND a_8730_16341# a_8688_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5387 VGND tdc0.w_dly_sig\[69\] tdc0.w_dly_sig_n\[69\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5389 VGND clknet_4_5_0_clk a_2419_17461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5390 tdc0.w_dly_sig\[81\] tdc0.w_dly_sig\[79\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5391 VGND a_5123_13103# a_5291_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5392 VGND tdc0.w_dly_sig\[46\] tdc0.w_dly_sig\[48\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5393 VGND tdc0.w_dly_sig_n\[30\] tdc0.w_dly_sig_n\[32\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5394 _079_ a_9043_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5395 VGND a_3854_10495# a_3812_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5396 tdc0.w_dly_sig_n\[105\] tdc0.w_dly_sig_n\[103\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5397 VPWR tdc0.w_dly_sig\[60\] tdc0.w_dly_sig\[62\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5398 VPWR a_16923_14709# a_16930_15009# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5399 VPWR a_6119_4123# a_6035_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5400 VGND ui_in[0] a_18187_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5402 tdc0.o_result\[47\] a_2623_17179# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5403 VPWR tdc0.w_dly_sig\[98\] tdc0.w_dly_sig_n\[98\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5405 tdc0.w_dly_sig\[52\] tdc0.w_dly_sig_n\[51\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5406 VGND a_17463_14423# tdc0.o_result\[122\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5407 a_3762_5461# a_3594_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5408 a_4521_17455# tdc0.w_dly_sig\[43\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5409 a_11490_6005# a_12148_6005# a_12082_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X5411 tdc0.o_result\[34\] a_8051_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5412 a_11610_12292# a_11410_12137# a_11759_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5413 VPWR tdc0.w_dly_sig_n\[47\] tdc0.w_dly_sig_n\[49\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5414 tdc0.w_dly_sig_n\[73\] tdc0.w_dly_sig_n\[71\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5415 VGND tdc0.o_result\[5\] a_11290_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5416 VPWR net4 a_11122_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X5417 a_16934_1135# a_16661_1141# a_16849_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5419 VGND a_18050_14468# a_17979_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X5420 VGND clknet_4_5_0_clk a_1591_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5421 clknet_4_14_0_clk a_17314_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5422 a_9301_14191# a_8767_14197# a_9206_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5423 VGND ui_in[4] a_10423_591# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5424 a_13979_14709# clknet_4_13_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5425 VGND tdc0.w_dly_sig_n\[27\] tdc0.w_dly_sig\[28\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5426 VGND a_11456_10927# uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5428 a_2313_3311# tdc0.w_dly_sig\[81\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5429 clknet_4_8_0_clk a_12548_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5430 VGND clknet_4_13_0_clk a_14563_17461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5431 VGND _005_ a_16166_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5432 VGND clknet_4_8_0_clk a_10975_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5433 a_7263_17673# clknet_4_7_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5434 VPWR tdc0.w_dly_sig\[80\] tdc0.w_dly_sig_n\[80\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5435 a_18121_17833# a_17574_17577# a_17774_17732# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5436 clknet_4_8_0_clk a_12548_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5437 tdc0.w_dly_sig\[31\] tdc0.w_dly_sig_n\[30\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5438 VPWR tdc0.w_dly_sig_n\[40\] tdc0.w_dly_sig\[41\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5440 a_7458_7663# a_7019_7669# a_7373_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5441 tdc0.w_dly_sig_n\[18\] tdc0.w_dly_sig_n\[16\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5442 a_10226_6575# a_10446_6549# _023_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5443 VGND tdc0.w_dly_sig\[25\] tdc0.w_dly_sig_n\[25\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5445 VGND tdc0.w_dly_sig\[3\] a_15545_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5447 a_11290_11247# tdc0.o_result\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X5448 VGND tdc0.w_dly_sig_n\[10\] tdc0.w_dly_sig_n\[12\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5449 VPWR a_6855_11989# a_6771_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5450 a_16155_17687# tdc0.o_result\[22\] a_16301_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5451 a_4330_4399# a_3891_4405# a_4245_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5452 net1 a_18187_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5453 VGND tdc0.w_dly_sig_n\[1\] tdc0.w_dly_sig_n\[3\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5454 a_9975_4777# a_9846_4521# a_9555_4631# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5455 a_6503_14013# a_5805_13647# a_6246_13759# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5456 a_14650_15823# a_14335_15975# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5457 VGND clknet_0_clk a_3348_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5458 tdc0.w_dly_sig\[29\] tdc0.w_dly_sig_n\[28\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5459 a_10137_2223# tdc0.o_result\[95\] a_10055_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5460 VPWR a_17543_8751# a_17711_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5461 VPWR a_15170_17429# a_15097_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5462 VPWR clknet_0_clk a_14664_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5463 a_15419_7895# tdc0.o_result\[118\] a_15565_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5464 tdc0.w_dly_sig\[82\] tdc0.w_dly_sig_n\[81\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5465 a_8941_6281# tdc0.o_result\[108\] a_8859_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5466 a_17157_5309# a_16819_5095# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5467 VGND a_14664_6005# clknet_4_9_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5468 VGND a_7515_9661# a_7683_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5469 a_2566_3285# a_2398_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5470 a_4606_6575# a_4333_6581# a_4521_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5471 a_10239_10633# _026_ a_10321_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5472 a_7074_15935# a_6906_16189# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5473 VPWR a_15427_15279# a_15595_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5474 VPWR _002_ a_11343_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X5475 VGND tdc0.w_dly_sig_n\[17\] tdc0.w_dly_sig_n\[19\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5477 VPWR tdc0.w_dly_sig\[99\] tdc0.w_dly_sig_n\[99\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5478 clknet_4_4_0_clk a_3698_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5479 VGND a_15427_15279# a_15595_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5480 VPWR tdc0.w_dly_sig\[110\] tdc0.w_dly_sig_n\[110\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5481 VPWR tdc0.w_dly_sig\[89\] tdc0.w_dly_sig_n\[89\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5482 a_1205_11471# a_1039_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5483 VGND a_7856_14165# clknet_4_7_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5485 VGND tdc0.w_dly_sig_n\[36\] tdc0.w_dly_sig\[37\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5486 VPWR a_16332_12015# uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5487 tdc0.o_result\[88\] a_7131_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5488 VPWR a_15419_7895# _045_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X5489 a_11251_15279# _029_ a_11333_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5490 a_17378_1791# a_17210_2045# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5491 a_2087_9839# a_1389_9845# a_1830_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5492 VGND a_12548_14165# clknet_4_12_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5493 a_1938_10927# a_1665_10933# a_1853_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5494 VGND clknet_0_clk a_8500_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5495 a_16547_7093# a_16831_7093# a_16766_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5496 VGND clknet_4_4_0_clk a_1499_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5497 VGND _016_ a_12171_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X5498 a_12069_10633# _045_ a_11987_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X5499 VPWR tdc0.w_dly_sig_n\[92\] tdc0.w_dly_sig_n\[94\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5500 VPWR a_4295_10927# a_4463_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5502 a_11403_13321# clknet_4_12_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5503 VPWR tdc0.w_dly_sig\[53\] tdc0.w_dly_sig\[55\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5504 VPWR clknet_0_clk a_14388_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5505 tdc0.w_dly_sig\[109\] tdc0.w_dly_sig_n\[108\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5506 a_14358_2223# a_13919_2229# a_14273_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5507 a_2823_3311# a_2125_3317# a_2566_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5508 VPWR tdc0.w_dly_sig_n\[41\] tdc0.w_dly_sig\[42\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5509 a_9669_9955# _079_ a_9597_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5510 _019_ _002_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5511 VGND a_9431_1109# a_9389_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5512 tdc0.w_dly_sig_n\[84\] tdc0.w_dly_sig_n\[82\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5513 tdc0.w_dly_sig_n\[48\] tdc0.w_dly_sig\[48\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5514 _023_ a_10446_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5515 a_11214_7093# a_11872_7093# a_11806_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X5516 a_4571_14013# a_3707_13647# a_4314_13759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5517 a_17703_13647# a_17567_13621# a_17283_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5518 a_16589_17775# net9 a_16155_17687# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5519 a_18383_3677# a_18163_3689# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X5520 VGND tdc0.w_dly_sig_n\[4\] tdc0.w_dly_sig\[5\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5521 a_8565_15823# a_8399_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5522 VGND tdc0.w_dly_sig\[2\] tdc0.w_dly_sig_n\[2\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5523 a_15903_12533# a_16187_12533# a_16122_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5524 VPWR _087_ a_7085_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5525 a_6979_17687# a_7270_17577# a_7221_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5526 _077_ a_4535_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5527 tdc0.w_dly_sig\[66\] tdc0.w_dly_sig\[64\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5528 VPWR a_9374_14165# a_9301_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5529 VGND a_7607_3311# a_7775_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5530 VPWR clk a_11058_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5533 a_4333_17461# a_4167_17461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5534 a_14115_3855# a_13986_4129# a_13695_3829# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5535 VPWR a_2290_5055# a_2217_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5536 a_15235_5719# tdc0.o_result\[10\] a_15381_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X5537 a_6357_10933# a_6191_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5538 tdc0.w_dly_sig_n\[77\] tdc0.w_dly_sig\[77\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5539 a_4241_14013# a_3707_13647# a_4146_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5540 tdc0.w_dly_sig_n\[44\] tdc0.w_dly_sig_n\[42\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5541 a_8201_12015# tdc0.w_dly_sig\[64\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5542 VGND tdc0.w_dly_sig\[35\] tdc0.w_dly_sig_n\[35\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5543 VGND tdc0.w_dly_sig_n\[110\] tdc0.w_dly_sig_n\[112\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5544 VPWR tdc0.w_dly_sig_n\[76\] tdc0.w_dly_sig\[77\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5545 VGND a_9466_18111# a_9424_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5546 a_11609_4399# tdc0.o_result\[102\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5547 VGND _078_ a_9366_10071# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5548 VGND tdc0.w_dly_sig_n\[38\] tdc0.w_dly_sig_n\[40\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5550 a_18318_9839# a_18071_10217# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5551 tdc0.w_dly_sig_n\[3\] tdc0.w_dly_sig\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5552 a_14563_5487# _015_ a_14645_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5553 VPWR tdc0.w_dly_sig\[63\] tdc0.w_dly_sig\[65\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5554 tdc0.w_dly_sig\[126\] tdc0.w_dly_sig_n\[125\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5555 VPWR tdc0.w_dly_sig_n\[1\] tdc0.w_dly_sig\[2\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5556 a_6445_16687# tdc0.o_result\[19\] a_6099_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5557 a_7584_8041# a_7185_7669# a_7458_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5559 a_11596_7119# net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.114 ps=1 w=0.65 l=0.15
X5560 VGND a_11610_12292# a_11539_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X5561 tdc0.w_dly_sig_n\[88\] tdc0.w_dly_sig\[88\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5562 tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5563 VPWR tdc0.w_dly_sig\[112\] tdc0.w_dly_sig_n\[112\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5564 tdc0.w_dly_sig\[86\] tdc0.w_dly_sig\[84\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5565 VGND a_9834_3285# a_9792_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5566 VGND tdc0.w_dly_sig_n\[105\] tdc0.w_dly_sig_n\[107\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5567 a_4456_4777# a_4057_4405# a_4330_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5568 a_9631_4221# a_8933_3855# a_9374_3967# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5569 tdc0.w_dly_sig\[43\] tdc0.w_dly_sig\[41\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5570 a_10239_8751# _028_ a_10321_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5572 tdc0.w_dly_sig\[74\] tdc0.w_dly_sig_n\[73\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5573 VPWR a_9747_8181# _007_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.62 as=0.165 ps=1.33 w=1 l=0.15
X5574 a_14519_9447# a_14615_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5575 VGND a_5751_18267# a_5709_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5576 tdc0.o_result\[99\] a_14491_1109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5577 VPWR a_16412_6549# clknet_4_10_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5578 tdc0.w_dly_sig\[68\] tdc0.w_dly_sig_n\[67\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5579 tdc0.w_dly_sig_n\[14\] tdc0.w_dly_sig_n\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5580 a_6467_7369# net7 a_6549_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5581 a_4295_10927# a_3431_10933# a_4038_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5582 a_4617_8751# tdc0.o_result\[49\] a_4535_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5583 a_14510_12559# tdc0.o_result\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X5584 VPWR a_8051_7637# a_7967_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5585 tdc0.w_dly_sig_n\[40\] tdc0.w_dly_sig\[40\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5586 a_9043_8751# _028_ a_9125_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5587 tdc0.w_dly_sig\[108\] tdc0.w_dly_sig_n\[107\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5588 VGND tdc0.w_dly_sig_n\[3\] tdc0.w_dly_sig\[4\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5589 VGND tdc0.w_dly_sig_n\[40\] tdc0.w_dly_sig_n\[42\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5590 a_17036_5807# tdc0.o_result\[112\] a_16733_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X5591 VPWR tdc0.w_dly_sig_n\[12\] tdc0.w_dly_sig\[13\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5592 VPWR a_12323_17673# a_12330_17577# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5593 tdc0.o_result\[85\] a_4923_1947# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5595 VPWR a_13863_3311# a_14031_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5596 tdc0.w_dly_sig_n\[85\] tdc0.w_dly_sig\[85\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5598 a_13717_8207# a_13551_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5599 _062_ a_8491_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5600 clknet_4_15_0_clk a_16578_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5601 VGND a_14675_6549# a_14633_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5602 a_6246_13759# a_6078_14013# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5603 a_2156_16911# a_1757_16911# a_2030_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5604 a_16819_5095# a_16915_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5606 a_9482_2045# a_9209_1679# a_9397_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5607 a_2511_10633# _026_ a_2593_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5608 a_14952_8751# _005_ a_14868_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5609 tdc0.w_dly_sig\[47\] tdc0.w_dly_sig_n\[46\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5610 VPWR a_17567_16585# a_17574_16489# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5611 VGND clknet_4_6_0_clk a_6743_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5612 a_8838_16189# a_8399_15823# a_8753_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5613 a_14484_2601# a_14085_2229# a_14358_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5614 a_9125_6895# tdc0.o_result\[76\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5615 VGND a_7699_4221# a_7867_4123# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5616 a_5639_6281# net7 a_5721_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5617 VPWR tdc0.w_dly_sig\[13\] tdc0.w_dly_sig_n\[13\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5618 VGND _021_ a_9043_8457# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5619 clknet_4_7_0_clk a_7856_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5620 a_15630_14847# a_15462_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5621 a_4697_4943# a_3707_4943# a_4571_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5622 tdc0.w_dly_sig\[17\] tdc0.w_dly_sig\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5623 VPWR tdc0.w_dly_sig\[111\] a_18121_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5624 a_8573_5487# tdc0.o_result\[88\] a_8491_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5625 a_8653_11305# a_7663_10933# a_8527_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5626 a_11403_12233# clknet_4_12_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5628 tdc0.w_dly_sig\[49\] tdc0.w_dly_sig\[47\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5629 VGND tdc0.o_result\[38\] a_6285_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5630 VPWR a_4314_13759# a_4241_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5631 VPWR tdc0.w_dly_sig_n\[97\] tdc0.w_dly_sig\[98\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5632 a_3854_18111# a_3686_18365# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5633 a_7626_5461# a_7458_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5634 tdc0.w_dly_sig\[103\] tdc0.w_dly_sig_n\[102\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5635 VGND tdc0.w_dly_sig\[9\] tdc0.w_dly_sig_n\[9\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5636 VGND tdc0.w_dly_sig_n\[93\] tdc0.w_dly_sig_n\[95\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5637 a_8178_8725# a_8010_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5638 VGND a_5199_17429# a_5157_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5639 tdc0.w_dly_sig_n\[60\] tdc0.w_dly_sig_n\[58\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5640 clknet_4_9_0_clk a_14664_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X5641 tdc0.w_dly_sig_n\[15\] tdc0.w_dly_sig_n\[13\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5642 VPWR tdc0.w_dly_sig\[90\] tdc0.w_dly_sig\[92\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5643 tdc0.w_dly_sig\[53\] tdc0.w_dly_sig_n\[52\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5644 a_6354_6575# a_5915_6581# a_6269_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5646 _013_ a_11159_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5647 _065_ a_14563_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5648 a_14195_8867# _017_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X5649 a_11965_1679# a_10975_1679# a_11839_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5650 a_17029_1135# a_16495_1141# a_16934_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5651 VPWR tdc0.o_result\[24\] a_16301_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X5652 a_8745_8207# tdc0.o_result\[92\] a_8399_8457# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5653 VGND tdc0.w_dly_sig\[127\] tdc0.w_dly_sig\[129\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5654 VGND tdc0.w_dly_sig_n\[92\] tdc0.w_dly_sig\[93\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5655 a_11892_11471# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5656 _027_ a_9043_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5657 VGND a_14952_8751# uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5658 VGND a_17647_3543# tdc0.o_result\[112\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5659 VPWR a_12792_6549# a_12134_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=2.12 as=0.165 ps=1.33 w=1 l=0.15
X5660 tdc0.w_dly_sig\[105\] tdc0.w_dly_sig\[103\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5661 VPWR _062_ a_15825_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5663 VPWR a_3175_14165# a_3091_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5664 VPWR tdc0.w_dly_sig\[36\] tdc0.w_dly_sig_n\[36\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5665 VPWR tdc0.w_dly_sig\[33\] tdc0.w_dly_sig\[35\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5666 VGND tdc0.w_dly_sig\[1\] a_16741_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5667 tdc0.w_dly_sig\[21\] tdc0.w_dly_sig_n\[20\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5668 VGND tdc0.w_dly_sig\[24\] a_14717_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5669 a_7607_9839# a_6743_9845# a_7350_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5670 VPWR tdc0.w_dly_sig\[29\] tdc0.w_dly_sig\[31\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5671 a_6154_17023# a_5986_17277# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5672 a_2087_15101# a_1389_14735# a_1830_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5673 a_13438_3311# a_13165_3317# a_13353_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5674 a_17335_4943# a_17199_4917# a_16915_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5675 _100_ a_2511_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5676 VPWR a_4038_10901# a_3965_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5677 a_8178_8725# a_8010_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5678 VGND tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5679 VGND tdc0.w_dly_sig_n\[99\] tdc0.w_dly_sig_n\[101\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5680 a_17559_14423# a_17850_14313# a_17801_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5681 VGND tdc0.w_dly_sig\[68\] tdc0.w_dly_sig_n\[68\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5682 a_6239_18151# a_6335_17973# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5683 VPWR a_4774_6549# a_4701_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5684 a_15738_10749# a_15299_10383# a_15653_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5685 VGND tdc0.w_dly_sig_n\[5\] tdc0.w_dly_sig_n\[7\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5686 tdc0.o_result\[29\] a_9799_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5687 a_2582_14191# a_2143_14197# a_2497_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5688 _044_ a_11146_4719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5689 VGND tdc0.w_dly_sig_n\[11\] tdc0.w_dly_sig\[12\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5690 tdc0.w_dly_sig\[98\] tdc0.w_dly_sig_n\[97\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5691 a_11714_7983# a_10975_7663# a_11600_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.137 ps=1.07 w=0.65 l=0.15
X5692 a_18027_12233# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5693 a_11361_14191# a_11023_14423# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5694 a_12134_6549# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.175 ps=1.35 w=1 l=0.15
X5695 a_12483_4221# a_11785_3855# a_12226_3967# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5696 tdc0.w_dly_sig\[79\] tdc0.w_dly_sig_n\[78\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5698 tdc0.w_dly_sig\[92\] tdc0.w_dly_sig\[90\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5699 tdc0.w_dly_sig\[103\] tdc0.w_dly_sig\[101\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5700 VGND a_8819_7637# net6 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5701 tdc0.w_dly_sig\[90\] tdc0.w_dly_sig\[88\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5702 tdc0.o_result\[78\] a_2623_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5703 a_8838_16189# a_8565_15823# a_8753_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5704 tdc0.w_dly_sig\[67\] tdc0.w_dly_sig\[65\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5705 VPWR a_11518_2741# a_11447_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5706 a_6361_8207# tdc0.w_dly_sig\[66\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5707 VPWR tdc0.o_result\[53\] a_9959_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5708 tdc0.o_result\[81\] a_2715_3035# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5709 tdc0.o_result\[41\] a_7499_16091# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5710 tdc0.w_dly_sig\[116\] tdc0.w_dly_sig\[114\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5711 a_16789_7485# a_16451_7271# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5712 a_4839_4399# a_4057_4405# a_4755_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5713 VGND a_2715_3035# a_2673_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5714 VPWR tdc0.w_dly_sig\[118\] tdc0.w_dly_sig\[120\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5716 tdc0.w_dly_sig_n\[124\] tdc0.w_dly_sig\[124\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5718 a_13937_4221# a_13599_4007# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5719 VPWR a_10259_3285# a_10175_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5720 tdc0.o_result\[85\] a_4923_1947# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5721 tdc0.w_dly_sig_n\[115\] tdc0.w_dly_sig_n\[113\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5722 _066_ a_15575_6281# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X5723 a_13165_3317# a_12999_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5724 _030_ a_8399_8457# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5725 a_5087_9545# _029_ a_5169_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5726 VGND a_7626_5461# a_7584_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5727 a_16301_14191# _007_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X5728 a_6480_6953# a_6081_6581# a_6354_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5729 a_4755_2045# a_4057_1679# a_4498_1791# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5730 VGND tdc0.w_dly_sig\[6\] tdc0.w_dly_sig\[8\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5731 a_1945_16911# tdc0.w_dly_sig\[48\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5732 VPWR a_17463_14423# tdc0.o_result\[122\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5733 a_12376_8751# _005_ a_12292_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5734 VGND a_16332_9839# uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5735 a_5970_12671# a_5802_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5736 a_18489_10217# a_17942_9961# a_18142_10116# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5737 a_11780_7637# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.312 ps=2.12 w=0.42 l=0.15
X5738 a_15561_17999# tdc0.w_dly_sig\[23\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5739 VPWR tdc0.w_dly_sig\[28\] tdc0.w_dly_sig_n\[28\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5740 VGND a_3790_7119# clknet_4_1_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5741 tdc0.o_result\[43\] a_4279_18267# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5742 VPWR a_9339_17429# a_9255_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5743 a_16155_6183# tdc0.o_result\[24\] a_16301_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X5745 a_2566_3285# a_2398_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5746 a_11943_17687# a_12039_17687# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5747 tdc0.w_dly_sig\[100\] tdc0.w_dly_sig\[98\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5748 VGND a_17314_12559# clknet_4_14_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5749 _059_ a_10791_16073# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5750 a_4701_6575# a_4167_6581# a_4606_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5751 a_4130_15253# a_3962_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5752 a_14867_2223# a_14085_2229# a_14783_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5753 VGND tdc0.w_dly_sig_n\[33\] tdc0.w_dly_sig\[34\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5754 a_3409_17833# a_2419_17461# a_3283_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5755 clknet_0_clk a_11058_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5756 tdc0.o_result\[75\] a_2071_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5757 VPWR a_8435_8751# a_8603_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5758 tdc0.w_dly_sig_n\[109\] tdc0.w_dly_sig\[109\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5759 a_6813_12393# a_5823_12021# a_6687_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5760 a_9217_5807# tdc0.o_result\[90\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5761 a_11597_8207# tdc0.o_result\[121\] a_11251_8457# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5762 tdc0.w_dly_sig\[15\] tdc0.w_dly_sig\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5763 VGND tdc0.w_dly_sig_n\[80\] tdc0.w_dly_sig\[81\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5764 VGND tdc0.w_dly_sig\[85\] tdc0.w_dly_sig\[87\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5765 VGND clknet_4_7_0_clk a_8307_17461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5766 tdc0.w_dly_sig\[128\] tdc0.w_dly_sig_n\[127\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5767 a_8477_16367# tdc0.w_dly_sig\[40\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5769 a_7274_4221# a_7001_3855# a_7189_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5770 VPWR tdc0.w_dly_sig\[24\] tdc0.w_dly_sig_n\[24\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5771 a_17187_16599# a_17283_16599# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5772 a_9581_3311# tdc0.w_dly_sig\[95\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5773 a_11582_1791# a_11414_2045# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5774 VGND a_18187_10901# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5775 tdc0.w_dly_sig_n\[0\] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5776 VPWR tdc0.w_dly_sig\[30\] tdc0.w_dly_sig\[32\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5777 a_16163_10749# a_15299_10383# a_15906_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5778 VPWR a_11214_7093# _022_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5779 VGND tdc0.w_dly_sig\[91\] tdc0.w_dly_sig\[93\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5780 VPWR clknet_4_6_0_clk a_7663_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5782 uo_out[1] a_12284_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5783 a_4535_8751# _022_ a_4617_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5784 a_11973_3855# tdc0.w_dly_sig\[106\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5785 tdc0.w_dly_sig\[37\] tdc0.w_dly_sig\[35\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5786 VGND a_2014_6549# a_1972_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5787 tdc0.w_dly_sig_n\[71\] tdc0.w_dly_sig\[71\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5788 a_12039_17687# a_12323_17673# a_12258_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5789 tdc0.w_dly_sig_n\[30\] tdc0.w_dly_sig_n\[28\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5790 tdc0.w_dly_sig\[97\] tdc0.w_dly_sig\[95\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5792 VPWR tdc0.w_dly_sig_n\[60\] tdc0.w_dly_sig\[61\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5793 a_17130_14709# a_16930_15009# a_17279_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5794 VPWR a_9650_1791# a_9577_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5795 VPWR clknet_4_8_0_clk a_13459_1141# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5796 a_3329_12335# tdc0.o_result\[74\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5797 VPWR a_6619_17973# a_6626_18273# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5798 VPWR a_6779_6575# a_6947_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5799 a_14373_8867# _014_ a_14277_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X5800 VGND a_4095_8725# a_4053_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5801 a_6335_17973# a_6619_17973# a_6554_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5803 a_1113_12021# a_947_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5804 a_9006_15935# a_8838_16189# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5805 _082_ a_9135_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5806 tdc0.w_dly_sig\[39\] tdc0.w_dly_sig_n\[38\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5807 VPWR tdc0.w_dly_sig\[89\] tdc0.w_dly_sig\[91\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5808 _005_ a_10759_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5809 a_18187_10901# ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5810 a_14250_14165# a_14082_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5811 VGND tdc0.w_dly_sig\[76\] tdc0.w_dly_sig_n\[76\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5812 VPWR tdc0.w_dly_sig_n\[121\] tdc0.w_dly_sig_n\[123\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5813 VGND net1 tdc0.w_dly_sig_n\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5814 tdc0.w_dly_sig_n\[37\] tdc0.w_dly_sig_n\[35\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5815 a_7626_5461# a_7458_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5816 tdc0.w_dly_sig\[63\] tdc0.w_dly_sig\[61\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5817 a_7089_4777# a_6099_4405# a_6963_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5818 a_9411_12809# _013_ a_9493_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5819 tdc0.w_dly_sig_n\[49\] tdc0.w_dly_sig_n\[47\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5820 a_11517_10633# _040_ a_11435_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X5821 a_4387_15279# a_3689_15285# a_4130_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5822 tdc0.o_result\[86\] a_6119_4123# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5823 VGND tdc0.w_dly_sig\[95\] tdc0.w_dly_sig_n\[95\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5824 net1 a_18187_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5825 VGND tdc0.w_dly_sig\[128\] tdc0.w_dly_sig_n\[128\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5827 VPWR clknet_4_6_0_clk a_5363_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5828 VGND tdc0.w_dly_sig_n\[86\] tdc0.w_dly_sig_n\[88\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5829 a_3670_8725# a_3502_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5830 tdc0.w_dly_sig_n\[31\] tdc0.w_dly_sig\[31\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5831 VPWR clknet_4_0_0_clk a_5179_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5832 a_7457_15823# a_6467_15823# a_7331_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5833 a_5951_4221# a_5253_3855# a_5694_3967# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5834 a_14917_17455# tdc0.w_dly_sig\[25\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5835 tdc0.w_dly_sig\[28\] tdc0.w_dly_sig_n\[27\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5836 a_1846_6575# a_1407_6581# a_1761_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5837 VGND _020_ a_13908_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5838 tdc0.w_dly_sig\[95\] tdc0.w_dly_sig\[93\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5839 a_14591_14191# a_13809_14197# a_14507_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5840 VPWR a_7699_4221# a_7867_4123# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5841 tdc0.w_dly_sig_n\[96\] tdc0.w_dly_sig_n\[94\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5842 VPWR a_7263_17673# a_7270_17577# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5843 VGND tdc0.w_dly_sig_n\[100\] tdc0.w_dly_sig\[101\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5844 _075_ a_11251_8457# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5845 a_7366_1135# a_7093_1141# a_7281_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5846 a_15128_17833# a_14729_17461# a_15002_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5847 VGND tdc0.w_dly_sig\[37\] tdc0.w_dly_sig\[39\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5849 tdc0.w_dly_sig_n\[25\] tdc0.w_dly_sig\[25\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5850 a_16166_12335# _071_ a_16332_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5851 VGND a_4463_1109# a_4421_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5852 VPWR a_7775_9813# a_7691_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5853 a_14917_4399# tdc0.w_dly_sig\[108\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5854 VPWR a_13606_3285# a_13533_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5855 VGND tdc0.w_dly_sig\[39\] tdc0.w_dly_sig_n\[39\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5856 VPWR tdc0.o_result\[3\] a_16248_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X5857 tdc0.w_dly_sig_n\[3\] tdc0.w_dly_sig_n\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5858 tdc0.w_dly_sig\[91\] tdc0.w_dly_sig\[89\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5859 VPWR a_9650_7637# _025_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5860 a_5621_15101# a_5087_14735# a_5526_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5861 a_2014_6549# a_1846_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5862 VGND _010_ a_6169_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X5863 a_11456_10927# _041_ a_11290_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5864 tdc0.w_dly_sig_n\[102\] tdc0.w_dly_sig_n\[100\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5865 a_15906_10495# a_15738_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5866 a_5802_2045# a_5529_1679# a_5717_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5867 tdc0.w_dly_sig_n\[59\] tdc0.w_dly_sig\[59\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5868 VGND tdc0.w_dly_sig_n\[104\] tdc0.w_dly_sig_n\[106\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5869 VGND a_7442_6143# a_7400_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5870 a_11333_8457# tdc0.o_result\[73\] a_11251_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5871 VGND tdc0.w_dly_sig\[15\] a_11957_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5872 a_3670_8725# a_3502_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5873 a_12345_4399# _015_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X5874 VPWR clknet_4_2_0_clk a_6927_1141# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5875 a_1987_11837# a_1205_11471# a_1903_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5876 a_5694_14847# a_5526_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5877 tdc0.w_dly_sig_n\[19\] tdc0.w_dly_sig_n\[17\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5878 a_8753_1135# tdc0.w_dly_sig\[94\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5879 a_14519_9447# a_14615_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5880 a_6863_6575# a_6081_6581# a_6779_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5881 VGND a_4739_5211# a_4697_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5882 a_13541_8751# tdc0.o_result\[20\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5884 a_17060_1513# a_16661_1141# a_16934_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5885 VPWR _022_ a_2593_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5886 VGND a_4295_10927# a_4463_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5888 tdc0.w_dly_sig_n\[23\] tdc0.w_dly_sig\[23\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5889 VGND a_11122_7637# _029_ VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X5890 VGND tdc0.w_dly_sig\[53\] tdc0.w_dly_sig_n\[53\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5891 VPWR tdc0.w_dly_sig\[109\] a_8921_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5892 _041_ a_11435_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X5893 VPWR a_14066_1109# a_13993_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5894 tdc0.o_result\[75\] a_2071_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5895 VPWR a_3790_7119# clknet_4_1_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5896 VPWR tdc0.w_dly_sig_n\[62\] tdc0.w_dly_sig_n\[64\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5898 tdc0.w_dly_sig\[101\] tdc0.w_dly_sig\[99\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5900 a_2585_17461# a_2419_17461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5902 a_7185_7669# a_7019_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5903 a_16967_7119# a_16831_7093# a_16547_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5904 VPWR a_3348_13077# clknet_4_5_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5905 VGND tdc0.w_dly_sig\[52\] tdc0.w_dly_sig\[54\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5906 VPWR a_11403_13321# a_11410_13225# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5907 a_17774_16644# a_17567_16585# a_17950_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5908 a_8819_7637# _023_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X5909 a_9006_1109# a_8838_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5910 a_1903_9661# a_1205_9295# a_1646_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5911 a_14002_10116# a_13802_9961# a_14151_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5912 VPWR a_11058_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5913 a_17843_14409# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5914 tdc0.w_dly_sig_n\[93\] tdc0.w_dly_sig_n\[91\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5915 a_8367_4617# clknet_4_2_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5916 VPWR tdc0.w_dly_sig_n\[22\] tdc0.w_dly_sig_n\[24\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5917 tdc0.w_dly_sig_n\[69\] tdc0.w_dly_sig\[69\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5918 tdc0.w_dly_sig_n\[47\] tdc0.w_dly_sig_n\[45\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5919 tdc0.w_dly_sig\[8\] tdc0.w_dly_sig_n\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5920 tdc0.w_dly_sig_n\[2\] tdc0.w_dly_sig\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5922 a_7001_3855# a_6835_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5923 a_16661_1141# a_16495_1141# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5925 VPWR clknet_4_5_0_clk a_4167_17461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5926 VPWR tdc0.w_dly_sig\[16\] tdc0.w_dly_sig\[18\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5927 VPWR tdc0.w_dly_sig\[57\] tdc0.w_dly_sig\[59\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5928 a_11159_4943# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.21 ps=1.42 w=1 l=0.15
X5929 a_1995_13103# a_1131_13109# a_1738_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5930 VGND tdc0.w_dly_sig\[104\] tdc0.w_dly_sig\[106\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5931 a_1938_10927# a_1499_10933# a_1853_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5932 tdc0.w_dly_sig_n\[35\] tdc0.w_dly_sig\[35\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5934 VGND tdc0.w_dly_sig_n\[44\] tdc0.w_dly_sig_n\[46\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5935 a_1972_6953# a_1573_6581# a_1846_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5936 a_13533_3311# a_12999_3317# a_13438_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5937 a_14002_10116# a_13795_10057# a_14178_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5938 _078_ a_9319_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5939 VGND tdc0.w_dly_sig\[105\] tdc0.w_dly_sig\[107\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5940 VGND tdc0.w_dly_sig\[111\] tdc0.w_dly_sig\[113\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5941 a_7373_5487# tdc0.w_dly_sig\[35\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5942 a_1665_13103# a_1131_13109# a_1570_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5943 VPWR net4 a_10446_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5944 VPWR a_5694_14847# a_5621_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5945 a_9650_9407# a_9482_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5946 VPWR _096_ a_16600_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X5947 a_8565_1141# a_8399_1141# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5948 a_17157_10749# a_16819_10535# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5949 a_2750_14165# a_2582_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5950 a_13997_6575# tdc0.w_dly_sig\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5951 VPWR a_7442_3967# a_7369_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5953 a_16013_14735# a_15023_14735# a_15887_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5954 a_13695_3829# a_13986_4129# a_13937_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5955 tdc0.o_result\[104\] a_16331_1947# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5956 VPWR tdc0.w_dly_sig\[83\] tdc0.w_dly_sig_n\[83\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5957 VGND a_17038_7093# a_16967_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X5958 tdc0.o_result\[69\] a_4739_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5959 a_2582_14191# a_2309_14197# a_2497_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5960 a_9723_18365# a_8859_17999# a_9466_18111# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5961 VPWR tdc0.w_dly_sig_n\[2\] tdc0.w_dly_sig_n\[4\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5962 tdc0.w_dly_sig_n\[42\] tdc0.w_dly_sig_n\[40\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5963 VPWR tdc0.w_dly_sig_n\[82\] tdc0.w_dly_sig\[83\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5964 VGND tdc0.w_dly_sig_n\[75\] tdc0.w_dly_sig_n\[77\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5965 VGND tdc0.w_dly_sig_n\[118\] tdc0.w_dly_sig_n\[120\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5966 VGND net3 a_11938_8253# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5967 tdc0.w_dly_sig_n\[122\] tdc0.w_dly_sig\[122\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5968 VGND tdc0.w_dly_sig_n\[23\] tdc0.w_dly_sig\[24\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5969 VGND a_4279_10651# a_4237_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5970 a_8102_10927# a_7663_10933# a_8017_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5971 VPWR tdc0.w_dly_sig_n\[0\] tdc0.w_dly_sig\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5972 a_9393_18365# a_8859_17999# a_9298_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5973 a_14250_6549# a_14082_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5974 a_5989_12021# a_5823_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5975 tdc0.w_dly_sig_n\[57\] tdc0.w_dly_sig_n\[55\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5976 a_12200_9545# _005_ a_12284_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5977 a_15657_6281# _065_ a_15575_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X5978 VPWR tdc0.w_dly_sig\[62\] tdc0.w_dly_sig_n\[62\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5979 VGND net8 a_11146_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X5981 VPWR a_2271_6575# a_2439_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5982 VGND a_6119_15003# a_6077_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5983 a_9466_18111# a_9298_18365# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5984 VGND clknet_4_4_0_clk a_1223_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5985 VGND a_3451_17429# a_3409_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5986 a_9206_4221# a_8767_3855# a_9121_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5987 tdc0.w_dly_sig_n\[13\] tdc0.w_dly_sig\[13\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5988 VPWR _007_ a_10229_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5989 VGND tdc0.w_dly_sig_n\[122\] tdc0.w_dly_sig\[123\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5990 VGND a_2750_14165# a_2708_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5991 VPWR a_11403_12233# a_11410_12137# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5992 a_10598_14709# a_10398_15009# a_10747_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5993 tdc0.o_result\[80\] a_2991_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5994 tdc0.o_result\[109\] a_9799_4123# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5995 VGND tdc0.w_dly_sig_n\[54\] tdc0.w_dly_sig_n\[56\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5996 a_9761_7119# _000_ a_9661_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X5998 tdc0.w_dly_sig_n\[38\] tdc0.w_dly_sig\[38\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5999 a_2823_3311# a_1959_3317# a_2566_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6000 a_11619_8867# _073_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6001 a_15669_5807# _015_ a_15235_5719# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6002 a_16831_7093# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6003 VPWR tdc0.w_dly_sig\[56\] tdc0.w_dly_sig_n\[56\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6004 a_7001_3855# a_6835_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6005 a_10239_12015# _026_ a_10321_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6006 VPWR a_1738_13077# a_1665_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6007 tdc0.w_dly_sig_n\[35\] tdc0.w_dly_sig_n\[33\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6008 a_6821_15823# tdc0.w_dly_sig\[42\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6009 a_10423_5193# _020_ a_10505_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6011 a_1301_12015# tdc0.w_dly_sig\[75\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6012 a_17443_1135# a_16661_1141# a_17359_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6013 a_13809_6581# a_13643_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6014 a_10226_6575# _003_ a_10029_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6015 VGND tdc0.o_result\[4\] a_14786_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6016 a_6756_11305# a_6357_10933# a_6630_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6017 tdc0.w_dly_sig_n\[65\] tdc0.w_dly_sig_n\[63\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6018 a_17335_10383# a_17206_10657# a_16915_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6019 VGND a_2623_17179# a_2581_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6020 VPWR a_5291_13077# a_5207_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6021 VGND tdc0.o_result\[7\] a_11892_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X6022 VPWR tdc0.w_dly_sig\[41\] tdc0.w_dly_sig_n\[41\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6023 VPWR a_12548_4917# clknet_4_8_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6025 a_3927_8751# a_3063_8757# a_3670_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6026 VPWR a_7534_1109# a_7461_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6027 VGND a_15595_17429# a_15553_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6029 tdc0.o_result\[36\] a_6671_13915# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6030 a_6979_17687# a_7263_17673# a_7198_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6031 a_2539_8751# a_1757_8757# a_2455_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6032 VPWR tdc0.w_dly_sig\[10\] a_11957_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6033 tdc0.w_dly_sig_n\[36\] tdc0.w_dly_sig\[36\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6034 VGND tdc0.w_dly_sig\[80\] tdc0.w_dly_sig\[82\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6035 VPWR a_7258_9407# a_7185_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6036 a_18187_10901# ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6037 tdc0.w_dly_sig_n\[28\] tdc0.w_dly_sig\[28\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6038 a_18121_17833# a_17567_17673# a_17774_17732# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6039 VPWR a_13605_4917# _074_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6040 a_10046_4676# a_9846_4521# a_10195_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6041 a_18326_7940# a_18119_7881# a_18502_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6042 a_7350_9813# a_7182_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6043 a_8746_17455# a_8473_17461# a_8661_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6044 tdc0.o_result\[86\] a_6119_4123# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6045 a_10107_14709# a_10391_14709# a_10326_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6047 tdc0.w_dly_sig_n\[22\] tdc0.w_dly_sig\[22\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6048 VPWR a_5970_1791# a_5897_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6049 a_16117_8457# tdc0.o_result\[27\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6050 tdc0.w_dly_sig_n\[1\] tdc0.w_dly_sig\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6051 tdc0.w_dly_sig\[44\] tdc0.w_dly_sig\[42\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6052 VPWR tdc0.w_dly_sig_n\[117\] tdc0.w_dly_sig\[118\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6053 a_9389_9071# tdc0.o_result\[33\] a_9043_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6054 a_14715_15797# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6055 VPWR a_9466_18111# a_9393_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6056 a_6645_10633# _099_ a_6549_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6057 tdc0.w_dly_sig_n\[86\] tdc0.w_dly_sig\[86\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6058 a_9834_3285# a_9666_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6059 uo_out[7] a_11504_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6060 tdc0.w_dly_sig_n\[101\] tdc0.w_dly_sig\[101\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6061 VGND tdc0.w_dly_sig\[111\] tdc0.w_dly_sig_n\[111\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6062 a_9209_1679# a_9043_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6063 a_12518_7119# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X6064 a_13358_11204# a_13158_11049# a_13507_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6065 tdc0.w_dly_sig_n\[55\] tdc0.w_dly_sig_n\[53\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6067 a_7883_5487# a_7019_5493# a_7626_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6068 VGND _019_ a_9205_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6069 a_7189_6031# tdc0.w_dly_sig\[33\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6070 VPWR tdc0.w_dly_sig\[37\] tdc0.w_dly_sig_n\[37\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6071 a_5115_6575# a_4333_6581# a_5031_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6072 a_4054_3311# a_3615_3317# a_3969_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6073 a_13997_14191# tdc0.w_dly_sig\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6074 a_13813_1135# tdc0.w_dly_sig\[100\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6075 tdc0.w_dly_sig_n\[121\] tdc0.w_dly_sig\[121\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6076 VPWR tdc0.w_dly_sig_n\[31\] tdc0.w_dly_sig_n\[33\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6077 VPWR tdc0.w_dly_sig_n\[111\] tdc0.w_dly_sig\[112\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6078 VPWR tdc0.w_dly_sig_n\[87\] tdc0.w_dly_sig\[88\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6079 VGND a_18326_7940# a_18255_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6080 VGND tdc0.w_dly_sig_n\[106\] tdc0.w_dly_sig_n\[108\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6081 _023_ _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6082 VPWR tdc0.w_dly_sig\[14\] tdc0.w_dly_sig\[16\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6083 a_18163_3689# a_18027_3529# a_17743_3543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6084 a_9332_3855# a_8933_3855# a_9206_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6085 tdc0.w_dly_sig_n\[78\] tdc0.w_dly_sig\[78\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6086 a_2673_1513# a_1683_1141# a_2547_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6087 tdc0.o_result\[104\] a_16331_1947# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6088 VPWR tdc0.w_dly_sig_n\[62\] tdc0.w_dly_sig\[63\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6089 VGND clknet_4_6_0_clk a_5363_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6090 VGND a_2531_10901# a_2489_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6091 VPWR a_17647_12247# tdc0.o_result\[120\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6092 VGND tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6093 a_18121_2767# a_17567_2741# a_17774_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6094 a_8399_12809# _013_ a_8481_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6095 tdc0.w_dly_sig_n\[12\] tdc0.w_dly_sig\[12\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6097 VGND tdc0.w_dly_sig_n\[125\] tdc0.w_dly_sig\[126\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6098 VGND tdc0.w_dly_sig_n\[74\] tdc0.w_dly_sig_n\[76\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6099 VPWR a_11504_11445# uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6100 tdc0.w_dly_sig_n\[74\] tdc0.w_dly_sig\[74\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6101 a_10046_4676# a_9839_4617# a_10222_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6102 VGND clknet_4_3_0_clk a_6835_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6103 VGND a_7039_8475# a_6997_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6104 a_8746_17455# a_8307_17461# a_8661_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6105 VGND net28 a_12893_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6107 a_14944_12809# _091_ a_14676_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6108 VPWR tdc0.w_dly_sig_n\[120\] tdc0.w_dly_sig\[121\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6109 VPWR tdc0.w_dly_sig\[100\] tdc0.w_dly_sig\[102\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6110 a_9650_1791# a_9482_2045# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6112 VGND tdc0.w_dly_sig\[54\] tdc0.w_dly_sig\[56\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6113 tdc0.w_dly_sig\[27\] tdc0.w_dly_sig\[25\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6114 VGND a_5970_12671# a_5928_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6115 a_10107_14709# a_10398_15009# a_10349_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6116 a_7461_1135# a_6927_1141# a_7366_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6118 a_11058_9839# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6119 VPWR tdc0.o_result\[97\] a_12345_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X6120 a_12058_4221# a_11619_3855# a_11973_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6123 VPWR a_15595_15253# a_15511_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6124 a_5441_14735# tdc0.w_dly_sig\[39\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6125 VPWR _009_ a_13541_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6127 VPWR a_15235_5719# _085_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X6128 a_7185_9661# a_6651_9295# a_7090_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6129 tdc0.w_dly_sig_n\[44\] tdc0.w_dly_sig\[44\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6130 tdc0.w_dly_sig_n\[0\] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6131 VGND clknet_4_0_0_clk a_1959_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6132 VGND a_17314_12559# clknet_4_14_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6133 VPWR tdc0.w_dly_sig\[55\] tdc0.w_dly_sig\[57\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6134 a_18502_7663# a_18255_8041# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6135 VPWR a_12771_11159# tdc0.o_result\[5\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6136 a_14707_13335# a_14998_13225# a_14949_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6137 VPWR a_4111_18365# a_4279_18267# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6138 a_2271_6575# a_1407_6581# a_2014_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6139 tdc0.o_result\[37\] a_9431_16091# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6140 uo_out[2] a_14676_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6142 VPWR tdc0.w_dly_sig_n\[58\] tdc0.w_dly_sig\[59\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6143 tdc0.w_dly_sig\[40\] tdc0.w_dly_sig\[38\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6144 VGND a_4111_10749# a_4279_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6145 VPWR tdc0.w_dly_sig_n\[79\] tdc0.w_dly_sig\[80\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6146 VGND tdc0.w_dly_sig\[87\] tdc0.w_dly_sig\[89\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6147 a_6449_6575# a_5915_6581# a_6354_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6148 a_8399_6575# _028_ a_8481_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6149 a_8013_12021# a_7847_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6150 tdc0.w_dly_sig\[34\] tdc0.w_dly_sig_n\[33\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6151 VPWR tdc0.w_dly_sig\[102\] tdc0.w_dly_sig_n\[102\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6152 VPWR tdc0.w_dly_sig\[101\] tdc0.w_dly_sig\[103\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6153 a_10393_4777# a_9839_4617# a_10046_4676# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6154 a_9595_11721# _013_ a_9677_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6155 tdc0.w_dly_sig_n\[79\] tdc0.w_dly_sig_n\[77\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6156 VGND a_16155_14423# _089_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6157 VPWR a_7055_10927# a_7223_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6158 a_17865_8457# _025_ a_17719_8359# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X6159 VGND clknet_4_7_0_clk a_8399_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6160 VGND a_9485_7485# _028_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0991 ps=0.955 w=0.65 l=0.15
X6161 VGND a_17187_16599# tdc0.o_result\[125\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6162 VGND tdc0.w_dly_sig\[121\] tdc0.w_dly_sig\[123\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6163 tdc0.w_dly_sig_n\[54\] tdc0.w_dly_sig_n\[52\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6164 tdc0.w_dly_sig_n\[24\] tdc0.w_dly_sig\[24\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6165 a_7733_3689# a_6743_3317# a_7607_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6167 VPWR clknet_4_13_0_clk a_13643_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6168 VPWR clknet_4_1_0_clk a_4167_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6169 VPWR tdc0.w_dly_sig_n\[67\] tdc0.w_dly_sig_n\[69\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6170 tdc0.w_dly_sig\[32\] tdc0.w_dly_sig\[30\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6171 a_15235_5719# tdc0.o_result\[98\] a_15381_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6172 VGND net1 tdc0.w_dly_sig_n\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6173 a_6549_7369# tdc0.o_result\[64\] a_6467_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6174 a_4330_2045# a_3891_1679# a_4245_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6175 tdc0.w_dly_sig_n\[74\] tdc0.w_dly_sig_n\[72\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6176 a_12323_17673# clknet_4_13_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6177 a_11023_12247# a_11119_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6178 VPWR a_14507_14191# a_14675_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6179 VGND _092_ a_16127_7779# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6180 VGND _012_ a_10585_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6181 VPWR a_15106_9269# a_15035_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6182 a_14460_4943# tdc0.o_result\[100\] a_14157_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X6183 VGND clknet_0_clk a_7856_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X6184 a_9209_9295# a_9043_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6185 a_13879_17973# a_14163_17973# a_14098_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6186 a_4180_3689# a_3781_3317# a_4054_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6187 a_9907_9661# a_9043_9295# a_9650_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6188 VGND a_11058_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6189 VGND _010_ a_6813_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6190 VGND clknet_0_clk a_16762_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6191 tdc0.w_dly_sig_n\[59\] tdc0.w_dly_sig_n\[57\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6192 VGND a_11058_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X6194 VGND clknet_0_clk a_12548_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X6195 a_13091_7779# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X6196 a_16858_14735# a_16543_14887# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6197 a_16155_17687# tdc0.o_result\[126\] a_16301_17775# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X6198 VGND _012_ a_14081_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6199 a_10222_4399# a_9975_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6200 a_5897_12925# a_5363_12559# a_5802_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6201 VGND a_9374_3967# a_9332_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6202 VGND a_6550_13103# clknet_4_6_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6203 a_13937_15101# a_13599_14887# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6204 VPWR a_12134_6549# _010_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6205 a_8270_10901# a_8102_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6206 a_16451_7271# a_16547_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6207 a_9401_12015# tdc0.o_result\[57\] a_9319_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6208 VPWR net1 tdc0.w_dly_sig_n\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6209 VGND a_7775_9813# a_7733_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6210 VGND a_9282_13077# a_9240_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6211 tdc0.w_dly_sig\[80\] tdc0.w_dly_sig_n\[79\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6212 tdc0.o_result\[30\] a_10075_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6213 tdc0.w_dly_sig_n\[123\] tdc0.w_dly_sig_n\[121\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6214 VGND tdc0.w_dly_sig\[122\] tdc0.w_dly_sig\[124\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6215 VGND tdc0.w_dly_sig_n\[126\] tdc0.w_dly_sig_n\[128\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6216 a_4019_5487# a_3321_5493# a_3762_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6217 VPWR tdc0.w_dly_sig_n\[118\] tdc0.w_dly_sig\[119\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6218 a_8399_11721# _013_ a_8481_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6219 a_11957_14569# a_11410_14313# a_11610_14468# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6220 VPWR tdc0.w_dly_sig\[16\] tdc0.w_dly_sig_n\[16\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6221 _013_ a_11159_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.327 ps=1.65 w=1 l=0.15
X6222 VPWR a_3698_12559# clknet_4_4_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6223 VPWR a_2991_3285# a_2907_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6224 VGND a_8367_4617# a_8374_4521# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6225 VGND tdc0.w_dly_sig_n\[117\] tdc0.w_dly_sig_n\[119\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6226 a_18226_14191# a_17979_14569# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6227 a_18199_14557# a_17979_14569# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6228 VGND tdc0.w_dly_sig\[76\] tdc0.w_dly_sig\[78\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6229 a_9539_13103# a_8841_13109# a_9282_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6230 a_3781_3317# a_3615_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6231 a_7055_10927# a_6191_10933# a_6798_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6232 VGND tdc0.w_dly_sig_n\[115\] tdc0.w_dly_sig_n\[117\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6233 a_12184_3855# a_11785_3855# a_12058_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6234 a_3785_1135# tdc0.w_dly_sig\[85\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6235 a_14922_15797# a_14715_15797# a_15098_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6236 VGND tdc0.w_dly_sig_n\[77\] tdc0.w_dly_sig\[78\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6238 a_9114_13103# a_8675_13109# a_9029_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6239 a_2593_10633# tdc0.o_result\[51\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6240 VGND a_14388_13621# clknet_4_13_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6241 tdc0.o_result\[99\] a_14491_1109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6242 VPWR a_11610_14468# a_11539_14569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6243 VPWR a_14664_6005# clknet_4_9_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6244 tdc0.w_dly_sig_n\[101\] tdc0.w_dly_sig_n\[99\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6245 _003_ a_14287_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X6246 VGND tdc0.w_dly_sig_n\[93\] tdc0.w_dly_sig\[94\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6247 VGND a_14664_6005# clknet_4_9_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6248 VGND a_2547_3133# a_2715_3035# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6249 VGND tdc0.w_dly_sig_n\[19\] tdc0.w_dly_sig_n\[21\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6250 _016_ _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6251 tdc0.w_dly_sig\[120\] tdc0.w_dly_sig\[118\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6253 VGND clknet_4_14_0_clk a_15299_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6254 tdc0.w_dly_sig\[18\] tdc0.w_dly_sig\[16\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6255 a_16589_6031# _020_ a_16155_6183# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6256 tdc0.w_dly_sig\[117\] tdc0.w_dly_sig_n\[116\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6257 a_14507_14191# a_13643_14197# a_14250_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6259 VPWR tdc0.w_dly_sig\[58\] tdc0.w_dly_sig_n\[58\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6260 VGND a_13863_3311# a_14031_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6261 a_13879_17973# a_14170_18273# a_14121_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6262 tdc0.w_dly_sig_n\[65\] tdc0.w_dly_sig\[65\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6264 VPWR a_4739_5211# a_4655_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6265 _092_ a_8399_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X6266 _073_ a_10975_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X6267 VPWR net3 a_11938_8253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X6268 a_15646_18365# a_15207_17999# a_15561_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6269 a_4038_1109# a_3870_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6270 tdc0.w_dly_sig\[39\] tdc0.w_dly_sig\[37\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6271 tdc0.o_result\[109\] a_9799_4123# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6272 VPWR _000_ a_10147_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6273 VPWR a_8730_16341# a_8657_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6274 VPWR tdc0.w_dly_sig_n\[107\] tdc0.w_dly_sig_n\[109\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6275 VPWR a_17199_10357# a_17206_10657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6276 a_14177_14191# a_13643_14197# a_14082_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6277 tdc0.w_dly_sig_n\[124\] tdc0.w_dly_sig_n\[122\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6278 a_1853_10927# tdc0.w_dly_sig\[52\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6279 tdc0.o_result\[64\] a_6027_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6281 a_13990_8573# a_13717_8207# a_13905_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6282 tdc0.w_dly_sig_n\[39\] tdc0.w_dly_sig_n\[37\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6283 a_11290_11247# _041_ a_11456_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6284 tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6285 a_4456_1679# a_4057_1679# a_4330_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6286 VPWR a_17406_4917# a_17335_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6287 VGND tdc0.w_dly_sig\[119\] tdc0.w_dly_sig\[121\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6288 a_7653_17161# tdc0.o_result\[40\] a_7571_17161# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6289 a_5526_4221# a_5087_3855# a_5441_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6290 VPWR tdc0.w_dly_sig\[70\] tdc0.w_dly_sig_n\[70\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6291 a_6446_8573# a_6173_8207# a_6361_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6292 a_6099_16367# _029_ a_6181_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6293 VGND tdc0.w_dly_sig_n\[14\] tdc0.w_dly_sig_n\[16\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6294 tdc0.w_dly_sig\[81\] tdc0.w_dly_sig_n\[80\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6295 tdc0.w_dly_sig\[87\] tdc0.w_dly_sig\[85\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6296 a_17125_1679# tdc0.w_dly_sig\[104\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6297 tdc0.w_dly_sig\[25\] tdc0.w_dly_sig_n\[24\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6298 VGND net10 a_9665_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6299 VPWR a_16727_18151# tdc0.o_result\[126\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6300 VGND a_11518_2741# a_11447_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6301 tdc0.w_dly_sig_n\[53\] tdc0.w_dly_sig\[53\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6302 VPWR tdc0.w_dly_sig\[34\] tdc0.w_dly_sig\[36\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6303 VPWR a_18142_6852# a_18071_6953# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6304 tdc0.w_dly_sig_n\[75\] tdc0.w_dly_sig_n\[73\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6305 a_13415_10071# a_13511_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6306 a_16831_7093# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6308 tdc0.w_dly_sig\[84\] tdc0.w_dly_sig_n\[83\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6309 VGND tdc0.w_dly_sig\[109\] tdc0.w_dly_sig_n\[109\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6310 VGND tdc0.w_dly_sig_n\[23\] tdc0.w_dly_sig_n\[25\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6311 VPWR a_4555_15253# a_4471_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6312 a_3597_1141# a_3431_1141# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6313 a_12165_10633# _044_ a_12069_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6314 a_18050_14468# a_17843_14409# a_18226_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6315 _014_ a_13735_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6316 VGND a_16819_10535# tdc0.o_result\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6317 VPWR a_17843_14409# a_17850_14313# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6318 a_9411_2223# _028_ a_9493_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6319 VPWR tdc0.w_dly_sig_n\[71\] tdc0.w_dly_sig\[72\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6320 VPWR tdc0.w_dly_sig\[20\] tdc0.w_dly_sig_n\[20\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6321 VGND tdc0.w_dly_sig\[128\] a_18121_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6322 tdc0.w_dly_sig_n\[109\] tdc0.w_dly_sig_n\[107\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6323 tdc0.w_dly_sig\[35\] tdc0.w_dly_sig_n\[34\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6324 tdc0.w_dly_sig_n\[52\] tdc0.w_dly_sig_n\[50\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6325 a_7987_4631# a_8083_4631# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6326 VGND a_4774_6549# a_4732_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6327 a_13783_18151# a_13879_17973# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6328 VGND a_12226_3967# a_12184_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6329 a_14250_6549# a_14082_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6330 VGND clknet_4_5_0_clk a_3523_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6331 VPWR a_4176_6005# clknet_4_0_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6332 VPWR a_14370_17973# a_14299_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6333 tdc0.w_dly_sig_n\[82\] tdc0.w_dly_sig_n\[80\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6334 a_6629_13647# a_5639_13647# a_6503_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6335 tdc0.w_dly_sig\[87\] tdc0.w_dly_sig_n\[86\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6336 a_1696_13481# a_1297_13109# a_1570_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6337 a_18673_8041# a_18126_7785# a_18326_7940# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6338 a_9623_13103# a_8841_13109# a_9539_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6339 tdc0.w_dly_sig_n\[46\] tdc0.w_dly_sig_n\[44\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6340 VPWR clknet_4_0_0_clk a_3891_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6341 VPWR a_15807_12711# tdc0.o_result\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6342 a_12679_17821# a_12459_17833# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6343 clknet_4_1_0_clk a_3790_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6344 VPWR a_14415_8573# a_14583_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6345 VGND net7 a_5433_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6346 a_7093_1141# a_6927_1141# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6347 VGND tdc0.w_dly_sig\[20\] tdc0.w_dly_sig\[22\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6348 VPWR a_17314_12559# clknet_4_14_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6349 tdc0.w_dly_sig\[110\] tdc0.w_dly_sig\[108\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6350 a_1478_9661# a_1039_9295# a_1393_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6351 a_9209_1679# a_9043_1679# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6352 a_17703_17833# a_17567_17673# a_17283_17687# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6353 VGND tdc0.w_dly_sig\[97\] tdc0.w_dly_sig_n\[97\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6354 a_5529_1679# a_5363_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6355 VPWR a_11058_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6356 tdc0.w_dly_sig\[31\] tdc0.w_dly_sig\[29\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6357 VPWR a_6871_8573# a_7039_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6358 a_15327_13799# tdc0.o_result\[12\] a_15473_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X6359 VPWR tdc0.w_dly_sig_n\[84\] tdc0.w_dly_sig\[85\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6360 a_17923_16733# a_17703_16745# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6362 tdc0.w_dly_sig_n\[86\] tdc0.w_dly_sig_n\[84\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6364 VGND clknet_4_7_0_clk a_8859_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6366 VGND a_4498_1791# a_4456_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6367 VPWR a_9263_1135# a_9431_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6368 a_9263_1135# a_8565_1141# a_9006_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6369 tdc0.w_dly_sig\[12\] tdc0.w_dly_sig\[10\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6370 a_9807_17687# tdc0.o_result\[21\] a_9953_17775# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X6371 a_5652_3855# a_5253_3855# a_5526_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6372 tdc0.o_result\[95\] a_10075_1947# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6374 VPWR tdc0.w_dly_sig\[69\] tdc0.w_dly_sig\[71\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6375 a_18326_7940# a_18126_7785# a_18475_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6376 VPWR tdc0.w_dly_sig\[124\] tdc0.w_dly_sig\[126\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6377 VGND a_7286_7119# clknet_4_3_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X6378 tdc0.w_dly_sig\[30\] tdc0.w_dly_sig_n\[29\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6379 VGND tdc0.w_dly_sig\[93\] tdc0.w_dly_sig\[95\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6380 VPWR tdc0.w_dly_sig\[66\] tdc0.w_dly_sig\[68\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6381 tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6382 tdc0.w_dly_sig_n\[111\] tdc0.w_dly_sig_n\[109\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6383 tdc0.w_dly_sig_n\[26\] tdc0.w_dly_sig\[26\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6384 tdc0.w_dly_sig_n\[83\] tdc0.w_dly_sig_n\[81\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6386 a_10393_4777# a_9846_4521# a_10046_4676# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6387 VPWR net2 a_13919_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X6388 a_12284_9545# _081_ a_12118_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6389 a_6817_9295# a_6651_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6390 tdc0.w_dly_sig_n\[106\] tdc0.w_dly_sig_n\[104\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6391 VGND tdc0.w_dly_sig\[9\] tdc0.w_dly_sig\[11\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6392 VPWR _007_ a_8481_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6393 VGND a_13979_14709# a_13986_15009# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6394 VPWR net9 a_11057_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6396 VGND _010_ a_4881_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6397 VGND a_2455_8751# a_2623_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6398 clknet_4_6_0_clk a_6550_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6399 a_14834_9295# a_14519_9447# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6400 a_4774_6549# a_4606_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6401 VGND clknet_4_2_0_clk a_9227_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6402 VGND a_4571_5309# a_4739_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6403 a_5652_14735# a_5253_14735# a_5526_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6404 tdc0.w_dly_sig\[60\] tdc0.w_dly_sig\[58\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6405 VGND a_7591_2197# a_7549_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6406 _038_ a_9411_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X6407 tdc0.o_result\[46\] a_4279_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6409 _029_ a_11122_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6410 VGND tdc0.w_dly_sig\[32\] tdc0.w_dly_sig\[34\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6411 tdc0.w_dly_sig\[20\] tdc0.w_dly_sig_n\[19\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6412 a_5169_9545# tdc0.o_result\[46\] a_5087_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6413 a_17739_7895# a_17835_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6414 a_8454_11989# a_8286_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6415 a_17187_17687# a_17283_17687# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6416 a_16849_1135# tdc0.w_dly_sig\[102\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6417 a_2037_2767# tdc0.w_dly_sig\[82\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6418 tdc0.w_dly_sig\[85\] tdc0.w_dly_sig_n\[84\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6419 tdc0.w_dly_sig\[89\] tdc0.w_dly_sig_n\[88\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6420 tdc0.w_dly_sig\[102\] tdc0.w_dly_sig_n\[101\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6421 VGND tdc0.w_dly_sig_n\[99\] tdc0.w_dly_sig\[100\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6423 VGND tdc0.w_dly_sig\[49\] tdc0.w_dly_sig\[51\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6424 VGND a_4755_4399# a_4923_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6425 VGND tdc0.w_dly_sig\[126\] tdc0.w_dly_sig\[128\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6426 VPWR tdc0.w_dly_sig_n\[96\] tdc0.w_dly_sig_n\[98\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6427 tdc0.w_dly_sig\[38\] tdc0.w_dly_sig\[36\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6428 VGND a_7791_1135# a_7959_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6429 a_3502_8751# a_3063_8757# a_3417_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6430 a_3965_10927# a_3431_10933# a_3870_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6431 a_9953_17775# net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X6432 VGND tdc0.w_dly_sig\[99\] tdc0.w_dly_sig\[101\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6433 VGND a_14922_15797# a_14851_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6434 VPWR tdc0.w_dly_sig_n\[89\] tdc0.w_dly_sig_n\[91\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6435 a_7263_17673# clknet_4_7_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6436 tdc0.w_dly_sig\[74\] tdc0.w_dly_sig\[72\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6437 a_15002_15279# a_14729_15285# a_14917_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6439 VPWR tdc0.w_dly_sig\[45\] tdc0.w_dly_sig\[47\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6440 a_1604_9295# a_1205_9295# a_1478_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6441 VGND a_8914_17429# a_8872_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6442 VPWR a_14507_6575# a_14675_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6443 VPWR tdc0.w_dly_sig\[66\] tdc0.w_dly_sig_n\[66\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6444 a_14507_6575# a_13809_6581# a_14250_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6445 VGND a_6779_6575# a_6947_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6446 a_8838_1135# a_8565_1141# a_8753_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6447 a_4885_17999# a_4719_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6448 tdc0.w_dly_sig\[107\] tdc0.w_dly_sig\[105\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6449 tdc0.w_dly_sig\[113\] tdc0.w_dly_sig\[111\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6450 VGND a_18119_4617# a_18126_4521# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6451 VPWR tdc0.w_dly_sig\[59\] tdc0.w_dly_sig_n\[59\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6454 VGND a_3698_12559# clknet_4_4_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6455 a_15473_13897# _007_ a_15327_13799# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X6456 a_8753_15823# tdc0.w_dly_sig\[38\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6457 VPWR a_16239_18267# a_16155_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6458 tdc0.o_result\[56\] a_6395_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6459 VGND a_14715_15797# a_14722_16097# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6460 VPWR a_2547_3133# a_2715_3035# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6461 VGND a_5694_3967# a_5652_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6462 VPWR a_6614_8319# a_6541_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6463 VPWR tdc0.w_dly_sig\[21\] a_12877_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6464 VGND _003_ a_10975_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6465 VPWR a_6550_13103# clknet_4_6_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6466 a_18673_8041# a_18119_7881# a_18326_7940# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6467 clknet_4_0_0_clk a_4176_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6468 VPWR net11 a_14829_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6469 a_6311_2045# a_5529_1679# a_6227_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6470 VGND tdc0.w_dly_sig_n\[68\] tdc0.w_dly_sig_n\[70\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6471 VPWR a_4187_5461# a_4103_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6472 a_14195_8867# _011_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6473 tdc0.w_dly_sig_n\[37\] tdc0.w_dly_sig\[37\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6474 tdc0.w_dly_sig_n\[90\] tdc0.w_dly_sig\[90\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6475 a_12318_7637# a_12171_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.331 ps=1.71 w=0.42 l=0.15
X6476 tdc0.w_dly_sig\[16\] tdc0.w_dly_sig\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6478 VPWR tdc0.w_dly_sig_n\[97\] tdc0.w_dly_sig_n\[99\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6479 tdc0.w_dly_sig_n\[28\] tdc0.w_dly_sig_n\[26\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6480 a_12548_4917# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6481 VPWR a_4571_5309# a_4739_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6482 a_1297_13109# a_1131_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6483 tdc0.w_dly_sig_n\[43\] tdc0.w_dly_sig_n\[41\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6484 VPWR clknet_4_0_0_clk a_3615_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6486 VPWR a_13979_14709# a_13986_15009# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6487 VPWR _007_ a_8481_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6488 tdc0.w_dly_sig_n\[103\] tdc0.w_dly_sig_n\[101\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6489 a_3601_17999# tdc0.w_dly_sig\[44\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6490 clknet_0_clk a_11058_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6491 a_10057_10927# tdc0.o_result\[55\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X6492 VPWR tdc0.w_dly_sig_n\[8\] tdc0.w_dly_sig\[9\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6493 VPWR a_11711_591# net5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6494 a_16166_12335# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6495 VPWR clknet_4_9_0_clk a_12999_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6496 VPWR net1 tdc0.w_dly_sig\[2\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6497 _015_ a_12318_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X6498 VGND a_17543_8751# a_17711_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6499 clknet_0_clk a_11058_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6500 tdc0.o_result\[50\] a_2163_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6501 VPWR _002_ a_8543_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0662 ps=0.735 w=0.42 l=0.15
X6502 tdc0.w_dly_sig_n\[66\] tdc0.w_dly_sig\[66\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6503 a_17559_14423# a_17843_14409# a_17778_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6504 tdc0.o_result\[50\] a_2163_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6505 tdc0.w_dly_sig\[121\] tdc0.w_dly_sig_n\[120\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6508 a_4333_17461# a_4167_17461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6509 VPWR tdc0.w_dly_sig_n\[25\] tdc0.w_dly_sig\[26\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6510 a_1945_8751# tdc0.w_dly_sig\[74\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6511 VGND _005_ a_11290_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6513 a_14592_12809# tdc0.o_result\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X6514 VGND clknet_0_clk a_17314_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6515 VPWR tdc0.w_dly_sig_n\[125\] tdc0.w_dly_sig_n\[127\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6516 VPWR tdc0.w_dly_sig\[19\] tdc0.w_dly_sig_n\[19\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6517 VPWR _023_ a_9217_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6518 a_3628_9129# a_3229_8757# a_3502_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6519 a_16332_9839# _101_ a_16600_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6520 VPWR a_12376_8751# uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X6521 VPWR net5 a_11067_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X6522 tdc0.w_dly_sig\[32\] tdc0.w_dly_sig_n\[31\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6523 a_18325_9071# _015_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X6524 VPWR a_6671_13915# a_6587_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6525 tdc0.w_dly_sig\[63\] tdc0.w_dly_sig_n\[62\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6526 _028_ a_9485_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.104 ps=1 w=0.65 l=0.15
X6527 VPWR a_14676_12809# uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6528 VGND a_7055_10927# a_7223_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6529 VGND a_1646_9407# a_1604_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6531 VGND a_13183_6583# _002_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X6532 VPWR tdc0.w_dly_sig\[5\] tdc0.w_dly_sig\[7\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6533 VPWR clknet_4_6_0_clk a_7847_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6534 VPWR _032_ a_9753_11043# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X6535 VGND tdc0.w_dly_sig_n\[119\] tdc0.w_dly_sig_n\[121\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6536 VGND tdc0.w_dly_sig\[40\] tdc0.w_dly_sig\[42\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6537 a_6541_8573# a_6007_8207# a_6446_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6538 tdc0.w_dly_sig\[37\] tdc0.w_dly_sig_n\[36\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6539 uo_out[0] a_16332_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X6540 a_11329_1679# tdc0.w_dly_sig\[98\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6541 a_11333_15279# tdc0.o_result\[41\] a_11251_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6543 a_15738_2045# a_15299_1679# a_15653_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6544 _005_ a_10759_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X6545 VPWR tdc0.w_dly_sig\[65\] tdc0.w_dly_sig_n\[65\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6546 VPWR tdc0.w_dly_sig_n\[7\] tdc0.w_dly_sig\[8\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6547 VGND clknet_4_8_0_clk a_11619_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6548 tdc0.w_dly_sig\[123\] tdc0.w_dly_sig\[121\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6549 a_17739_4631# a_17835_4631# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6550 VGND tdc0.w_dly_sig_n\[9\] tdc0.w_dly_sig\[10\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6551 a_14991_13321# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6552 VGND tdc0.w_dly_sig\[68\] tdc0.w_dly_sig\[70\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6553 tdc0.w_dly_sig\[42\] tdc0.w_dly_sig_n\[41\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6554 VPWR tdc0.w_dly_sig\[100\] tdc0.w_dly_sig_n\[100\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6555 VGND tdc0.w_dly_sig_n\[85\] tdc0.w_dly_sig\[86\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6556 VGND a_11058_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6557 VGND a_1646_11583# a_1604_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6558 a_2079_13103# a_1297_13109# a_1995_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6559 VGND a_12323_17673# a_12330_17577# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6561 tdc0.o_result\[68\] a_6211_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6562 VPWR clknet_4_4_0_clk a_1223_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6563 VGND a_12548_14165# clknet_4_12_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6564 a_15565_7983# _020_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X6565 a_4245_1679# tdc0.w_dly_sig\[86\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6566 a_10401_7369# _002_ a_10595_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6567 VGND a_10046_4676# a_9975_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6568 a_18410_12015# a_18163_12393# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6569 a_4038_1109# a_3870_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
R26 tt_um_hpretl_tt06_tdc_26.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
R27 VPWR tt_um_hpretl_tt06_tdc_27.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6571 a_2290_5055# a_2122_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6572 VPWR a_16332_12015# uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X6573 a_11067_9545# _013_ a_11149_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6574 uo_out[5] a_11456_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X6575 tdc0.w_dly_sig_n\[115\] tdc0.w_dly_sig\[115\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6576 net10 a_13603_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6577 VGND a_17567_16585# a_17574_16489# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6578 VPWR _010_ a_5721_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6579 a_16484_5807# tdc0.o_result\[114\] a_16181_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X6580 VPWR net5 a_11490_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X6581 VPWR tdc0.w_dly_sig_n\[114\] tdc0.w_dly_sig_n\[116\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6583 tdc0.w_dly_sig\[24\] tdc0.w_dly_sig\[22\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6584 a_12237_10633# _043_ a_12165_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6585 a_15373_17999# a_15207_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6586 clknet_4_5_0_clk a_3348_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6587 tdc0.o_result\[119\] a_18171_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6588 VGND a_2255_9813# a_2213_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6589 a_10229_15823# tdc0.o_result\[37\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6590 tdc0.w_dly_sig_n\[110\] tdc0.w_dly_sig\[110\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6591 tdc0.w_dly_sig_n\[128\] tdc0.w_dly_sig_n\[126\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6593 a_7619_17821# a_7399_17833# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6595 VGND tdc0.w_dly_sig\[67\] tdc0.w_dly_sig_n\[67\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6597 VGND a_6798_10901# a_6756_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6598 a_14615_9269# a_14899_9269# a_14834_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6599 a_17243_17999# a_17114_18273# a_16823_17973# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6600 VGND clknet_4_0_0_clk a_3891_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6601 VPWR a_16412_6549# clknet_4_10_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6602 tdc0.w_dly_sig_n\[119\] tdc0.w_dly_sig_n\[117\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6603 VGND a_14388_13621# clknet_4_13_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6604 a_10607_12809# _060_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X6605 VGND tdc0.w_dly_sig\[64\] tdc0.w_dly_sig_n\[64\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6606 a_3962_15279# a_3689_15285# a_3877_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6607 a_11613_10633# _039_ a_11517_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6608 VPWR a_17635_2045# a_17803_1947# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6609 a_7733_10217# a_6743_9845# a_7607_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6610 tdc0.w_dly_sig\[80\] tdc0.w_dly_sig\[78\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6611 VPWR tdc0.w_dly_sig\[75\] tdc0.w_dly_sig\[77\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6612 VPWR tdc0.w_dly_sig\[122\] tdc0.w_dly_sig_n\[122\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6613 tdc0.w_dly_sig_n\[84\] tdc0.w_dly_sig\[84\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6614 VPWR a_11456_10927# uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X6615 a_5529_1679# a_5363_1679# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6616 a_5905_5487# tdc0.o_result\[67\] a_5823_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6618 tdc0.w_dly_sig_n\[21\] tdc0.w_dly_sig_n\[19\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6619 VPWR tdc0.w_dly_sig_n\[64\] tdc0.w_dly_sig\[65\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6620 VGND tdc0.w_dly_sig\[8\] tdc0.w_dly_sig_n\[8\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6621 a_8688_16745# a_8289_16373# a_8562_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6622 tdc0.w_dly_sig\[119\] tdc0.w_dly_sig\[117\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6623 VGND a_6579_17179# a_6537_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6624 a_9125_8751# tdc0.o_result\[33\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6625 VGND a_6871_8573# a_7039_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6626 VGND tdc0.w_dly_sig\[23\] tdc0.w_dly_sig_n\[23\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6627 tdc0.w_dly_sig\[13\] tdc0.w_dly_sig_n\[12\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6628 VGND tdc0.w_dly_sig\[86\] tdc0.w_dly_sig\[88\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6629 a_15833_10749# a_15299_10383# a_15738_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6630 VGND tdc0.w_dly_sig_n\[48\] tdc0.w_dly_sig_n\[50\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6631 VGND _002_ _009_ VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X6632 a_12459_17833# a_12330_17577# a_12039_17687# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6633 tdc0.o_result\[88\] a_7131_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6634 a_8527_10927# a_7829_10933# a_8270_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6635 a_12600_7119# a_12263_7119# a_12518_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6636 VPWR tdc0.w_dly_sig\[109\] tdc0.w_dly_sig\[111\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6637 VPWR tdc0.w_dly_sig_n\[89\] tdc0.w_dly_sig\[90\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6638 tdc0.w_dly_sig\[119\] tdc0.w_dly_sig_n\[118\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6639 VPWR a_3790_7119# clknet_4_1_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6640 VGND tdc0.w_dly_sig_n\[0\] tdc0.w_dly_sig_n\[2\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6642 a_14729_15285# a_14563_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6643 tdc0.w_dly_sig\[95\] tdc0.w_dly_sig_n\[94\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6644 a_2064_11305# a_1665_10933# a_1938_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6645 tdc0.w_dly_sig\[62\] tdc0.w_dly_sig\[60\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6646 a_15864_1679# a_15465_1679# a_15738_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6647 _090_ a_3247_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6648 a_12495_12247# a_12591_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6649 tdc0.w_dly_sig_n\[125\] tdc0.w_dly_sig_n\[123\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6650 VPWR tdc0.w_dly_sig_n\[70\] tdc0.w_dly_sig_n\[72\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6651 VGND _006_ a_12574_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6652 a_14507_14191# a_13809_14197# a_14250_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6653 VPWR net10 a_6273_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6654 VGND net4 a_12263_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X6655 clknet_4_14_0_clk a_17314_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6656 a_11786_13103# a_11539_13481# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6657 VPWR clk a_11058_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6658 a_17703_16745# a_17574_16489# a_17283_16599# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6659 VGND tdc0.w_dly_sig_n\[75\] tdc0.w_dly_sig\[76\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6662 VPWR clknet_4_8_0_clk a_11619_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6663 VGND a_11311_2741# a_11318_3041# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6664 tdc0.w_dly_sig_n\[45\] tdc0.w_dly_sig\[45\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6665 a_17950_16367# a_17703_16745# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6666 a_7442_3967# a_7274_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6667 tdc0.w_dly_sig\[5\] tdc0.w_dly_sig_n\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6668 a_18234_12292# a_18027_12233# a_18410_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6669 clknet_4_13_0_clk a_14388_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6670 tdc0.w_dly_sig\[121\] tdc0.w_dly_sig\[119\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6671 VPWR a_2071_11739# a_1987_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6672 clknet_4_9_0_clk a_14664_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6673 VGND a_4571_14013# a_4739_13915# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6674 tdc0.w_dly_sig_n\[89\] tdc0.w_dly_sig\[89\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6675 VGND tdc0.w_dly_sig_n\[66\] tdc0.w_dly_sig\[67\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6676 tdc0.w_dly_sig\[102\] tdc0.w_dly_sig\[100\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6677 tdc0.w_dly_sig_n\[16\] tdc0.w_dly_sig_n\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6678 tdc0.w_dly_sig\[23\] tdc0.w_dly_sig\[21\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6679 a_18163_12393# a_18027_12233# a_17743_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6680 tdc0.w_dly_sig_n\[15\] tdc0.w_dly_sig\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6681 a_5441_3855# tdc0.w_dly_sig\[87\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6682 VGND a_11490_6005# _026_ VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X6684 VGND tdc0.w_dly_sig\[7\] tdc0.w_dly_sig\[9\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6685 VPWR a_17555_6807# tdc0.o_result\[116\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6686 a_8009_8041# a_7019_7669# a_7883_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6687 tdc0.w_dly_sig_n\[9\] tdc0.w_dly_sig\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6688 tdc0.w_dly_sig\[36\] tdc0.w_dly_sig\[34\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6690 VGND a_5326_18111# a_5284_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6692 a_9677_4943# _019_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X6693 tdc0.w_dly_sig_n\[94\] tdc0.w_dly_sig_n\[92\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6694 tdc0.w_dly_sig_n\[25\] tdc0.w_dly_sig_n\[23\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6695 a_6495_17277# a_5713_16911# a_6411_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6697 a_7373_7663# tdc0.w_dly_sig\[36\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6698 a_12281_17455# a_11943_17687# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6699 VPWR _003_ a_9650_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X6700 VGND a_6395_12827# a_6353_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6701 VGND a_3348_13077# clknet_4_5_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6702 tdc0.w_dly_sig\[90\] tdc0.w_dly_sig_n\[89\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6703 VPWR tdc0.w_dly_sig\[125\] tdc0.w_dly_sig\[127\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6704 VGND tdc0.w_dly_sig\[42\] tdc0.w_dly_sig\[44\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R28 uio_oe[3] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6705 tdc0.w_dly_sig_n\[20\] tdc0.w_dly_sig\[20\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6708 VPWR tdc0.w_dly_sig_n\[106\] tdc0.w_dly_sig\[107\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6709 VPWR a_4295_1135# a_4463_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6710 a_3969_3311# tdc0.w_dly_sig\[84\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6711 a_4295_1135# a_3597_1141# a_4038_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6712 VGND tdc0.w_dly_sig_n\[59\] tdc0.w_dly_sig\[60\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6713 VPWR a_13783_18151# tdc0.o_result\[23\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6714 tdc0.w_dly_sig_n\[66\] tdc0.w_dly_sig_n\[64\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6715 tdc0.w_dly_sig_n\[72\] tdc0.w_dly_sig_n\[70\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6716 a_5434_7485# a_4995_7119# a_5349_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6717 a_13287_11305# a_13151_11145# a_12867_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6718 a_3026_17429# a_2858_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6719 tdc0.w_dly_sig\[94\] tdc0.w_dly_sig\[92\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6720 VPWR tdc0.w_dly_sig\[123\] tdc0.w_dly_sig\[125\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6721 clknet_4_1_0_clk a_3790_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6722 a_13795_10057# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6723 a_11892_11471# _056_ a_11504_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X6724 a_8933_1135# a_8399_1141# a_8838_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6725 VPWR a_15906_10495# a_15833_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6726 VPWR tdc0.w_dly_sig_n\[126\] tdc0.w_dly_sig\[127\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6727 a_9907_2045# a_9043_1679# a_9650_1791# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6729 a_8481_12809# tdc0.o_result\[120\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6730 VPWR tdc0.w_dly_sig\[121\] tdc0.w_dly_sig_n\[121\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6731 a_1485_13103# tdc0.w_dly_sig\[51\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6732 VPWR a_2255_15003# a_2171_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6733 tdc0.w_dly_sig_n\[7\] tdc0.w_dly_sig_n\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6734 a_14909_2601# a_13919_2229# a_14783_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6735 VGND a_9631_14191# a_9799_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6736 VPWR tdc0.w_dly_sig\[17\] a_7817_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6737 VPWR a_12649_7814# a_12318_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X6738 VGND _022_ a_2949_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6739 tdc0.o_result\[39\] a_9155_16341# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6740 tdc0.o_result\[119\] a_18171_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6741 VPWR a_14388_13621# clknet_4_13_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6742 tdc0.w_dly_sig\[38\] tdc0.w_dly_sig_n\[37\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6743 tdc0.w_dly_sig\[46\] tdc0.w_dly_sig\[44\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6744 VPWR tdc0.w_dly_sig\[21\] tdc0.w_dly_sig_n\[21\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6745 a_9209_13103# a_8675_13109# a_9114_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6746 tdc0.w_dly_sig\[91\] tdc0.w_dly_sig_n\[90\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6747 tdc0.w_dly_sig\[94\] tdc0.w_dly_sig_n\[93\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6748 a_11610_13380# a_11403_13321# a_11786_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6749 VGND a_15906_1791# a_15864_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6750 tdc0.w_dly_sig\[76\] tdc0.w_dly_sig\[74\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6751 VGND tdc0.w_dly_sig\[121\] a_18581_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6752 VPWR a_16578_13103# clknet_4_15_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6753 a_16639_14709# a_16930_15009# a_16881_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6755 a_12199_4631# tdc0.o_result\[97\] a_12345_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X6756 a_1393_9295# tdc0.w_dly_sig\[76\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6757 VGND _094_ a_16127_7779# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X6758 tdc0.w_dly_sig_n\[64\] tdc0.w_dly_sig\[64\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6759 a_18003_9661# a_17305_9295# a_17746_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6761 VGND a_17635_2045# a_17803_1947# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6762 tdc0.w_dly_sig_n\[63\] tdc0.w_dly_sig\[63\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6763 a_13070_8207# a_12893_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X6764 a_11539_13481# a_11403_13321# a_11119_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6765 tdc0.w_dly_sig\[84\] tdc0.w_dly_sig\[82\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6766 VPWR a_17647_3543# tdc0.o_result\[112\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6767 VGND a_9431_16091# a_9389_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6768 a_4563_3311# a_3781_3317# a_4479_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6769 VGND tdc0.w_dly_sig_n\[95\] tdc0.w_dly_sig\[96\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6770 VPWR a_11311_2741# a_11318_3041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6772 tdc0.w_dly_sig\[126\] tdc0.w_dly_sig\[124\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6773 a_17865_8207# _015_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X6774 tdc0.w_dly_sig_n\[33\] tdc0.w_dly_sig_n\[31\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6775 VPWR clknet_4_0_0_clk a_1683_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6776 a_2593_10383# tdc0.o_result\[75\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6777 VGND clknet_4_8_0_clk a_13459_1141# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6778 a_15646_18365# a_15373_17999# a_15561_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6779 VGND tdc0.w_dly_sig_n\[87\] tdc0.w_dly_sig_n\[89\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6780 VGND tdc0.w_dly_sig_n\[69\] tdc0.w_dly_sig\[70\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6781 VGND tdc0.w_dly_sig_n\[100\] tdc0.w_dly_sig_n\[102\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6782 VPWR tdc0.w_dly_sig\[18\] tdc0.w_dly_sig\[20\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6783 VPWR tdc0.w_dly_sig_n\[80\] tdc0.w_dly_sig_n\[82\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6784 VPWR tdc0.w_dly_sig\[7\] a_14349_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6785 a_12345_4399# _025_ a_12199_4631# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X6786 clknet_4_6_0_clk a_6550_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6787 clknet_4_11_0_clk a_16762_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6788 VGND tdc0.w_dly_sig\[38\] tdc0.w_dly_sig\[40\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6789 VGND a_12999_591# net2 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6790 tdc0.w_dly_sig_n\[94\] tdc0.w_dly_sig\[94\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6791 tdc0.w_dly_sig\[106\] tdc0.w_dly_sig\[104\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6792 VGND tdc0.w_dly_sig_n\[123\] tdc0.w_dly_sig\[124\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6793 tdc0.w_dly_sig\[8\] tdc0.w_dly_sig\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6794 a_13082_12292# a_12875_12233# a_13258_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6795 a_6687_12015# a_5989_12021# a_6430_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6796 VGND a_6411_17277# a_6579_17179# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6797 VGND a_8435_8751# a_8603_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6798 a_10239_10633# _026_ a_10321_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6799 uo_out[3] a_16332_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6800 a_9071_16367# a_8289_16373# a_8987_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6801 VPWR a_8270_10901# a_8197_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6802 tdc0.w_dly_sig_n\[72\] tdc0.w_dly_sig\[72\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6803 VGND _064_ a_15575_6281# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X6804 VPWR tdc0.w_dly_sig_n\[49\] tdc0.w_dly_sig_n\[51\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6806 a_13011_12393# a_12875_12233# a_12591_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6807 tdc0.o_result\[24\] a_15595_17429# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6808 a_1830_9813# a_1662_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6809 VGND tdc0.w_dly_sig_n\[52\] tdc0.w_dly_sig_n\[54\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6810 tdc0.w_dly_sig_n\[43\] tdc0.w_dly_sig\[43\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6811 a_1987_9661# a_1205_9295# a_1903_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6812 a_5560_7119# a_5161_7119# a_5434_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6813 tdc0.w_dly_sig\[99\] tdc0.w_dly_sig_n\[98\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6814 a_8661_17455# tdc0.w_dly_sig\[18\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6815 VPWR net10 a_7653_17161# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6816 VGND a_11023_13335# tdc0.o_result\[13\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6818 a_4111_18365# a_3413_17999# a_3854_18111# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6819 tdc0.w_dly_sig_n\[83\] tdc0.w_dly_sig\[83\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6820 a_3689_15285# a_3523_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6821 a_14786_9071# tdc0.o_result\[4\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X6822 tdc0.w_dly_sig\[128\] tdc0.w_dly_sig\[126\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6823 VPWR a_13690_7895# _004_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X6824 clknet_4_15_0_clk a_16578_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6825 a_14664_6005# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6826 VPWR a_14186_3829# a_14115_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6827 a_16819_10535# a_16915_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6828 tdc0.w_dly_sig_n\[81\] tdc0.w_dly_sig\[81\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6829 VPWR _025_ a_15853_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6830 a_4866_13077# a_4698_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6831 VGND a_16332_9839# uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6833 net7 a_11027_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6834 _096_ a_16127_7779# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6836 a_8481_11721# tdc0.o_result\[123\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6837 VGND a_7263_17673# a_7270_17577# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6839 VGND a_16331_10651# a_16289_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6840 a_11490_6005# a_11343_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X6841 a_4617_8751# tdc0.o_result\[81\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6842 VPWR tdc0.w_dly_sig_n\[18\] tdc0.w_dly_sig\[19\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6844 tdc0.w_dly_sig_n\[79\] tdc0.w_dly_sig\[79\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6845 VGND a_7987_4631# tdc0.o_result\[108\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6846 VGND clknet_0_clk a_3698_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6848 tdc0.o_result\[78\] a_2623_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6849 tdc0.w_dly_sig_n\[34\] tdc0.w_dly_sig_n\[32\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6850 VGND _019_ a_10769_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6851 clknet_4_12_0_clk a_12548_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6852 VGND a_17406_4917# a_17335_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6853 VGND tdc0.w_dly_sig_n\[79\] tdc0.w_dly_sig_n\[81\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6854 VGND tdc0.w_dly_sig_n\[81\] tdc0.w_dly_sig_n\[83\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6855 _050_ a_11527_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6856 a_6883_17687# a_6979_17687# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6857 a_6905_6953# a_5915_6581# a_6779_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6858 a_15511_17455# a_14729_17461# a_15427_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6859 VPWR tdc0.w_dly_sig\[27\] tdc0.w_dly_sig\[29\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6860 tdc0.w_dly_sig\[71\] tdc0.w_dly_sig_n\[70\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6861 a_14445_8867# _011_ a_14373_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6862 VPWR a_16155_6183# _063_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X6863 tdc0.w_dly_sig_n\[0\] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6864 a_13863_5487# a_13165_5493# a_13606_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6865 VGND clknet_4_2_0_clk a_6927_1141# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6866 _356_.X a_16732_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X6867 VPWR tdc0.w_dly_sig\[73\] tdc0.w_dly_sig\[75\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6868 tdc0.w_dly_sig_n\[120\] tdc0.w_dly_sig_n\[118\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6869 VGND tdc0.w_dly_sig\[8\] a_13429_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6870 a_16301_17775# _007_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X6871 VPWR tdc0.w_dly_sig_n\[3\] tdc0.w_dly_sig_n\[5\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6872 VPWR a_6503_14013# a_6671_13915# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6873 clknet_4_7_0_clk a_7856_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6874 a_13695_3829# a_13979_3829# a_13914_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6875 a_8573_5487# tdc0.o_result\[32\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6876 VPWR net6 a_9125_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6877 a_14186_14709# a_13986_15009# a_14335_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6878 a_15128_4777# a_14729_4405# a_15002_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6879 clknet_0_clk a_11058_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6880 a_5253_14735# a_5087_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6881 a_6191_17455# _029_ a_6273_17775# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6882 clknet_0_clk a_11058_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6883 a_2585_17461# a_2419_17461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6884 VPWR a_11839_2045# a_12007_1947# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6885 a_14082_6575# a_13643_6581# a_13997_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6886 a_9747_8181# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0746 pd=0.775 as=0.0777 ps=0.79 w=0.42 l=0.15
X6887 VPWR tdc0.w_dly_sig\[57\] tdc0.w_dly_sig_n\[57\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6888 VGND a_16578_13103# clknet_4_15_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6889 VPWR tdc0.w_dly_sig\[75\] tdc0.w_dly_sig_n\[75\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6890 VPWR net4 a_13183_6583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X6891 a_6550_13103# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X6892 a_7699_4221# a_6835_3855# a_7442_3967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6893 tdc0.w_dly_sig\[9\] tdc0.w_dly_sig_n\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6894 a_17843_14409# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6895 VGND tdc0.o_result\[0\] a_16166_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6896 VPWR tdc0.w_dly_sig\[119\] a_18673_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6897 a_12118_9295# tdc0.o_result\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X6898 VGND tdc0.w_dly_sig_n\[51\] tdc0.w_dly_sig\[52\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6899 a_17463_14423# a_17559_14423# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6900 a_16155_6183# tdc0.o_result\[104\] a_16301_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R29 uio_out[4] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6901 a_7399_17833# a_7270_17577# a_6979_17687# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6902 a_1554_11989# a_1386_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6903 a_7646_17455# a_7399_17833# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6904 a_11685_10633# _038_ a_11613_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6905 VGND clknet_4_5_0_clk a_4167_17461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6906 a_14786_9071# _018_ a_14952_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6907 a_18255_8041# a_18126_7785# a_17835_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6908 a_11290_11247# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6909 a_9715_14191# a_8933_14197# a_9631_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6910 tdc0.w_dly_sig\[26\] tdc0.w_dly_sig_n\[25\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6911 a_9459_4631# a_9555_4631# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6912 tdc0.w_dly_sig_n\[39\] tdc0.w_dly_sig\[39\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6914 net1 a_18187_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6915 a_10527_14735# a_10398_15009# a_10107_14709# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6916 VGND a_4555_15253# a_4513_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6917 a_14729_4405# a_14563_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6918 tdc0.w_dly_sig_n\[91\] tdc0.w_dly_sig\[91\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6919 a_7097_3311# tdc0.w_dly_sig\[91\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6920 tdc0.w_dly_sig_n\[92\] tdc0.w_dly_sig\[92\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6921 a_1757_16911# a_1591_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6923 net28 a_12574_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6924 a_6725_2229# a_6559_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6925 VPWR a_14157_4917# _017_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6926 VGND tdc0.w_dly_sig\[27\] tdc0.w_dly_sig_n\[27\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6927 tdc0.w_dly_sig\[106\] tdc0.w_dly_sig_n\[105\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6929 VGND _002_ a_11987_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6931 tdc0.w_dly_sig_n\[121\] tdc0.w_dly_sig_n\[119\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6932 tdc0.w_dly_sig\[42\] tdc0.w_dly_sig\[40\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6933 VGND tdc0.w_dly_sig_n\[30\] tdc0.w_dly_sig\[31\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6934 VGND tdc0.w_dly_sig_n\[47\] tdc0.w_dly_sig\[48\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6935 a_11241_4943# a_11154_5095# a_11159_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
X6936 a_8565_1141# a_8399_1141# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6938 VPWR tdc0.w_dly_sig_n\[16\] tdc0.w_dly_sig_n\[18\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6939 VPWR clknet_4_2_0_clk a_6099_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6940 a_16166_12335# _066_ a_16332_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6941 VGND a_4019_5487# a_4187_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6942 tdc0.w_dly_sig_n\[112\] tdc0.w_dly_sig_n\[110\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6943 VPWR tdc0.w_dly_sig_n\[78\] tdc0.w_dly_sig_n\[80\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6944 tdc0.w_dly_sig_n\[106\] tdc0.w_dly_sig\[106\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6945 VGND a_6706_4373# a_6664_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6946 VPWR a_18187_10901# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6947 VPWR tdc0.w_dly_sig_n\[8\] tdc0.w_dly_sig_n\[10\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6948 VPWR tdc0.w_dly_sig_n\[101\] tdc0.w_dly_sig\[102\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6949 a_11057_8751# tdc0.o_result\[65\] a_10975_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6950 VGND tdc0.w_dly_sig_n\[50\] tdc0.w_dly_sig_n\[52\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6951 VGND tdc0.w_dly_sig\[116\] tdc0.w_dly_sig_n\[116\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6952 tdc0.w_dly_sig\[10\] tdc0.w_dly_sig_n\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6953 VPWR tdc0.w_dly_sig\[112\] a_10393_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6954 VPWR tdc0.w_dly_sig_n\[101\] tdc0.w_dly_sig_n\[103\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6955 tdc0.o_result\[98\] a_13479_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6956 a_12567_4221# a_11785_3855# a_12483_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6957 a_15653_1679# tdc0.w_dly_sig\[105\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6958 a_7221_17455# a_6883_17687# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6959 a_8454_11989# a_8286_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6960 a_9665_12335# tdc0.o_result\[17\] a_9319_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6961 VGND a_9891_18267# a_9849_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6962 tdc0.w_dly_sig\[5\] tdc0.w_dly_sig\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6963 VGND tdc0.w_dly_sig\[41\] tdc0.w_dly_sig\[43\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6964 clknet_4_10_0_clk a_16412_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6965 a_11609_4719# tdc0.o_result\[78\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6966 VPWR a_14952_8751# uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6967 VPWR a_14664_6005# clknet_4_9_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6968 tdc0.w_dly_sig\[18\] tdc0.w_dly_sig_n\[17\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6970 VPWR a_10423_591# net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6971 a_16117_8207# tdc0.o_result\[107\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6973 a_11701_8867# _075_ a_11619_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X6974 a_8286_12015# a_8013_12021# a_8201_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6975 tdc0.w_dly_sig_n\[12\] tdc0.w_dly_sig_n\[10\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6976 uo_out[0] a_16332_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6977 a_11957_12393# a_11403_12233# a_11610_12292# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6978 VGND a_7166_2197# a_7124_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6979 a_14208_6953# a_13809_6581# a_14082_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6982 clknet_4_3_0_clk a_7286_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6984 a_7182_9839# a_6743_9845# a_7097_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6985 a_1665_10933# a_1499_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6986 a_13695_14709# a_13986_15009# a_13937_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6987 a_5253_14735# a_5087_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6988 a_15887_15101# a_15189_14735# a_15630_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6989 a_6273_17455# tdc0.o_result\[18\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6990 VPWR clknet_4_15_0_clk a_15207_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6991 _018_ a_14195_8867# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X6992 tdc0.o_result\[55\] a_4463_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6993 VGND _022_ a_3593_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6994 VGND a_14388_13621# clknet_4_13_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6995 VPWR tdc0.w_dly_sig\[119\] tdc0.w_dly_sig_n\[119\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6996 tdc0.w_dly_sig_n\[22\] tdc0.w_dly_sig_n\[20\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6997 a_2631_3133# a_1849_2767# a_2547_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6998 a_7470_17732# a_7263_17673# a_7646_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6999 VGND tdc0.w_dly_sig_n\[73\] tdc0.w_dly_sig\[74\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7000 VGND tdc0.w_dly_sig_n\[114\] tdc0.w_dly_sig\[115\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7001 VPWR a_10759_8181# _005_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7002 VGND tdc0.w_dly_sig\[48\] tdc0.w_dly_sig_n\[48\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7003 a_4655_14013# a_3873_13647# a_4571_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7004 a_3686_18365# a_3247_17999# a_3601_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7005 a_4839_2045# a_4057_1679# a_4755_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7006 VPWR tdc0.w_dly_sig\[10\] tdc0.w_dly_sig\[12\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7007 a_17485_1513# a_16495_1141# a_17359_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7008 tdc0.w_dly_sig\[46\] tdc0.w_dly_sig_n\[45\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7009 _093_ a_16035_8457# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X7010 tdc0.w_dly_sig\[96\] tdc0.w_dly_sig\[94\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7011 _069_ a_8399_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X7012 a_13809_6581# a_13643_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7013 tdc0.w_dly_sig_n\[8\] tdc0.w_dly_sig\[8\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7014 VGND tdc0.w_dly_sig_n\[42\] tdc0.w_dly_sig_n\[44\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7015 VGND tdc0.w_dly_sig\[117\] tdc0.w_dly_sig_n\[117\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7016 VPWR tdc0.w_dly_sig\[127\] a_17661_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7017 VGND tdc0.w_dly_sig\[77\] tdc0.w_dly_sig\[79\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7018 VGND a_11839_2045# a_12007_1947# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7019 VGND a_9263_1135# a_9431_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7020 tdc0.w_dly_sig_n\[4\] tdc0.w_dly_sig_n\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7021 a_4149_3311# a_3615_3317# a_4054_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7022 a_9366_10071# _079_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X7023 VGND a_17774_16644# a_17703_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X7024 tdc0.w_dly_sig\[54\] tdc0.w_dly_sig_n\[53\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7025 VPWR tdc0.w_dly_sig\[3\] tdc0.w_dly_sig_n\[3\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7026 a_6706_4373# a_6538_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7027 a_13091_7779# _048_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7028 a_10029_6575# _001_ a_9779_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7029 a_14299_17999# a_14170_18273# a_13879_17973# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7030 a_15473_13647# net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X7031 VPWR a_11780_7637# a_11122_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=2.12 as=0.165 ps=1.33 w=1 l=0.15
X7032 tdc0.w_dly_sig_n\[120\] tdc0.w_dly_sig\[120\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7034 clknet_4_14_0_clk a_17314_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7035 VPWR a_17378_1791# a_17305_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7036 a_12801_2223# tdc0.w_dly_sig\[99\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7037 tdc0.w_dly_sig\[66\] tdc0.w_dly_sig_n\[65\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7038 VPWR a_14611_13335# tdc0.o_result\[2\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7039 a_1662_15101# a_1389_14735# a_1577_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7040 tdc0.w_dly_sig_n\[11\] tdc0.w_dly_sig_n\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7041 clknet_4_13_0_clk a_14388_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7042 VPWR a_2071_9563# a_1987_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7043 a_6909_9845# a_6743_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7044 a_5970_1791# a_5802_2045# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7045 VPWR a_14158_8319# a_14085_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7046 VPWR tdc0.w_dly_sig\[19\] tdc0.w_dly_sig\[21\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7047 a_9347_1135# a_8565_1141# a_9263_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7048 a_4379_10927# a_3597_10933# a_4295_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7049 VPWR tdc0.w_dly_sig\[107\] tdc0.w_dly_sig_n\[107\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7050 _002_ a_13183_6583# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X7051 VPWR tdc0.w_dly_sig_n\[21\] tdc0.w_dly_sig\[22\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7052 VGND a_12631_591# net4 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7053 VPWR tdc0.w_dly_sig_n\[74\] tdc0.w_dly_sig\[75\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7054 a_3965_1135# a_3431_1141# a_3870_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7055 VGND _001_ _019_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7056 VPWR _012_ a_9677_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7057 VGND a_13082_12292# a_13011_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X7058 VGND tdc0.w_dly_sig\[84\] tdc0.w_dly_sig\[86\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7059 tdc0.w_dly_sig_n\[128\] tdc0.w_dly_sig\[128\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7060 a_16589_14511# _012_ a_16155_14423# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7061 VPWR a_4176_6005# clknet_4_0_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7062 VPWR a_2087_15101# a_2255_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7063 a_7189_6031# tdc0.w_dly_sig\[33\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7064 a_11122_7637# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.175 ps=1.35 w=1 l=0.15
X7065 a_17743_12247# a_18034_12137# a_17985_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7067 VPWR tdc0.w_dly_sig_n\[0\] tdc0.w_dly_sig\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7068 a_4245_4399# tdc0.w_dly_sig\[68\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7069 VPWR tdc0.w_dly_sig_n\[25\] tdc0.w_dly_sig_n\[27\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7070 VPWR net28 a_10321_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7071 VPWR tdc0.w_dly_sig\[1\] a_16741_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7073 VPWR tdc0.o_result\[69\] a_9677_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X7075 a_14851_15823# a_14715_15797# a_14431_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7076 tdc0.w_dly_sig_n\[82\] tdc0.w_dly_sig\[82\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7077 tdc0.w_dly_sig\[86\] tdc0.w_dly_sig_n\[85\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7078 VPWR a_8500_4917# clknet_4_2_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7079 VPWR clknet_4_0_0_clk a_1683_1141# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7080 tdc0.w_dly_sig_n\[118\] tdc0.w_dly_sig\[118\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7081 VGND a_2439_6549# a_2397_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7082 a_17567_16585# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7083 VPWR a_7867_4123# a_7783_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7084 a_6043_5309# a_5345_4943# a_5786_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7085 VPWR a_16762_8207# clknet_4_11_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7088 a_6909_9845# a_6743_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7089 VGND clknet_0_clk a_12548_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X7090 a_7561_13103# tdc0.o_result\[36\] a_7479_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7091 VGND net8 a_16022_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X7092 VPWR _012_ a_11333_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7093 tdc0.w_dly_sig_n\[87\] tdc0.w_dly_sig\[87\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7094 VPWR a_11058_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7095 VGND a_14507_6575# a_14675_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7096 VPWR a_12376_8751# uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7097 a_13459_8751# _010_ a_13541_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7098 tdc0.w_dly_sig\[56\] tdc0.w_dly_sig_n\[55\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7099 tdc0.w_dly_sig_n\[117\] tdc0.w_dly_sig_n\[115\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7100 VPWR a_17935_6793# a_17942_6697# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7101 VPWR tdc0.w_dly_sig\[72\] tdc0.w_dly_sig_n\[72\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7102 a_2581_9129# a_1591_8757# a_2455_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7103 a_5583_18365# a_4719_17999# a_5326_18111# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7104 VPWR tdc0.w_dly_sig_n\[13\] tdc0.w_dly_sig_n\[15\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7105 a_4425_13109# a_4259_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7106 VGND a_3026_17429# a_2984_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7107 VGND _025_ a_9389_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X7108 net6 a_8819_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7109 a_18326_4676# a_18126_4521# a_18475_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7110 a_14273_2223# tdc0.w_dly_sig\[97\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7111 VGND tdc0.w_dly_sig_n\[52\] tdc0.w_dly_sig\[53\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7112 a_17305_2045# a_16771_1679# a_17210_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7113 VPWR _023_ a_8573_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7115 VPWR a_8987_16367# a_9155_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7116 a_11361_12015# a_11023_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X7117 VPWR tdc0.w_dly_sig_n\[108\] tdc0.w_dly_sig_n\[110\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7118 _099_ a_8399_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X7119 a_9411_12809# _013_ a_9493_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7120 a_5253_18365# a_4719_17999# a_5158_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7121 tdc0.w_dly_sig\[25\] tdc0.w_dly_sig\[23\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7122 VPWR tdc0.w_dly_sig\[7\] tdc0.w_dly_sig_n\[7\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7123 VGND a_8987_16367# a_9155_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7124 a_11923_2045# a_11141_1679# a_11839_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7125 VGND _005_ a_11892_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7126 VPWR clknet_0_clk a_16578_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7127 a_14085_8573# a_13551_8207# a_13990_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7128 VPWR tdc0.w_dly_sig_n\[26\] tdc0.w_dly_sig_n\[28\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7129 VGND tdc0.w_dly_sig\[114\] tdc0.w_dly_sig_n\[114\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7130 VGND a_15106_9269# a_15035_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X7131 VPWR tdc0.w_dly_sig_n\[39\] tdc0.w_dly_sig\[40\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R30 VPWR tt_um_hpretl_tt06_tdc_19.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7132 VPWR _046_ a_12644_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X7133 VGND tdc0.w_dly_sig\[26\] a_15269_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7134 a_1849_2767# a_1683_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7135 VGND tdc0.w_dly_sig_n\[57\] tdc0.w_dly_sig\[58\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7136 a_11269_3133# a_10931_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X7138 VGND tdc0.w_dly_sig_n\[20\] tdc0.w_dly_sig\[21\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7139 a_18613_9071# _025_ a_18179_8983# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7140 a_18119_7881# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7141 VPWR clknet_4_0_0_clk a_1591_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7142 a_7925_8751# tdc0.w_dly_sig\[34\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7143 a_7653_17161# tdc0.o_result\[16\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X7144 VGND clknet_4_13_0_clk a_13643_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7145 a_2455_17277# a_1591_16911# a_2198_17023# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7146 VGND a_2198_17023# a_2156_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7147 VGND clknet_4_1_0_clk a_4167_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7148 VGND net3 _023_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7149 a_8017_10927# tdc0.w_dly_sig\[62\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7150 VGND tdc0.w_dly_sig\[6\] a_13705_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7151 VPWR tdc0.w_dly_sig\[8\] tdc0.w_dly_sig\[10\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7152 a_17979_14569# a_17843_14409# a_17559_14423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7153 a_17283_16599# a_17574_16489# a_17525_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7154 tdc0.w_dly_sig\[129\] tdc0.w_dly_sig\[127\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7155 a_6453_4399# tdc0.w_dly_sig\[89\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7156 a_15553_15657# a_14563_15285# a_15427_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7157 a_9747_8181# _003_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.28 ps=1.62 w=0.42 l=0.15
X7158 a_10975_8751# net7 a_11057_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7159 a_8964_15823# a_8565_15823# a_8838_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7160 a_11806_7119# a_11067_7119# a_11692_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.137 ps=1.07 w=0.65 l=0.15
X7161 a_16967_7119# a_16838_7393# a_16547_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7162 tdc0.o_result\[11\] a_14583_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7163 tdc0.w_dly_sig_n\[13\] tdc0.w_dly_sig_n\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7164 tdc0.o_result\[32\] a_7867_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7165 _051_ a_13091_7779# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X7166 VGND tdc0.w_dly_sig_n\[127\] tdc0.w_dly_sig\[128\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7167 VPWR a_7959_1109# a_7875_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7168 VPWR net5 a_11642_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7169 a_3854_14847# a_3686_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7170 a_2949_3689# a_1959_3317# a_2823_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7172 VPWR tdc0.w_dly_sig\[92\] tdc0.w_dly_sig\[94\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7173 tdc0.w_dly_sig\[20\] tdc0.w_dly_sig\[18\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7174 a_18326_4676# a_18119_4617# a_18502_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7175 _006_ net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X7177 VPWR tdc0.w_dly_sig_n\[70\] tdc0.w_dly_sig\[71\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7178 VPWR a_7856_14165# clknet_4_7_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7179 tdc0.w_dly_sig_n\[8\] tdc0.w_dly_sig_n\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7180 tdc0.w_dly_sig\[124\] tdc0.w_dly_sig_n\[123\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7181 VPWR a_7883_7663# a_8051_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7182 VGND tdc0.w_dly_sig_n\[14\] tdc0.w_dly_sig\[15\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7184 tdc0.w_dly_sig\[83\] tdc0.w_dly_sig\[81\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7185 VGND _025_ a_16484_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7186 _000_ a_10515_7671# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7187 a_4774_17429# a_4606_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7188 a_10055_2223# _028_ a_10137_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7189 VGND tdc0.w_dly_sig\[83\] tdc0.w_dly_sig\[85\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7190 a_15853_7983# _025_ a_15419_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7192 tdc0.w_dly_sig_n\[105\] tdc0.w_dly_sig\[105\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7193 a_17578_9661# a_17139_9295# a_17493_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7194 tdc0.w_dly_sig_n\[51\] tdc0.w_dly_sig_n\[49\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7195 VGND a_2991_3285# a_2949_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7196 a_9555_4631# a_9846_4521# a_9797_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7197 tdc0.w_dly_sig\[108\] tdc0.w_dly_sig\[106\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7198 tdc0.w_dly_sig\[112\] tdc0.w_dly_sig_n\[111\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7199 VGND net28 a_11413_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X7200 a_17774_13621# a_17567_13621# a_17950_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7201 VGND tdc0.w_dly_sig_n\[83\] tdc0.w_dly_sig\[84\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7202 a_16412_6549# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7203 VPWR a_16055_15003# a_15971_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7204 tdc0.w_dly_sig_n\[31\] tdc0.w_dly_sig_n\[29\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7205 _007_ a_9747_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7206 tdc0.w_dly_sig_n\[10\] tdc0.w_dly_sig\[10\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7207 tdc0.w_dly_sig_n\[34\] tdc0.w_dly_sig\[34\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7208 VPWR a_5326_18111# a_5253_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7209 a_18673_4777# a_18119_4617# a_18326_4676# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7210 VGND tdc0.w_dly_sig\[95\] tdc0.w_dly_sig\[97\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7211 VPWR tdc0.w_dly_sig_n\[76\] tdc0.w_dly_sig_n\[78\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7212 VGND a_2106_10901# a_2064_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7213 VGND tdc0.w_dly_sig_n\[47\] tdc0.w_dly_sig_n\[49\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7214 VPWR a_4279_18267# a_4195_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7215 uo_out[3] a_16332_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7216 a_18581_3689# a_18034_3433# a_18234_3588# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X7217 tdc0.w_dly_sig\[14\] tdc0.w_dly_sig\[12\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7218 clknet_4_0_0_clk a_4176_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7219 a_9757_3855# a_8767_3855# a_9631_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7220 a_12877_17833# a_12330_17577# a_12530_17732# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X7221 VPWR tdc0.w_dly_sig\[96\] tdc0.w_dly_sig\[98\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7222 VGND a_17199_4917# a_17206_5217# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7223 a_7166_2197# a_6998_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7224 VPWR a_16332_9839# uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7225 VPWR clknet_4_2_0_clk a_6743_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7226 VGND tdc0.w_dly_sig\[16\] a_10945_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7227 a_15864_10383# a_15465_10383# a_15738_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7228 a_2708_14569# a_2309_14197# a_2582_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7229 VPWR a_12530_17732# a_12459_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X7230 a_17739_7895# a_17835_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7231 a_1849_2767# a_1683_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7232 clknet_4_8_0_clk a_12548_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7233 VGND tdc0.w_dly_sig\[60\] tdc0.w_dly_sig_n\[60\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7236 VPWR clknet_4_1_0_clk a_1039_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7238 VGND a_11490_6005# _026_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7239 a_18502_4399# a_18255_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7240 clknet_0_clk a_11058_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7241 a_15427_17455# a_14563_17461# a_15170_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7242 a_6975_17999# a_6755_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X7243 tdc0.w_dly_sig_n\[18\] tdc0.w_dly_sig_n\[16\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7244 VPWR clknet_4_9_0_clk a_14563_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7245 VGND net1 tdc0.w_dly_sig_n\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7246 a_4606_17455# a_4167_17461# a_4521_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7247 VGND net11 a_14909_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X7248 VGND tdc0.w_dly_sig\[108\] tdc0.w_dly_sig_n\[108\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7250 a_16247_10749# a_15465_10383# a_16163_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7251 tdc0.w_dly_sig\[75\] tdc0.w_dly_sig\[73\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7252 a_11058_9839# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7253 a_7458_7663# a_7185_7669# a_7373_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7254 a_2217_1135# a_1683_1141# a_2122_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7255 tdc0.w_dly_sig_n\[61\] tdc0.w_dly_sig_n\[59\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7256 VPWR tdc0.w_dly_sig\[35\] tdc0.w_dly_sig\[37\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7257 VGND tdc0.w_dly_sig\[50\] tdc0.w_dly_sig\[52\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7258 a_15097_17455# a_14563_17461# a_15002_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7259 VGND tdc0.w_dly_sig_n\[84\] tdc0.w_dly_sig_n\[86\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7260 a_16951_5487# net8 a_16733_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7261 a_6173_8207# a_6007_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7262 VPWR a_6027_7387# a_5943_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7263 a_6619_17973# clknet_4_7_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7264 VGND tdc0.w_dly_sig\[123\] tdc0.w_dly_sig_n\[123\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7265 VGND clknet_4_5_0_clk a_5087_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7266 tdc0.w_dly_sig\[96\] tdc0.w_dly_sig_n\[95\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7267 a_8481_12559# tdc0.o_result\[56\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7268 VPWR a_13054_2197# a_12981_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7269 a_3597_1141# a_3431_1141# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7270 a_7987_4631# a_8083_4631# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7271 a_3348_13077# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7272 a_15814_18111# a_15646_18365# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7273 a_17704_9295# a_17305_9295# a_17578_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7274 a_17306_15101# a_17059_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7275 VGND tdc0.w_dly_sig_n\[38\] tdc0.w_dly_sig\[39\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7276 VGND clknet_4_6_0_clk a_5823_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7278 VGND a_17843_14409# a_17850_14313# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7279 VGND tdc0.w_dly_sig_n\[113\] tdc0.w_dly_sig\[114\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7280 a_6577_18365# a_6239_18151# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X7281 tdc0.w_dly_sig_n\[89\] tdc0.w_dly_sig_n\[87\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7282 a_12134_6549# a_11987_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X7283 VGND a_12518_7119# _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X7284 a_1738_13077# a_1570_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7286 VGND tdc0.w_dly_sig_n\[104\] tdc0.w_dly_sig\[105\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7287 a_10321_8751# tdc0.o_result\[94\] a_10239_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7288 VGND a_4187_5461# a_4145_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7289 a_15825_6281# _063_ a_15753_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7290 clknet_4_2_0_clk a_8500_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7291 a_1830_9813# a_1662_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7292 VGND a_13783_18151# tdc0.o_result\[23\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7293 a_9965_4943# _020_ a_9531_5095# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7294 VGND tdc0.w_dly_sig_n\[22\] tdc0.w_dly_sig\[23\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7295 VPWR tdc0.w_dly_sig\[45\] tdc0.w_dly_sig_n\[45\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7296 a_6963_4399# a_6099_4405# a_6706_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7297 tdc0.w_dly_sig\[73\] tdc0.w_dly_sig_n\[72\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7298 a_13438_5487# a_12999_5493# a_13353_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7299 VGND a_1903_11837# a_2071_11739# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7300 VGND clknet_4_0_0_clk a_5087_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7301 VPWR tdc0.w_dly_sig_n\[32\] tdc0.w_dly_sig\[33\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7302 _043_ a_11067_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7303 a_4605_3689# a_3615_3317# a_4479_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7304 a_3873_4943# a_3707_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7305 VPWR a_18187_10901# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7306 tdc0.o_result\[52\] a_4739_13915# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7307 a_4038_10901# a_3870_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7308 VGND a_3790_7119# clknet_4_1_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X7309 VGND a_7350_9813# a_7308_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7310 tdc0.w_dly_sig_n\[9\] tdc0.w_dly_sig_n\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7311 VPWR tdc0.w_dly_sig\[31\] tdc0.w_dly_sig_n\[31\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7312 a_6081_6581# a_5915_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7314 tdc0.w_dly_sig_n\[27\] tdc0.w_dly_sig\[27\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7315 VPWR tdc0.w_dly_sig\[115\] tdc0.w_dly_sig\[117\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7316 a_11251_15279# _029_ a_11333_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7318 a_16301_14191# _012_ a_16155_14423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X7319 VPWR a_10091_3311# a_10259_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7321 a_12318_7637# net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X7322 tdc0.w_dly_sig\[48\] tdc0.w_dly_sig_n\[47\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7323 a_7350_9813# a_7182_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7324 a_10975_17455# _029_ a_11057_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7325 a_11447_2767# a_11311_2741# a_11027_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7326 uo_out[1] a_12284_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X7327 clknet_4_10_0_clk a_16412_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X7328 a_16332_12015# _071_ a_16166_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7329 a_15170_15253# a_15002_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7330 a_12609_3855# a_11619_3855# a_12483_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7331 a_12649_7814# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X7332 tdc0.w_dly_sig\[98\] tdc0.w_dly_sig\[96\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7333 tdc0.w_dly_sig_n\[10\] tdc0.w_dly_sig_n\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7334 tdc0.w_dly_sig\[126\] tdc0.w_dly_sig_n\[125\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7335 a_17477_14735# a_16923_14709# a_17130_14709# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7336 a_15381_5807# net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X7337 tdc0.w_dly_sig\[72\] tdc0.w_dly_sig\[70\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7338 tdc0.w_dly_sig\[57\] tdc0.w_dly_sig_n\[56\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7339 a_6078_14013# a_5639_13647# a_5993_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7340 net5 a_11711_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X7341 _094_ a_16022_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7342 a_3413_17999# a_3247_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7343 a_11290_11247# _036_ a_11456_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7344 tdc0.w_dly_sig\[112\] tdc0.w_dly_sig\[110\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7345 a_14676_12809# _091_ a_14944_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7346 tdc0.w_dly_sig\[43\] tdc0.w_dly_sig\[41\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7347 a_17979_14569# a_17850_14313# a_17559_14423# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7348 a_1945_4399# tdc0.w_dly_sig\[79\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7349 VGND a_4295_1135# a_4463_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7350 a_17703_13647# a_17574_13921# a_17283_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7351 a_16600_12015# _066_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7352 a_17130_14709# a_16923_14709# a_17306_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7353 VGND tdc0.w_dly_sig\[79\] tdc0.w_dly_sig_n\[79\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7354 tdc0.o_result\[55\] a_4463_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7355 VGND a_11214_7093# _022_ VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X7356 VPWR a_16762_8207# clknet_4_11_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7357 VPWR tdc0.w_dly_sig_n\[37\] tdc0.w_dly_sig\[38\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7358 VPWR a_13919_7119# _001_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7359 VGND tdc0.w_dly_sig\[44\] tdc0.w_dly_sig\[46\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7360 a_11780_7637# _000_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.176 ps=1.68 w=0.42 l=0.15
X7361 a_2673_2767# a_1683_2767# a_2547_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7362 VGND a_17746_9407# a_17704_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7363 VPWR clknet_4_5_0_clk a_5087_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7364 a_8481_11471# tdc0.o_result\[59\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7365 a_17059_14735# a_16923_14709# a_16639_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7366 VPWR _042_ a_12237_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7367 VPWR a_4279_10651# a_4195_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7369 _060_ a_10055_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7370 a_11509_2045# a_10975_1679# a_11414_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7371 VPWR tdc0.w_dly_sig_n\[115\] tdc0.w_dly_sig\[116\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7372 VGND tdc0.w_dly_sig\[71\] tdc0.w_dly_sig\[73\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7373 a_4379_1135# a_3597_1141# a_4295_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7374 clknet_4_5_0_clk a_3348_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7375 tdc0.w_dly_sig_n\[6\] tdc0.w_dly_sig_n\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7376 a_13564_5865# a_13165_5493# a_13438_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7377 VPWR tdc0.w_dly_sig_n\[45\] tdc0.w_dly_sig_n\[47\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7378 VGND tdc0.w_dly_sig_n\[85\] tdc0.w_dly_sig_n\[87\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7379 VGND _059_ a_10607_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X7380 VGND a_16239_18267# a_16197_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7381 a_5618_5309# a_5345_4943# a_5533_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7382 a_11724_10927# _036_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7383 a_18142_10116# a_17935_10057# a_18318_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7384 VPWR clknet_4_0_0_clk a_5087_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7385 tdc0.w_dly_sig\[118\] tdc0.w_dly_sig\[116\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7386 VPWR _012_ a_9493_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7387 a_10321_10633# tdc0.o_result\[13\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X7388 VPWR a_8574_4676# a_8503_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X7389 a_11027_6005# _019_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X7390 a_13341_7779# _048_ a_13269_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7391 tdc0.w_dly_sig_n\[98\] tdc0.w_dly_sig\[98\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7392 tdc0.w_dly_sig_n\[100\] tdc0.w_dly_sig\[100\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7393 tdc0.w_dly_sig_n\[78\] tdc0.w_dly_sig_n\[76\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7395 a_9747_8181# _000_ a_10228_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0619 ps=0.715 w=0.42 l=0.15
X7396 a_17314_12559# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7397 VGND a_11642_5461# _019_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7398 VPWR clknet_4_8_0_clk a_13919_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7399 a_11333_15279# tdc0.o_result\[25\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X7400 VPWR a_9631_4221# a_9799_4123# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7401 clknet_4_13_0_clk a_14388_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7402 a_17378_1791# a_17210_2045# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7403 _013_ a_11159_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7406 a_14277_8867# _017_ a_14195_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X7407 a_16163_2045# a_15299_1679# a_15906_1791# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7408 a_11872_7093# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.312 ps=2.12 w=0.42 l=0.15
X7409 VPWR clknet_4_6_0_clk a_6651_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7410 a_11610_14468# a_11410_14313# a_11759_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7411 tdc0.w_dly_sig\[26\] tdc0.w_dly_sig\[24\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7412 a_18027_3529# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7413 VPWR tdc0.w_dly_sig\[104\] tdc0.w_dly_sig_n\[104\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7414 VGND tdc0.w_dly_sig\[43\] tdc0.w_dly_sig_n\[43\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7415 tdc0.w_dly_sig\[124\] tdc0.w_dly_sig\[122\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7416 a_18673_4777# a_18126_4521# a_18326_4676# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X7417 VGND tdc0.w_dly_sig_n\[36\] tdc0.w_dly_sig_n\[38\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7419 a_18054_8029# a_17739_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7420 a_1761_6575# tdc0.w_dly_sig\[77\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7421 VPWR a_4176_6005# clknet_4_0_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7422 VPWR tdc0.w_dly_sig\[24\] a_14717_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7423 tdc0.w_dly_sig\[22\] tdc0.w_dly_sig_n\[21\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7424 VGND tdc0.w_dly_sig\[91\] tdc0.w_dly_sig_n\[91\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7425 a_12258_17821# a_11943_17687# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7426 a_15162_5095# _085_ a_15465_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X7427 VPWR tdc0.w_dly_sig_n\[65\] tdc0.w_dly_sig_n\[67\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7428 a_1554_11989# a_1386_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7429 a_9807_18365# a_9025_17999# a_9723_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7430 VPWR a_7626_7637# a_7553_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7431 a_14899_9269# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7432 a_16819_5095# a_16915_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7433 tdc0.w_dly_sig\[82\] tdc0.w_dly_sig\[80\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7434 VPWR tdc0.w_dly_sig_n\[113\] tdc0.w_dly_sig_n\[115\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7435 VPWR a_7607_9839# a_7775_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
R31 tt_um_hpretl_tt06_tdc_20.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7436 tdc0.w_dly_sig\[61\] tdc0.w_dly_sig_n\[60\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7437 VPWR a_17187_17687# tdc0.o_result\[127\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7438 tdc0.w_dly_sig\[17\] tdc0.w_dly_sig_n\[16\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7439 a_18234_12292# a_18034_12137# a_18383_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7440 a_10091_3311# a_9227_3317# a_9834_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7441 VGND tdc0.w_dly_sig_n\[46\] tdc0.w_dly_sig_n\[48\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7442 clknet_4_1_0_clk a_3790_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7443 tdc0.w_dly_sig\[1\] tdc0.w_dly_sig_n\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7444 a_1386_12015# a_1113_12021# a_1301_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7445 tdc0.o_result\[29\] a_9799_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7446 tdc0.w_dly_sig_n\[27\] tdc0.w_dly_sig_n\[25\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7447 a_6998_2223# a_6559_2229# a_6913_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7448 a_17502_16733# a_17187_16599# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7449 VPWR clknet_4_1_0_clk a_4995_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7450 a_12118_9295# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7451 a_14431_15797# a_14722_16097# a_14673_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7452 a_2014_6549# a_1846_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7453 VGND a_11938_8253# _009_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7454 VPWR a_11058_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X7455 tdc0.w_dly_sig_n\[126\] tdc0.w_dly_sig\[126\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7456 VPWR a_9503_7663# a_9650_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.22 ps=1.44 w=1 l=0.15
X7457 a_1389_9845# a_1223_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7458 tdc0.w_dly_sig\[78\] tdc0.w_dly_sig_n\[77\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7459 a_14786_9071# _031_ a_14952_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7460 VPWR tdc0.w_dly_sig_n\[32\] tdc0.w_dly_sig_n\[34\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7461 _056_ a_10883_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7462 VGND a_6619_17973# a_6626_18273# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7463 VGND clknet_4_9_0_clk a_12999_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7464 tdc0.w_dly_sig\[61\] tdc0.w_dly_sig\[59\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7465 VGND a_9799_4123# a_9757_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7466 tdc0.w_dly_sig\[47\] tdc0.w_dly_sig\[45\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7467 a_7166_2197# a_6998_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7468 a_7691_3311# a_6909_3317# a_7607_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7470 tdc0.w_dly_sig\[24\] tdc0.w_dly_sig_n\[23\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7471 tdc0.w_dly_sig_n\[108\] tdc0.w_dly_sig_n\[106\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7472 VPWR a_10075_9563# a_9991_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7473 VGND tdc0.w_dly_sig_n\[81\] tdc0.w_dly_sig\[82\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7474 a_2685_12015# tdc0.o_result\[72\] a_2603_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7475 VGND tdc0.w_dly_sig\[86\] tdc0.w_dly_sig_n\[86\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 uio_in[4] VGND 0.182f
C1 uio_in[5] VGND 0.182f
C2 uio_in[6] VGND 0.182f
C3 uio_in[7] VGND 0.182f
C4 uio_in[0] VGND 0.182f
C5 uio_in[1] VGND 0.182f
C6 uio_in[2] VGND 0.182f
C7 uio_in[3] VGND 0.182f
C8 rst_n VGND 0.182f
C9 ui_in[1] VGND 0.182f
C10 ui_in[2] VGND 0.182f
C11 ui_in[7] VGND 0.182f
C12 ena VGND 0.182f
C13 uio_oe[6] VGND 1.05f
C14 uio_oe[3] VGND 1.57f
C15 ui_in[3] VGND 0.749f
C16 ui_in[5] VGND 0.877f
C17 ui_in[6] VGND 0.747f
C18 ui_in[4] VGND 0.768f
C19 uio_out[3] VGND 1.14f
C20 uio_out[7] VGND 0.927f
C21 uio_oe[7] VGND 0.955f
C22 uio_oe[5] VGND 1.22f
C23 uio_out[1] VGND 1.12f
C24 uo_out[4] VGND 2.5f
C25 uo_out[6] VGND 3.82f
C26 uo_out[1] VGND 4.38f
C27 uo_out[3] VGND 2.21f
C28 clk VGND 8.2f
C29 uo_out[5] VGND 4.29f
C30 ui_in[0] VGND 1.38f
C31 uo_out[7] VGND 3.89f
C32 uo_out[0] VGND 1.91f
C33 uo_out[2] VGND 2.74f
C34 uio_oe[0] VGND 1.22f
C35 uio_oe[2] VGND 1.04f
C36 uio_out[2] VGND 1.22f
C37 uio_out[4] VGND 1.21f
C38 uio_oe[4] VGND 1.12f
C39 uio_out[5] VGND 1.46f
C40 uio_out[6] VGND 1.39f
C41 uio_oe[1] VGND 1.56f
C42 uio_out[0] VGND 1.1f
C43 VPWR VGND 1.32p
C44 tt_um_hpretl_tt06_tdc_18.HI VGND 0.415f $ **FLOATING
C45 tt_um_hpretl_tt06_tdc_15.HI VGND 0.415f $ **FLOATING
C46 a_12999_591# VGND 0.698f $ **FLOATING
C47 a_12631_591# VGND 0.698f $ **FLOATING
C48 a_11711_591# VGND 0.698f $ **FLOATING
C49 a_10423_591# VGND 0.648f $ **FLOATING
C50 tt_um_hpretl_tt06_tdc_23.HI VGND 0.415f $ **FLOATING
C51 tt_um_hpretl_tt06_tdc_27.HI VGND 0.415f $ **FLOATING
C52 tt_um_hpretl_tt06_tdc_19.HI VGND 0.415f $ **FLOATING
C53 a_16849_1135# VGND 0.23f $ **FLOATING
C54 a_13813_1135# VGND 0.23f $ **FLOATING
C55 tdc0.w_dly_sig_n\[99\] VGND 2.26f $ **FLOATING
C56 a_8753_1135# VGND 0.23f $ **FLOATING
C57 a_7281_1135# VGND 0.23f $ **FLOATING
C58 a_3785_1135# VGND 0.23f $ **FLOATING
C59 a_2037_1135# VGND 0.23f $ **FLOATING
C60 a_17359_1135# VGND 0.609f $ **FLOATING
C61 a_17527_1109# VGND 0.817f $ **FLOATING
C62 a_16934_1135# VGND 0.626f $ **FLOATING
C63 a_17102_1109# VGND 0.581f $ **FLOATING
C64 a_16661_1141# VGND 1.43f $ **FLOATING
C65 a_16495_1141# VGND 1.81f $ **FLOATING
C66 tdc0.w_dly_sig\[102\] VGND 3.5f $ **FLOATING
C67 a_14323_1135# VGND 0.609f $ **FLOATING
C68 a_14491_1109# VGND 0.817f $ **FLOATING
C69 a_13898_1135# VGND 0.626f $ **FLOATING
C70 a_14066_1109# VGND 0.581f $ **FLOATING
C71 a_13625_1141# VGND 1.43f $ **FLOATING
C72 tdc0.w_dly_sig\[100\] VGND 2.97f $ **FLOATING
C73 a_13459_1141# VGND 1.81f $ **FLOATING
C74 a_9263_1135# VGND 0.609f $ **FLOATING
C75 a_9431_1109# VGND 0.817f $ **FLOATING
C76 a_8838_1135# VGND 0.626f $ **FLOATING
C77 a_9006_1109# VGND 0.581f $ **FLOATING
C78 a_8565_1141# VGND 1.43f $ **FLOATING
C79 a_8399_1141# VGND 1.81f $ **FLOATING
C80 a_7791_1135# VGND 0.609f $ **FLOATING
C81 a_7959_1109# VGND 0.817f $ **FLOATING
C82 a_7366_1135# VGND 0.626f $ **FLOATING
C83 a_7534_1109# VGND 0.581f $ **FLOATING
C84 a_7093_1141# VGND 1.43f $ **FLOATING
C85 a_6927_1141# VGND 1.81f $ **FLOATING
C86 a_4295_1135# VGND 0.609f $ **FLOATING
C87 a_4463_1109# VGND 0.817f $ **FLOATING
C88 a_3870_1135# VGND 0.626f $ **FLOATING
C89 a_4038_1109# VGND 0.581f $ **FLOATING
C90 a_3597_1141# VGND 1.43f $ **FLOATING
C91 a_3431_1141# VGND 1.81f $ **FLOATING
C92 a_2547_1135# VGND 0.609f $ **FLOATING
C93 a_2715_1109# VGND 0.817f $ **FLOATING
C94 a_2122_1135# VGND 0.626f $ **FLOATING
C95 a_2290_1109# VGND 0.581f $ **FLOATING
C96 a_1849_1141# VGND 1.43f $ **FLOATING
C97 a_1683_1141# VGND 1.81f $ **FLOATING
C98 tt_um_hpretl_tt06_tdc_17.HI VGND 0.415f $ **FLOATING
C99 a_17125_1679# VGND 0.23f $ **FLOATING
C100 a_17635_2045# VGND 0.609f $ **FLOATING
C101 a_17803_1947# VGND 0.817f $ **FLOATING
C102 a_17210_2045# VGND 0.626f $ **FLOATING
C103 a_17378_1791# VGND 0.581f $ **FLOATING
C104 a_16937_1679# VGND 1.43f $ **FLOATING
C105 a_16771_1679# VGND 1.81f $ **FLOATING
C106 a_15653_1679# VGND 0.23f $ **FLOATING
C107 a_16163_2045# VGND 0.609f $ **FLOATING
C108 a_16331_1947# VGND 0.817f $ **FLOATING
C109 a_15738_2045# VGND 0.626f $ **FLOATING
C110 a_15906_1791# VGND 0.581f $ **FLOATING
C111 a_15465_1679# VGND 1.43f $ **FLOATING
C112 a_15299_1679# VGND 1.81f $ **FLOATING
C113 tdc0.w_dly_sig_n\[103\] VGND 2.51f $ **FLOATING
C114 a_11329_1679# VGND 0.23f $ **FLOATING
C115 tdc0.w_dly_sig_n\[101\] VGND 2.61f $ **FLOATING
C116 tdc0.w_dly_sig_n\[102\] VGND 2.39f $ **FLOATING
C117 tdc0.w_dly_sig_n\[100\] VGND 2.53f $ **FLOATING
C118 tdc0.w_dly_sig_n\[98\] VGND 2.67f $ **FLOATING
C119 a_11839_2045# VGND 0.609f $ **FLOATING
C120 a_12007_1947# VGND 0.817f $ **FLOATING
C121 a_11414_2045# VGND 0.626f $ **FLOATING
C122 a_11582_1791# VGND 0.581f $ **FLOATING
C123 a_11141_1679# VGND 1.43f $ **FLOATING
C124 tdc0.w_dly_sig\[98\] VGND 2.96f $ **FLOATING
C125 a_10975_1679# VGND 1.81f $ **FLOATING
C126 a_9397_1679# VGND 0.23f $ **FLOATING
C127 a_9907_2045# VGND 0.609f $ **FLOATING
C128 a_10075_1947# VGND 0.817f $ **FLOATING
C129 a_9482_2045# VGND 0.626f $ **FLOATING
C130 a_9650_1791# VGND 0.581f $ **FLOATING
C131 a_9209_1679# VGND 1.43f $ **FLOATING
C132 a_9043_1679# VGND 1.81f $ **FLOATING
C133 tdc0.w_dly_sig_n\[96\] VGND 2.81f $ **FLOATING
C134 a_5717_1679# VGND 0.23f $ **FLOATING
C135 tdc0.w_dly_sig_n\[94\] VGND 1.79f $ **FLOATING
C136 tdc0.w_dly_sig\[92\] VGND 2.7f $ **FLOATING
C137 a_6227_2045# VGND 0.609f $ **FLOATING
C138 a_6395_1947# VGND 0.817f $ **FLOATING
C139 a_5802_2045# VGND 0.626f $ **FLOATING
C140 a_5970_1791# VGND 0.581f $ **FLOATING
C141 a_5529_1679# VGND 1.43f $ **FLOATING
C142 a_5363_1679# VGND 1.81f $ **FLOATING
C143 a_4245_1679# VGND 0.23f $ **FLOATING
C144 a_4755_2045# VGND 0.609f $ **FLOATING
C145 a_4923_1947# VGND 0.817f $ **FLOATING
C146 a_4330_2045# VGND 0.626f $ **FLOATING
C147 a_4498_1791# VGND 0.581f $ **FLOATING
C148 a_4057_1679# VGND 1.43f $ **FLOATING
C149 a_3891_1679# VGND 1.81f $ **FLOATING
C150 tdc0.w_dly_sig\[83\] VGND 3.44f $ **FLOATING
C151 tt_um_hpretl_tt06_tdc_21.HI VGND 0.415f $ **FLOATING
C152 a_14273_2223# VGND 0.23f $ **FLOATING
C153 a_10137_2223# VGND 0.206f $ **FLOATING
C154 a_9493_2223# VGND 0.206f $ **FLOATING
C155 a_12801_2223# VGND 0.23f $ **FLOATING
C156 tdc0.w_dly_sig_n\[97\] VGND 2.63f $ **FLOATING
C157 tdc0.w_dly_sig_n\[95\] VGND 2.76f $ **FLOATING
C158 tdc0.w_dly_sig\[96\] VGND 3.67f $ **FLOATING
C159 a_6913_2223# VGND 0.23f $ **FLOATING
C160 tdc0.w_dly_sig_n\[89\] VGND 2.18f $ **FLOATING
C161 tdc0.w_dly_sig_n\[82\] VGND 2.06f $ **FLOATING
C162 tdc0.w_dly_sig\[105\] VGND 3.07f $ **FLOATING
C163 a_14783_2223# VGND 0.609f $ **FLOATING
C164 a_14951_2197# VGND 0.817f $ **FLOATING
C165 a_14358_2223# VGND 0.626f $ **FLOATING
C166 a_14526_2197# VGND 0.581f $ **FLOATING
C167 a_14085_2229# VGND 1.43f $ **FLOATING
C168 a_13919_2229# VGND 1.81f $ **FLOATING
C169 a_13311_2223# VGND 0.609f $ **FLOATING
C170 a_13479_2197# VGND 0.817f $ **FLOATING
C171 a_12886_2223# VGND 0.626f $ **FLOATING
C172 a_13054_2197# VGND 0.581f $ **FLOATING
C173 a_12613_2229# VGND 1.43f $ **FLOATING
C174 a_12447_2229# VGND 1.81f $ **FLOATING
C175 tdc0.w_dly_sig\[97\] VGND 4.26f $ **FLOATING
C176 a_10055_2223# VGND 0.804f $ **FLOATING
C177 tdc0.o_result\[87\] VGND 2.61f $ **FLOATING
C178 tdc0.o_result\[95\] VGND 0.966f $ **FLOATING
C179 a_9411_2223# VGND 0.804f $ **FLOATING
C180 tdc0.o_result\[85\] VGND 2.91f $ **FLOATING
C181 tdc0.o_result\[93\] VGND 1.19f $ **FLOATING
C182 tdc0.w_dly_sig\[94\] VGND 3.13f $ **FLOATING
C183 tdc0.w_dly_sig_n\[93\] VGND 2.39f $ **FLOATING
C184 a_7423_2223# VGND 0.609f $ **FLOATING
C185 a_7591_2197# VGND 0.817f $ **FLOATING
C186 a_6998_2223# VGND 0.626f $ **FLOATING
C187 a_7166_2197# VGND 0.581f $ **FLOATING
C188 a_6725_2229# VGND 1.43f $ **FLOATING
C189 a_6559_2229# VGND 1.81f $ **FLOATING
C190 tdc0.w_dly_sig_n\[90\] VGND 2.58f $ **FLOATING
C191 tdc0.w_dly_sig_n\[88\] VGND 2.36f $ **FLOATING
C192 tdc0.w_dly_sig_n\[87\] VGND 3.17f $ **FLOATING
C193 tdc0.w_dly_sig_n\[86\] VGND 2.59f $ **FLOATING
C194 tdc0.w_dly_sig\[86\] VGND 3.05f $ **FLOATING
C195 tdc0.w_dly_sig\[85\] VGND 3.25f $ **FLOATING
C196 tdc0.w_dly_sig_n\[85\] VGND 3.32f $ **FLOATING
C197 tdc0.w_dly_sig_n\[84\] VGND 2.38f $ **FLOATING
C198 a_18121_2767# VGND 0.23f $ **FLOATING
C199 tdc0.w_dly_sig_n\[104\] VGND 2.51f $ **FLOATING
C200 tdc0.w_dly_sig\[111\] VGND 3.09f $ **FLOATING
C201 a_17703_2767# VGND 0.581f $ **FLOATING
C202 a_17774_2741# VGND 0.626f $ **FLOATING
C203 a_17567_2741# VGND 1.81f $ **FLOATING
C204 a_17574_3041# VGND 1.43f $ **FLOATING
C205 a_17283_2741# VGND 0.609f $ **FLOATING
C206 a_17187_2919# VGND 0.817f $ **FLOATING
C207 tdc0.w_dly_sig\[104\] VGND 3.67f $ **FLOATING
C208 tdc0.w_dly_sig_n\[106\] VGND 2.67f $ **FLOATING
C209 tdc0.w_dly_sig_n\[105\] VGND 2.91f $ **FLOATING
C210 tdc0.w_dly_sig\[99\] VGND 2.88f $ **FLOATING
C211 a_11865_2767# VGND 0.23f $ **FLOATING
C212 tdc0.w_dly_sig_n\[91\] VGND 3.12f $ **FLOATING
C213 tdc0.w_dly_sig\[90\] VGND 3.6f $ **FLOATING
C214 tdc0.w_dly_sig_n\[83\] VGND 2.95f $ **FLOATING
C215 a_2037_2767# VGND 0.23f $ **FLOATING
C216 tdc0.w_dly_sig\[103\] VGND 4.2f $ **FLOATING
C217 a_11447_2767# VGND 0.581f $ **FLOATING
C218 a_11518_2741# VGND 0.626f $ **FLOATING
C219 a_11311_2741# VGND 1.81f $ **FLOATING
C220 a_11318_3041# VGND 1.43f $ **FLOATING
C221 a_11027_2741# VGND 0.609f $ **FLOATING
C222 a_10931_2919# VGND 0.817f $ **FLOATING
C223 tdc0.w_dly_sig_n\[92\] VGND 2.99f $ **FLOATING
C224 tdc0.w_dly_sig\[88\] VGND 3.56f $ **FLOATING
C225 a_2547_3133# VGND 0.609f $ **FLOATING
C226 a_2715_3035# VGND 0.817f $ **FLOATING
C227 a_2122_3133# VGND 0.626f $ **FLOATING
C228 a_2290_2879# VGND 0.581f $ **FLOATING
C229 a_1849_2767# VGND 1.43f $ **FLOATING
C230 a_1683_2767# VGND 1.81f $ **FLOATING
C231 tdc0.w_dly_sig\[82\] VGND 2.71f $ **FLOATING
C232 tdc0.w_dly_sig_n\[81\] VGND 2.9f $ **FLOATING
C233 a_18581_3689# VGND 0.23f $ **FLOATING
C234 a_13353_3311# VGND 0.23f $ **FLOATING
C235 a_9581_3311# VGND 0.23f $ **FLOATING
C236 a_7097_3311# VGND 0.23f $ **FLOATING
C237 a_3969_3311# VGND 0.23f $ **FLOATING
C238 a_2313_3311# VGND 0.23f $ **FLOATING
C239 a_18163_3689# VGND 0.581f $ **FLOATING
C240 a_18234_3588# VGND 0.626f $ **FLOATING
C241 a_18034_3433# VGND 1.43f $ **FLOATING
C242 a_18027_3529# VGND 1.81f $ **FLOATING
C243 a_17743_3543# VGND 0.609f $ **FLOATING
C244 a_17647_3543# VGND 0.817f $ **FLOATING
C245 tdc0.w_dly_sig_n\[108\] VGND 2.15f $ **FLOATING
C246 tdc0.w_dly_sig_n\[107\] VGND 2.31f $ **FLOATING
C247 a_13863_3311# VGND 0.609f $ **FLOATING
C248 a_14031_3285# VGND 0.817f $ **FLOATING
C249 a_13438_3311# VGND 0.626f $ **FLOATING
C250 a_13606_3285# VGND 0.581f $ **FLOATING
C251 a_13165_3317# VGND 1.43f $ **FLOATING
C252 tdc0.w_dly_sig\[101\] VGND 3.16f $ **FLOATING
C253 a_12999_3317# VGND 1.81f $ **FLOATING
C254 a_10091_3311# VGND 0.609f $ **FLOATING
C255 a_10259_3285# VGND 0.817f $ **FLOATING
C256 a_9666_3311# VGND 0.626f $ **FLOATING
C257 a_9834_3285# VGND 0.581f $ **FLOATING
C258 a_9393_3317# VGND 1.43f $ **FLOATING
C259 tdc0.w_dly_sig\[95\] VGND 5.22f $ **FLOATING
C260 a_9227_3317# VGND 1.81f $ **FLOATING
C261 a_7607_3311# VGND 0.609f $ **FLOATING
C262 a_7775_3285# VGND 0.817f $ **FLOATING
C263 a_7182_3311# VGND 0.626f $ **FLOATING
C264 a_7350_3285# VGND 0.581f $ **FLOATING
C265 a_6909_3317# VGND 1.43f $ **FLOATING
C266 tdc0.w_dly_sig\[91\] VGND 3f $ **FLOATING
C267 a_6743_3317# VGND 1.81f $ **FLOATING
C268 a_4479_3311# VGND 0.609f $ **FLOATING
C269 a_4647_3285# VGND 0.817f $ **FLOATING
C270 a_4054_3311# VGND 0.626f $ **FLOATING
C271 a_4222_3285# VGND 0.581f $ **FLOATING
C272 a_3781_3317# VGND 1.43f $ **FLOATING
C273 tdc0.w_dly_sig\[84\] VGND 3.85f $ **FLOATING
C274 a_3615_3317# VGND 1.81f $ **FLOATING
C275 a_2823_3311# VGND 0.609f $ **FLOATING
C276 a_2991_3285# VGND 0.817f $ **FLOATING
C277 a_2398_3311# VGND 0.626f $ **FLOATING
C278 a_2566_3285# VGND 0.581f $ **FLOATING
C279 a_2125_3317# VGND 1.43f $ **FLOATING
C280 tdc0.w_dly_sig\[81\] VGND 3.33f $ **FLOATING
C281 a_1959_3317# VGND 1.81f $ **FLOATING
C282 tdc0.w_dly_sig\[113\] VGND 3.9f $ **FLOATING
C283 tdc0.w_dly_sig_n\[111\] VGND 2.51f $ **FLOATING
C284 tdc0.w_dly_sig_n\[110\] VGND 2.49f $ **FLOATING
C285 tdc0.w_dly_sig_n\[112\] VGND 1.75f $ **FLOATING
C286 tdc0.w_dly_sig_n\[109\] VGND 2.4f $ **FLOATING
C287 a_14533_3855# VGND 0.23f $ **FLOATING
C288 a_11973_3855# VGND 0.23f $ **FLOATING
C289 tdc0.w_dly_sig\[107\] VGND 4.07f $ **FLOATING
C290 a_14115_3855# VGND 0.581f $ **FLOATING
C291 a_14186_3829# VGND 0.626f $ **FLOATING
C292 a_13979_3829# VGND 1.81f $ **FLOATING
C293 a_13986_4129# VGND 1.43f $ **FLOATING
C294 a_13695_3829# VGND 0.609f $ **FLOATING
C295 a_13599_4007# VGND 0.817f $ **FLOATING
C296 a_12483_4221# VGND 0.609f $ **FLOATING
C297 a_12651_4123# VGND 0.817f $ **FLOATING
C298 a_12058_4221# VGND 0.626f $ **FLOATING
C299 a_12226_3967# VGND 0.581f $ **FLOATING
C300 a_11785_3855# VGND 1.43f $ **FLOATING
C301 tdc0.w_dly_sig\[106\] VGND 5.93f $ **FLOATING
C302 a_11619_3855# VGND 1.81f $ **FLOATING
C303 a_9121_3855# VGND 0.23f $ **FLOATING
C304 a_9631_4221# VGND 0.609f $ **FLOATING
C305 a_9799_4123# VGND 0.817f $ **FLOATING
C306 a_9206_4221# VGND 0.626f $ **FLOATING
C307 a_9374_3967# VGND 0.581f $ **FLOATING
C308 a_8933_3855# VGND 1.43f $ **FLOATING
C309 tdc0.w_dly_sig\[110\] VGND 5.02f $ **FLOATING
C310 a_8767_3855# VGND 1.81f $ **FLOATING
C311 a_7189_3855# VGND 0.23f $ **FLOATING
C312 a_7699_4221# VGND 0.609f $ **FLOATING
C313 a_7867_4123# VGND 0.817f $ **FLOATING
C314 a_7274_4221# VGND 0.626f $ **FLOATING
C315 a_7442_3967# VGND 0.581f $ **FLOATING
C316 a_7001_3855# VGND 1.43f $ **FLOATING
C317 tdc0.w_dly_sig\[93\] VGND 3.4f $ **FLOATING
C318 a_6835_3855# VGND 1.81f $ **FLOATING
C319 a_5441_3855# VGND 0.23f $ **FLOATING
C320 a_5951_4221# VGND 0.609f $ **FLOATING
C321 a_6119_4123# VGND 0.817f $ **FLOATING
C322 a_5526_4221# VGND 0.626f $ **FLOATING
C323 a_5694_3967# VGND 0.581f $ **FLOATING
C324 a_5253_3855# VGND 1.43f $ **FLOATING
C325 tdc0.w_dly_sig\[87\] VGND 4.12f $ **FLOATING
C326 a_5087_3855# VGND 1.81f $ **FLOATING
C327 tdc0.w_dly_sig_n\[80\] VGND 3.61f $ **FLOATING
C328 a_18673_4777# VGND 0.23f $ **FLOATING
C329 a_12345_4399# VGND 0.206f $ **FLOATING
C330 a_11609_4399# VGND 0.206f $ **FLOATING
C331 a_10977_4399# VGND 0.253f $ **FLOATING
C332 a_14917_4399# VGND 0.23f $ **FLOATING
C333 a_10393_4777# VGND 0.23f $ **FLOATING
C334 a_8921_4777# VGND 0.23f $ **FLOATING
C335 a_6453_4399# VGND 0.23f $ **FLOATING
C336 a_4245_4399# VGND 0.23f $ **FLOATING
C337 a_1945_4399# VGND 0.23f $ **FLOATING
C338 tdc0.w_dly_sig_n\[79\] VGND 2.5f $ **FLOATING
C339 a_18255_4777# VGND 0.581f $ **FLOATING
C340 a_18326_4676# VGND 0.626f $ **FLOATING
C341 a_18126_4521# VGND 1.43f $ **FLOATING
C342 a_18119_4617# VGND 1.81f $ **FLOATING
C343 a_17835_4631# VGND 0.609f $ **FLOATING
C344 a_17739_4631# VGND 0.817f $ **FLOATING
C345 a_15427_4399# VGND 0.609f $ **FLOATING
C346 a_15595_4373# VGND 0.817f $ **FLOATING
C347 a_15002_4399# VGND 0.626f $ **FLOATING
C348 a_15170_4373# VGND 0.581f $ **FLOATING
C349 a_14729_4405# VGND 1.43f $ **FLOATING
C350 tdc0.w_dly_sig\[108\] VGND 3.11f $ **FLOATING
C351 a_14563_4405# VGND 1.81f $ **FLOATING
C352 tdc0.o_result\[97\] VGND 1.99f $ **FLOATING
C353 a_12199_4631# VGND 0.804f $ **FLOATING
C354 a_11527_4399# VGND 0.804f $ **FLOATING
C355 tdc0.o_result\[102\] VGND 1.69f $ **FLOATING
C356 tdc0.o_result\[78\] VGND 4.39f $ **FLOATING
C357 a_11146_4719# VGND 0.55f $ **FLOATING
C358 tdc0.o_result\[86\] VGND 3.01f $ **FLOATING
C359 tdc0.w_dly_sig\[112\] VGND 5.79f $ **FLOATING
C360 a_9975_4777# VGND 0.581f $ **FLOATING
C361 a_10046_4676# VGND 0.626f $ **FLOATING
C362 a_9846_4521# VGND 1.43f $ **FLOATING
C363 a_9839_4617# VGND 1.81f $ **FLOATING
C364 a_9555_4631# VGND 0.609f $ **FLOATING
C365 a_9459_4631# VGND 0.817f $ **FLOATING
C366 tdc0.w_dly_sig\[109\] VGND 6.67f $ **FLOATING
C367 a_8503_4777# VGND 0.581f $ **FLOATING
C368 a_8574_4676# VGND 0.626f $ **FLOATING
C369 a_8374_4521# VGND 1.43f $ **FLOATING
C370 a_8367_4617# VGND 1.81f $ **FLOATING
C371 a_8083_4631# VGND 0.609f $ **FLOATING
C372 a_7987_4631# VGND 0.817f $ **FLOATING
C373 a_6963_4399# VGND 0.609f $ **FLOATING
C374 a_7131_4373# VGND 0.817f $ **FLOATING
C375 a_6538_4399# VGND 0.626f $ **FLOATING
C376 a_6706_4373# VGND 0.581f $ **FLOATING
C377 a_6265_4405# VGND 1.43f $ **FLOATING
C378 tdc0.w_dly_sig\[89\] VGND 3.53f $ **FLOATING
C379 a_6099_4405# VGND 1.81f $ **FLOATING
C380 a_4755_4399# VGND 0.609f $ **FLOATING
C381 a_4923_4373# VGND 0.817f $ **FLOATING
C382 a_4330_4399# VGND 0.626f $ **FLOATING
C383 a_4498_4373# VGND 0.581f $ **FLOATING
C384 a_4057_4405# VGND 1.43f $ **FLOATING
C385 a_3891_4405# VGND 1.81f $ **FLOATING
C386 a_2455_4399# VGND 0.609f $ **FLOATING
C387 a_2623_4373# VGND 0.817f $ **FLOATING
C388 a_2030_4399# VGND 0.626f $ **FLOATING
C389 a_2198_4373# VGND 0.581f $ **FLOATING
C390 a_1757_4405# VGND 1.43f $ **FLOATING
C391 a_1591_4405# VGND 1.81f $ **FLOATING
C392 a_17753_4943# VGND 0.23f $ **FLOATING
C393 tdc0.o_result\[113\] VGND 2.49f $ **FLOATING
C394 a_14375_5193# VGND 0.253f $ **FLOATING
C395 a_13823_5193# VGND 0.253f $ **FLOATING
C396 clknet_4_8_0_clk VGND 8.49f $ **FLOATING
C397 a_10505_5193# VGND 0.206f $ **FLOATING
C398 a_9677_5193# VGND 0.206f $ **FLOATING
C399 clknet_4_2_0_clk VGND 10f $ **FLOATING
C400 a_5533_4943# VGND 0.23f $ **FLOATING
C401 a_17335_4943# VGND 0.581f $ **FLOATING
C402 a_17406_4917# VGND 0.626f $ **FLOATING
C403 a_17199_4917# VGND 1.81f $ **FLOATING
C404 a_17206_5217# VGND 1.43f $ **FLOATING
C405 a_16915_4917# VGND 0.609f $ **FLOATING
C406 a_16819_5095# VGND 0.817f $ **FLOATING
C407 a_15162_5095# VGND 0.702f $ **FLOATING
C408 tdc0.o_result\[100\] VGND 1.25f $ **FLOATING
C409 a_14157_4917# VGND 0.55f $ **FLOATING
C410 tdc0.o_result\[105\] VGND 1.54f $ **FLOATING
C411 a_13605_4917# VGND 0.55f $ **FLOATING
C412 a_12548_4917# VGND 1.98f $ **FLOATING
C413 a_11159_4943# VGND 1.31f $ **FLOATING
C414 a_11154_5095# VGND 0.905f $ **FLOATING
C415 a_10423_5193# VGND 0.804f $ **FLOATING
C416 tdc0.o_result\[111\] VGND 1.2f $ **FLOATING
C417 tdc0.o_result\[109\] VGND 1.11f $ **FLOATING
C418 a_9531_5095# VGND 0.804f $ **FLOATING
C419 a_8500_4917# VGND 1.98f $ **FLOATING
C420 a_6043_5309# VGND 0.609f $ **FLOATING
C421 a_6211_5211# VGND 0.817f $ **FLOATING
C422 a_5618_5309# VGND 0.626f $ **FLOATING
C423 a_5786_5055# VGND 0.581f $ **FLOATING
C424 a_5345_4943# VGND 1.43f $ **FLOATING
C425 a_5179_4943# VGND 1.81f $ **FLOATING
C426 tdc0.o_result\[69\] VGND 2.65f $ **FLOATING
C427 a_4061_4943# VGND 0.23f $ **FLOATING
C428 a_4571_5309# VGND 0.609f $ **FLOATING
C429 a_4739_5211# VGND 0.817f $ **FLOATING
C430 a_4146_5309# VGND 0.626f $ **FLOATING
C431 a_4314_5055# VGND 0.581f $ **FLOATING
C432 a_3873_4943# VGND 1.43f $ **FLOATING
C433 a_3707_4943# VGND 1.81f $ **FLOATING
C434 a_2037_4943# VGND 0.23f $ **FLOATING
C435 a_2547_5309# VGND 0.609f $ **FLOATING
C436 a_2715_5211# VGND 0.817f $ **FLOATING
C437 a_2122_5309# VGND 0.626f $ **FLOATING
C438 a_2290_5055# VGND 0.581f $ **FLOATING
C439 a_1849_4943# VGND 1.43f $ **FLOATING
C440 a_1683_4943# VGND 1.81f $ **FLOATING
C441 tdc0.w_dly_sig\[79\] VGND 3.22f $ **FLOATING
C442 a_16951_5487# VGND 0.253f $ **FLOATING
C443 a_16399_5487# VGND 0.253f $ **FLOATING
C444 a_15381_5487# VGND 0.206f $ **FLOATING
C445 a_14645_5487# VGND 0.206f $ **FLOATING
C446 _084_ VGND 1.11f $ **FLOATING
C447 _085_ VGND 1.01f $ **FLOATING
C448 a_13353_5487# VGND 0.23f $ **FLOATING
C449 a_11422_5487# VGND 0.36f $ **FLOATING
C450 a_11225_5487# VGND 0.247f $ **FLOATING
C451 a_10975_5487# VGND 0.393f $ **FLOATING
C452 a_9217_5487# VGND 0.206f $ **FLOATING
C453 a_8573_5487# VGND 0.206f $ **FLOATING
C454 _082_ VGND 3.37f $ **FLOATING
C455 a_5905_5487# VGND 0.206f $ **FLOATING
C456 a_7373_5487# VGND 0.23f $ **FLOATING
C457 tdc0.o_result\[71\] VGND 3.85f $ **FLOATING
C458 a_3509_5487# VGND 0.23f $ **FLOATING
C459 tdc0.w_dly_sig\[80\] VGND 3.51f $ **FLOATING
C460 tdc0.w_dly_sig_n\[78\] VGND 2.81f $ **FLOATING
C461 tdc0.w_dly_sig_n\[113\] VGND 2.98f $ **FLOATING
C462 tdc0.w_dly_sig_n\[114\] VGND 2.88f $ **FLOATING
C463 tdc0.w_dly_sig\[114\] VGND 2.89f $ **FLOATING
C464 tdc0.o_result\[112\] VGND 1.8f $ **FLOATING
C465 a_16733_5461# VGND 0.55f $ **FLOATING
C466 tdc0.o_result\[114\] VGND 1.7f $ **FLOATING
C467 a_16181_5461# VGND 0.55f $ **FLOATING
C468 tdc0.o_result\[98\] VGND 2.74f $ **FLOATING
C469 tdc0.o_result\[10\] VGND 1.1f $ **FLOATING
C470 a_15235_5719# VGND 0.804f $ **FLOATING
C471 a_14563_5487# VGND 0.804f $ **FLOATING
C472 tdc0.o_result\[96\] VGND 2.54f $ **FLOATING
C473 a_13863_5487# VGND 0.609f $ **FLOATING
C474 a_14031_5461# VGND 0.817f $ **FLOATING
C475 a_13438_5487# VGND 0.626f $ **FLOATING
C476 a_13606_5461# VGND 0.581f $ **FLOATING
C477 a_13165_5493# VGND 1.43f $ **FLOATING
C478 a_12999_5493# VGND 1.81f $ **FLOATING
C479 a_12171_5487# VGND 0.698f $ **FLOATING
C480 a_11642_5461# VGND 0.649f $ **FLOATING
C481 a_9135_5487# VGND 0.804f $ **FLOATING
C482 tdc0.o_result\[34\] VGND 1.28f $ **FLOATING
C483 tdc0.o_result\[90\] VGND 1.86f $ **FLOATING
C484 a_8491_5487# VGND 0.804f $ **FLOATING
C485 tdc0.o_result\[88\] VGND 1.44f $ **FLOATING
C486 a_7883_5487# VGND 0.609f $ **FLOATING
C487 a_8051_5461# VGND 0.817f $ **FLOATING
C488 a_7458_5487# VGND 0.626f $ **FLOATING
C489 a_7626_5461# VGND 0.581f $ **FLOATING
C490 a_7185_5493# VGND 1.43f $ **FLOATING
C491 a_7019_5493# VGND 1.81f $ **FLOATING
C492 a_5823_5487# VGND 0.804f $ **FLOATING
C493 tdc0.o_result\[83\] VGND 2.06f $ **FLOATING
C494 tdc0.o_result\[67\] VGND 1.24f $ **FLOATING
C495 a_4019_5487# VGND 0.609f $ **FLOATING
C496 a_4187_5461# VGND 0.817f $ **FLOATING
C497 a_3594_5487# VGND 0.626f $ **FLOATING
C498 a_3762_5461# VGND 0.581f $ **FLOATING
C499 a_3321_5493# VGND 1.43f $ **FLOATING
C500 a_3155_5493# VGND 1.81f $ **FLOATING
C501 a_16301_6281# VGND 0.206f $ **FLOATING
C502 _062_ VGND 4.25f $ **FLOATING
C503 _064_ VGND 1.23f $ **FLOATING
C504 _065_ VGND 0.992f $ **FLOATING
C505 _063_ VGND 0.835f $ **FLOATING
C506 a_14093_6281# VGND 0.206f $ **FLOATING
C507 _083_ VGND 1.71f $ **FLOATING
C508 a_8941_6281# VGND 0.206f $ **FLOATING
C509 tdc0.o_result\[32\] VGND 1.03f $ **FLOATING
C510 a_7189_6031# VGND 0.23f $ **FLOATING
C511 tdc0.w_dly_sig\[115\] VGND 3.41f $ **FLOATING
C512 tdc0.w_dly_sig_n\[115\] VGND 1.99f $ **FLOATING
C513 tdc0.o_result\[104\] VGND 2.25f $ **FLOATING
C514 a_16155_6183# VGND 0.804f $ **FLOATING
C515 a_15575_6281# VGND 0.702f $ **FLOATING
C516 a_14664_6005# VGND 1.98f $ **FLOATING
C517 tdc0.o_result\[106\] VGND 2f $ **FLOATING
C518 a_13947_6183# VGND 0.804f $ **FLOATING
C519 a_12148_6005# VGND 0.619f $ **FLOATING
C520 a_11343_6031# VGND 0.897f $ **FLOATING
C521 a_11490_6005# VGND 1.24f $ **FLOATING
C522 a_11027_6005# VGND 0.698f $ **FLOATING
C523 a_8859_6281# VGND 0.804f $ **FLOATING
C524 _019_ VGND 4.57f $ **FLOATING
C525 tdc0.o_result\[68\] VGND 2.13f $ **FLOATING
C526 tdc0.o_result\[108\] VGND 1.73f $ **FLOATING
C527 a_7699_6397# VGND 0.609f $ **FLOATING
C528 a_7867_6299# VGND 0.817f $ **FLOATING
C529 a_7274_6397# VGND 0.626f $ **FLOATING
C530 a_7442_6143# VGND 0.581f $ **FLOATING
C531 a_7001_6031# VGND 1.43f $ **FLOATING
C532 a_6835_6031# VGND 1.81f $ **FLOATING
C533 a_5721_6281# VGND 0.206f $ **FLOATING
C534 clknet_4_0_0_clk VGND 14.5f $ **FLOATING
C535 tdc0.w_dly_sig_n\[77\] VGND 2.39f $ **FLOATING
C536 a_5639_6281# VGND 0.804f $ **FLOATING
C537 tdc0.o_result\[82\] VGND 3.81f $ **FLOATING
C538 a_4176_6005# VGND 1.98f $ **FLOATING
C539 tdc0.w_dly_sig\[70\] VGND 3.58f $ **FLOATING
C540 a_18489_6953# VGND 0.23f $ **FLOATING
C541 clknet_4_10_0_clk VGND 10.8f $ **FLOATING
C542 tdc0.o_result\[8\] VGND 1.26f $ **FLOATING
C543 a_13997_6575# VGND 0.23f $ **FLOATING
C544 a_10226_6575# VGND 0.36f $ **FLOATING
C545 a_10029_6575# VGND 0.247f $ **FLOATING
C546 a_9779_6575# VGND 0.393f $ **FLOATING
C547 a_9125_6575# VGND 0.206f $ **FLOATING
C548 a_8481_6575# VGND 0.206f $ **FLOATING
C549 tdc0.o_result\[58\] VGND 3.97f $ **FLOATING
C550 a_6269_6575# VGND 0.23f $ **FLOATING
C551 tdc0.o_result\[66\] VGND 0.847f $ **FLOATING
C552 a_4521_6575# VGND 0.23f $ **FLOATING
C553 a_1761_6575# VGND 0.23f $ **FLOATING
C554 tdc0.w_dly_sig_n\[76\] VGND 2.71f $ **FLOATING
C555 a_18071_6953# VGND 0.581f $ **FLOATING
C556 a_18142_6852# VGND 0.626f $ **FLOATING
C557 a_17942_6697# VGND 1.43f $ **FLOATING
C558 a_17935_6793# VGND 1.81f $ **FLOATING
C559 a_17651_6807# VGND 0.609f $ **FLOATING
C560 a_17555_6807# VGND 0.817f $ **FLOATING
C561 a_16412_6549# VGND 1.98f $ **FLOATING
C562 a_14507_6575# VGND 0.609f $ **FLOATING
C563 a_14675_6549# VGND 0.817f $ **FLOATING
C564 a_14082_6575# VGND 0.626f $ **FLOATING
C565 a_14250_6549# VGND 0.581f $ **FLOATING
C566 a_13809_6581# VGND 1.43f $ **FLOATING
C567 a_13643_6581# VGND 1.81f $ **FLOATING
C568 a_13183_6583# VGND 0.648f $ **FLOATING
C569 a_12792_6549# VGND 0.619f $ **FLOATING
C570 a_11987_6575# VGND 0.897f $ **FLOATING
C571 a_12134_6549# VGND 1.24f $ **FLOATING
C572 a_11386_6652# VGND 0.658f $ **FLOATING
C573 a_10446_6549# VGND 0.649f $ **FLOATING
C574 a_9043_6575# VGND 0.804f $ **FLOATING
C575 tdc0.o_result\[116\] VGND 4.42f $ **FLOATING
C576 tdc0.o_result\[76\] VGND 3.86f $ **FLOATING
C577 a_8399_6575# VGND 0.804f $ **FLOATING
C578 tdc0.o_result\[91\] VGND 2.74f $ **FLOATING
C579 a_6779_6575# VGND 0.609f $ **FLOATING
C580 a_6947_6549# VGND 0.817f $ **FLOATING
C581 a_6354_6575# VGND 0.626f $ **FLOATING
C582 a_6522_6549# VGND 0.581f $ **FLOATING
C583 a_6081_6581# VGND 1.43f $ **FLOATING
C584 a_5915_6581# VGND 1.81f $ **FLOATING
C585 a_5031_6575# VGND 0.609f $ **FLOATING
C586 a_5199_6549# VGND 0.817f $ **FLOATING
C587 a_4606_6575# VGND 0.626f $ **FLOATING
C588 a_4774_6549# VGND 0.581f $ **FLOATING
C589 a_4333_6581# VGND 1.43f $ **FLOATING
C590 a_4167_6581# VGND 1.81f $ **FLOATING
C591 tdc0.w_dly_sig_n\[68\] VGND 1.97f $ **FLOATING
C592 a_2271_6575# VGND 0.609f $ **FLOATING
C593 a_2439_6549# VGND 0.817f $ **FLOATING
C594 a_1846_6575# VGND 0.626f $ **FLOATING
C595 a_2014_6549# VGND 0.581f $ **FLOATING
C596 a_1573_6581# VGND 1.43f $ **FLOATING
C597 tdc0.w_dly_sig\[77\] VGND 3.46f $ **FLOATING
C598 a_1407_6581# VGND 1.81f $ **FLOATING
C599 tdc0.w_dly_sig\[117\] VGND 2.92f $ **FLOATING
C600 tdc0.w_dly_sig_n\[116\] VGND 2.36f $ **FLOATING
C601 a_17385_7119# VGND 0.23f $ **FLOATING
C602 a_15853_7369# VGND 0.253f $ **FLOATING
C603 a_16967_7119# VGND 0.581f $ **FLOATING
C604 a_17038_7093# VGND 0.626f $ **FLOATING
C605 a_16831_7093# VGND 1.81f $ **FLOATING
C606 a_16838_7393# VGND 1.43f $ **FLOATING
C607 a_16547_7093# VGND 0.609f $ **FLOATING
C608 a_16451_7271# VGND 0.817f $ **FLOATING
C609 a_16022_7119# VGND 0.55f $ **FLOATING
C610 net8 VGND 6.59f $ **FLOATING
C611 tdc0.o_result\[115\] VGND 0.798f $ **FLOATING
C612 a_14287_7119# VGND 0.648f $ **FLOATING
C613 a_13919_7119# VGND 0.648f $ **FLOATING
C614 a_10595_7369# VGND 0.35f $ **FLOATING
C615 a_10401_7369# VGND 0.249f $ **FLOATING
C616 a_10147_7369# VGND 0.381f $ **FLOATING
C617 a_6549_7369# VGND 0.206f $ **FLOATING
C618 a_5349_7119# VGND 0.23f $ **FLOATING
C619 a_13603_7093# VGND 0.698f $ **FLOATING
C620 a_12518_7119# VGND 1.24f $ **FLOATING
C621 a_12642_7271# VGND 0.897f $ **FLOATING
C622 a_12263_7119# VGND 0.619f $ **FLOATING
C623 a_11872_7093# VGND 0.619f $ **FLOATING
C624 a_11067_7119# VGND 0.897f $ **FLOATING
C625 a_11214_7093# VGND 1.24f $ **FLOATING
C626 a_9485_7485# VGND 0.85f $ **FLOATING
C627 a_9319_7485# VGND 0.604f $ **FLOATING
C628 a_8995_7093# VGND 0.604f $ **FLOATING
C629 a_8543_7093# VGND 0.85f $ **FLOATING
C630 a_7286_7119# VGND 1.98f $ **FLOATING
C631 a_6467_7369# VGND 0.804f $ **FLOATING
C632 tdc0.o_result\[80\] VGND 3.65f $ **FLOATING
C633 tdc0.o_result\[64\] VGND 0.63f $ **FLOATING
C634 a_5859_7485# VGND 0.609f $ **FLOATING
C635 a_6027_7387# VGND 0.817f $ **FLOATING
C636 a_5434_7485# VGND 0.626f $ **FLOATING
C637 a_5602_7231# VGND 0.581f $ **FLOATING
C638 a_5161_7119# VGND 1.43f $ **FLOATING
C639 a_4995_7119# VGND 1.81f $ **FLOATING
C640 a_3790_7119# VGND 1.98f $ **FLOATING
C641 tdc0.w_dly_sig\[69\] VGND 4.37f $ **FLOATING
C642 a_18673_8041# VGND 0.23f $ **FLOATING
C643 a_15565_7663# VGND 0.206f $ **FLOATING
C644 a_14829_7663# VGND 0.206f $ **FLOATING
C645 a_18255_8041# VGND 0.581f $ **FLOATING
C646 a_18326_7940# VGND 0.626f $ **FLOATING
C647 a_18126_7785# VGND 1.43f $ **FLOATING
C648 a_18119_7881# VGND 1.81f $ **FLOATING
C649 a_17835_7895# VGND 0.609f $ **FLOATING
C650 a_17739_7895# VGND 0.817f $ **FLOATING
C651 tdc0.w_dly_sig\[116\] VGND 3.11f $ **FLOATING
C652 a_16127_7779# VGND 0.702f $ **FLOATING
C653 _092_ VGND 5.49f $ **FLOATING
C654 _094_ VGND 0.832f $ **FLOATING
C655 _095_ VGND 1.11f $ **FLOATING
C656 tdc0.o_result\[118\] VGND 1.33f $ **FLOATING
C657 tdc0.o_result\[110\] VGND 3.35f $ **FLOATING
C658 a_15419_7895# VGND 0.804f $ **FLOATING
C659 a_14747_7663# VGND 0.804f $ **FLOATING
C660 tdc0.o_result\[99\] VGND 3.53f $ **FLOATING
C661 a_14195_7663# VGND 0.698f $ **FLOATING
C662 a_13690_7895# VGND 0.702f $ **FLOATING
C663 a_13091_7779# VGND 0.702f $ **FLOATING
C664 _050_ VGND 2.45f $ **FLOATING
C665 tdc0.o_result\[35\] VGND 1.12f $ **FLOATING
C666 a_7373_7663# VGND 0.23f $ **FLOATING
C667 tdc0.w_dly_sig\[67\] VGND 3.92f $ **FLOATING
C668 tdc0.w_dly_sig_n\[66\] VGND 2.61f $ **FLOATING
C669 tdc0.w_dly_sig\[68\] VGND 4.08f $ **FLOATING
C670 tdc0.w_dly_sig_n\[71\] VGND 2.49f $ **FLOATING
C671 net5 VGND 8.66f $ **FLOATING
C672 a_12649_7814# VGND 0.696f $ **FLOATING
C673 a_12171_7663# VGND 0.788f $ **FLOATING
C674 a_12318_7637# VGND 0.795f $ **FLOATING
C675 a_11780_7637# VGND 0.619f $ **FLOATING
C676 a_10975_7663# VGND 0.897f $ **FLOATING
C677 net4 VGND 9.24f $ **FLOATING
C678 a_11122_7637# VGND 1.24f $ **FLOATING
C679 a_10515_7671# VGND 0.648f $ **FLOATING
C680 a_9503_7663# VGND 0.905f $ **FLOATING
C681 a_9650_7637# VGND 1.31f $ **FLOATING
C682 _023_ VGND 3.6f $ **FLOATING
C683 a_8819_7637# VGND 0.698f $ **FLOATING
C684 a_7883_7663# VGND 0.609f $ **FLOATING
C685 a_8051_7637# VGND 0.817f $ **FLOATING
C686 a_7458_7663# VGND 0.626f $ **FLOATING
C687 a_7626_7637# VGND 0.581f $ **FLOATING
C688 a_7185_7669# VGND 1.43f $ **FLOATING
C689 a_7019_7669# VGND 1.81f $ **FLOATING
C690 tdc0.w_dly_sig_n\[67\] VGND 2.76f $ **FLOATING
C691 tdc0.w_dly_sig_n\[69\] VGND 2.49f $ **FLOATING
C692 tdc0.w_dly_sig_n\[70\] VGND 2.88f $ **FLOATING
C693 tdc0.w_dly_sig\[72\] VGND 4.59f $ **FLOATING
C694 tdc0.w_dly_sig_n\[73\] VGND 2.01f $ **FLOATING
C695 a_17865_8457# VGND 0.206f $ **FLOATING
C696 _093_ VGND 1.12f $ **FLOATING
C697 a_16117_8457# VGND 0.206f $ **FLOATING
C698 tdc0.o_result\[11\] VGND 0.831f $ **FLOATING
C699 a_13905_8207# VGND 0.23f $ **FLOATING
C700 tdc0.o_result\[103\] VGND 3.2f $ **FLOATING
C701 a_17719_8359# VGND 0.804f $ **FLOATING
C702 a_16762_8207# VGND 1.98f $ **FLOATING
C703 a_16035_8457# VGND 0.804f $ **FLOATING
C704 _020_ VGND 9.83f $ **FLOATING
C705 tdc0.o_result\[107\] VGND 2.08f $ **FLOATING
C706 a_14415_8573# VGND 0.609f $ **FLOATING
C707 a_14583_8475# VGND 0.817f $ **FLOATING
C708 a_13990_8573# VGND 0.626f $ **FLOATING
C709 a_14158_8319# VGND 0.581f $ **FLOATING
C710 a_13717_8207# VGND 1.43f $ **FLOATING
C711 a_13551_8207# VGND 1.81f $ **FLOATING
C712 clknet_4_9_0_clk VGND 6.71f $ **FLOATING
C713 a_13353_8207# VGND 0.227f $ **FLOATING
C714 net3 VGND 8.75f $ **FLOATING
C715 a_11333_8457# VGND 0.206f $ **FLOATING
C716 _021_ VGND 1.49f $ **FLOATING
C717 _027_ VGND 1.56f $ **FLOATING
C718 _030_ VGND 0.682f $ **FLOATING
C719 a_8481_8457# VGND 0.206f $ **FLOATING
C720 a_6361_8207# VGND 0.23f $ **FLOATING
C721 a_13176_8207# VGND 0.498f $ **FLOATING
C722 a_13070_8207# VGND 0.578f $ **FLOATING
C723 a_12893_8207# VGND 0.5f $ **FLOATING
C724 a_12574_8207# VGND 0.535f $ **FLOATING
C725 _006_ VGND 3.41f $ **FLOATING
C726 a_11938_8253# VGND 0.658f $ **FLOATING
C727 net2 VGND 8.66f $ **FLOATING
C728 a_11251_8457# VGND 0.804f $ **FLOATING
C729 _004_ VGND 2.08f $ **FLOATING
C730 a_10759_8181# VGND 1.2f $ **FLOATING
C731 _000_ VGND 9.47f $ **FLOATING
C732 _001_ VGND 10.5f $ **FLOATING
C733 _002_ VGND 9.59f $ **FLOATING
C734 _003_ VGND 11f $ **FLOATING
C735 a_9747_8181# VGND 0.887f $ **FLOATING
C736 a_9043_8457# VGND 0.702f $ **FLOATING
C737 a_8399_8457# VGND 0.804f $ **FLOATING
C738 tdc0.o_result\[92\] VGND 2.6f $ **FLOATING
C739 a_6871_8573# VGND 0.609f $ **FLOATING
C740 a_7039_8475# VGND 0.817f $ **FLOATING
C741 a_6446_8573# VGND 0.626f $ **FLOATING
C742 a_6614_8319# VGND 0.581f $ **FLOATING
C743 a_6173_8207# VGND 1.43f $ **FLOATING
C744 a_6007_8207# VGND 1.81f $ **FLOATING
C745 tdc0.w_dly_sig_n\[74\] VGND 2.77f $ **FLOATING
C746 tdc0.w_dly_sig\[65\] VGND 2.82f $ **FLOATING
C747 tdc0.w_dly_sig_n\[65\] VGND 1.93f $ **FLOATING
C748 tdc0.w_dly_sig_n\[72\] VGND 2.61f $ **FLOATING
C749 tdc0.w_dly_sig_n\[75\] VGND 3.09f $ **FLOATING
C750 a_18325_8751# VGND 0.206f $ **FLOATING
C751 a_15220_8751# VGND 0.14f $ **FLOATING
C752 a_14868_8751# VGND 0.171f $ **FLOATING
C753 a_13541_8751# VGND 0.206f $ **FLOATING
C754 a_12644_8751# VGND 0.14f $ **FLOATING
C755 a_12292_8751# VGND 0.171f $ **FLOATING
C756 a_11057_8751# VGND 0.206f $ **FLOATING
C757 a_10321_8751# VGND 0.206f $ **FLOATING
C758 a_9125_8751# VGND 0.206f $ **FLOATING
C759 a_17033_8751# VGND 0.23f $ **FLOATING
C760 a_14786_9071# VGND 0.482f $ **FLOATING
C761 tdc0.w_dly_sig_n\[118\] VGND 2.65f $ **FLOATING
C762 tdc0.o_result\[117\] VGND 0.867f $ **FLOATING
C763 _025_ VGND 11.4f $ **FLOATING
C764 tdc0.o_result\[101\] VGND 3.82f $ **FLOATING
C765 _015_ VGND 9.04f $ **FLOATING
C766 a_18179_8983# VGND 0.804f $ **FLOATING
C767 a_17543_8751# VGND 0.609f $ **FLOATING
C768 a_17711_8725# VGND 0.817f $ **FLOATING
C769 a_17118_8751# VGND 0.626f $ **FLOATING
C770 a_17286_8725# VGND 0.581f $ **FLOATING
C771 a_16845_8757# VGND 1.43f $ **FLOATING
C772 a_16679_8757# VGND 1.81f $ **FLOATING
C773 a_14952_8751# VGND 1.37f $ **FLOATING
C774 _031_ VGND 3.54f $ **FLOATING
C775 _018_ VGND 1.27f $ **FLOATING
C776 a_14195_8867# VGND 0.702f $ **FLOATING
C777 _017_ VGND 2.16f $ **FLOATING
C778 _011_ VGND 0.796f $ **FLOATING
C779 a_12210_9071# VGND 0.482f $ **FLOATING
C780 a_13459_8751# VGND 0.804f $ **FLOATING
C781 _009_ VGND 2.49f $ **FLOATING
C782 tdc0.o_result\[84\] VGND 7.68f $ **FLOATING
C783 a_12376_8751# VGND 1.37f $ **FLOATING
C784 _051_ VGND 1.62f $ **FLOATING
C785 a_11619_8867# VGND 0.702f $ **FLOATING
C786 _074_ VGND 2.86f $ **FLOATING
C787 _075_ VGND 0.928f $ **FLOATING
C788 _073_ VGND 0.757f $ **FLOATING
C789 _049_ VGND 2.15f $ **FLOATING
C790 a_4617_8751# VGND 0.206f $ **FLOATING
C791 a_7925_8751# VGND 0.23f $ **FLOATING
C792 tdc0.w_dly_sig\[66\] VGND 3.79f $ **FLOATING
C793 tdc0.w_dly_sig_n\[64\] VGND 2.7f $ **FLOATING
C794 a_3417_8751# VGND 0.23f $ **FLOATING
C795 tdc0.o_result\[73\] VGND 4.54f $ **FLOATING
C796 a_1945_8751# VGND 0.23f $ **FLOATING
C797 a_10975_8751# VGND 0.804f $ **FLOATING
C798 tdc0.o_result\[65\] VGND 2.42f $ **FLOATING
C799 a_10239_8751# VGND 0.804f $ **FLOATING
C800 tdc0.o_result\[94\] VGND 2.87f $ **FLOATING
C801 a_9043_8751# VGND 0.804f $ **FLOATING
C802 tdc0.o_result\[33\] VGND 0.878f $ **FLOATING
C803 _028_ VGND 8.07f $ **FLOATING
C804 tdc0.o_result\[89\] VGND 3.79f $ **FLOATING
C805 a_8435_8751# VGND 0.609f $ **FLOATING
C806 a_8603_8725# VGND 0.817f $ **FLOATING
C807 a_8010_8751# VGND 0.626f $ **FLOATING
C808 a_8178_8725# VGND 0.581f $ **FLOATING
C809 a_7737_8757# VGND 1.43f $ **FLOATING
C810 a_7571_8757# VGND 1.81f $ **FLOATING
C811 a_4535_8751# VGND 0.804f $ **FLOATING
C812 _010_ VGND 13f $ **FLOATING
C813 tdc0.o_result\[81\] VGND 3.7f $ **FLOATING
C814 a_3927_8751# VGND 0.609f $ **FLOATING
C815 a_4095_8725# VGND 0.817f $ **FLOATING
C816 a_3502_8751# VGND 0.626f $ **FLOATING
C817 a_3670_8725# VGND 0.581f $ **FLOATING
C818 a_3229_8757# VGND 1.43f $ **FLOATING
C819 tdc0.w_dly_sig\[71\] VGND 3.25f $ **FLOATING
C820 a_3063_8757# VGND 1.81f $ **FLOATING
C821 a_2455_8751# VGND 0.609f $ **FLOATING
C822 a_2623_8725# VGND 0.817f $ **FLOATING
C823 a_2030_8751# VGND 0.626f $ **FLOATING
C824 a_2198_8725# VGND 0.581f $ **FLOATING
C825 a_1757_8757# VGND 1.43f $ **FLOATING
C826 tdc0.w_dly_sig\[74\] VGND 2.9f $ **FLOATING
C827 a_1591_8757# VGND 1.81f $ **FLOATING
C828 tdc0.o_result\[119\] VGND 1.13f $ **FLOATING
C829 a_17493_9295# VGND 0.23f $ **FLOATING
C830 a_18003_9661# VGND 0.609f $ **FLOATING
C831 a_18171_9563# VGND 0.817f $ **FLOATING
C832 a_17578_9661# VGND 0.626f $ **FLOATING
C833 a_17746_9407# VGND 0.581f $ **FLOATING
C834 a_17305_9295# VGND 1.43f $ **FLOATING
C835 a_17139_9295# VGND 1.81f $ **FLOATING
C836 a_12118_9295# VGND 0.482f $ **FLOATING
C837 tdc0.w_dly_sig\[118\] VGND 3.54f $ **FLOATING
C838 clknet_4_11_0_clk VGND 6.88f $ **FLOATING
C839 a_15453_9295# VGND 0.23f $ **FLOATING
C840 tdc0.o_result\[4\] VGND 1.27f $ **FLOATING
C841 _014_ VGND 0.89f $ **FLOATING
C842 a_13817_9545# VGND 0.206f $ **FLOATING
C843 a_12552_9545# VGND 0.14f $ **FLOATING
C844 a_12200_9545# VGND 0.171f $ **FLOATING
C845 a_11149_9545# VGND 0.206f $ **FLOATING
C846 tdc0.o_result\[30\] VGND 0.966f $ **FLOATING
C847 a_9397_9295# VGND 0.23f $ **FLOATING
C848 a_15035_9295# VGND 0.581f $ **FLOATING
C849 a_15106_9269# VGND 0.626f $ **FLOATING
C850 a_14899_9269# VGND 1.81f $ **FLOATING
C851 a_14906_9569# VGND 1.43f $ **FLOATING
C852 a_14615_9269# VGND 0.609f $ **FLOATING
C853 a_14519_9447# VGND 0.817f $ **FLOATING
C854 a_13735_9545# VGND 0.804f $ **FLOATING
C855 a_12284_9545# VGND 1.37f $ **FLOATING
C856 _076_ VGND 1.32f $ **FLOATING
C857 a_11067_9545# VGND 0.804f $ **FLOATING
C858 a_9907_9661# VGND 0.609f $ **FLOATING
C859 a_10075_9563# VGND 0.817f $ **FLOATING
C860 a_9482_9661# VGND 0.626f $ **FLOATING
C861 a_9650_9407# VGND 0.581f $ **FLOATING
C862 a_9209_9295# VGND 1.43f $ **FLOATING
C863 a_9043_9295# VGND 1.81f $ **FLOATING
C864 clknet_4_3_0_clk VGND 8.55f $ **FLOATING
C865 tdc0.o_result\[60\] VGND 3.13f $ **FLOATING
C866 a_7005_9295# VGND 0.23f $ **FLOATING
C867 a_7515_9661# VGND 0.609f $ **FLOATING
C868 a_7683_9563# VGND 0.817f $ **FLOATING
C869 a_7090_9661# VGND 0.626f $ **FLOATING
C870 a_7258_9407# VGND 0.581f $ **FLOATING
C871 a_6817_9295# VGND 1.43f $ **FLOATING
C872 a_6651_9295# VGND 1.81f $ **FLOATING
C873 _048_ VGND 4.86f $ **FLOATING
C874 a_5169_9545# VGND 0.206f $ **FLOATING
C875 a_1393_9295# VGND 0.23f $ **FLOATING
C876 a_5087_9545# VGND 0.804f $ **FLOATING
C877 net7 VGND 8.06f $ **FLOATING
C878 tdc0.o_result\[70\] VGND 1.47f $ **FLOATING
C879 tdc0.w_dly_sig_n\[63\] VGND 2.46f $ **FLOATING
C880 a_1903_9661# VGND 0.609f $ **FLOATING
C881 a_2071_9563# VGND 0.817f $ **FLOATING
C882 a_1478_9661# VGND 0.626f $ **FLOATING
C883 a_1646_9407# VGND 0.581f $ **FLOATING
C884 a_1205_9295# VGND 1.43f $ **FLOATING
C885 tdc0.w_dly_sig\[76\] VGND 3.37f $ **FLOATING
C886 a_1039_9295# VGND 1.81f $ **FLOATING
C887 clknet_4_1_0_clk VGND 10.2f $ **FLOATING
C888 a_18489_10217# VGND 0.23f $ **FLOATING
C889 a_16600_9839# VGND 0.14f $ **FLOATING
C890 a_16248_9839# VGND 0.171f $ **FLOATING
C891 tdc0.o_result\[121\] VGND 3.8f $ **FLOATING
C892 a_16166_10159# VGND 0.482f $ **FLOATING
C893 a_14349_10217# VGND 0.23f $ **FLOATING
C894 tdc0.o_result\[6\] VGND 1.83f $ **FLOATING
C895 a_18071_10217# VGND 0.581f $ **FLOATING
C896 a_18142_10116# VGND 0.626f $ **FLOATING
C897 a_17942_9961# VGND 1.43f $ **FLOATING
C898 a_17935_10057# VGND 1.81f $ **FLOATING
C899 a_17651_10071# VGND 0.609f $ **FLOATING
C900 a_17555_10071# VGND 0.817f $ **FLOATING
C901 a_16332_9839# VGND 1.37f $ **FLOATING
C902 _096_ VGND 1.73f $ **FLOATING
C903 a_13931_10217# VGND 0.581f $ **FLOATING
C904 a_14002_10116# VGND 0.626f $ **FLOATING
C905 a_13802_9961# VGND 1.43f $ **FLOATING
C906 a_13795_10057# VGND 1.81f $ **FLOATING
C907 a_13511_10071# VGND 0.609f $ **FLOATING
C908 a_13415_10071# VGND 0.817f $ **FLOATING
C909 a_11058_9839# VGND 4.03f $ **FLOATING
C910 _080_ VGND 3.9f $ **FLOATING
C911 _079_ VGND 1.05f $ **FLOATING
C912 _077_ VGND 3.14f $ **FLOATING
C913 _081_ VGND 2.67f $ **FLOATING
C914 tdc0.o_result\[62\] VGND 2.07f $ **FLOATING
C915 a_7097_9839# VGND 0.23f $ **FLOATING
C916 tdc0.w_dly_sig_n\[62\] VGND 2.06f $ **FLOATING
C917 a_1577_9839# VGND 0.23f $ **FLOATING
C918 a_9366_10071# VGND 0.702f $ **FLOATING
C919 a_7607_9839# VGND 0.609f $ **FLOATING
C920 a_7775_9813# VGND 0.817f $ **FLOATING
C921 a_7182_9839# VGND 0.626f $ **FLOATING
C922 a_7350_9813# VGND 0.581f $ **FLOATING
C923 a_6909_9845# VGND 1.43f $ **FLOATING
C924 tdc0.w_dly_sig\[63\] VGND 3.96f $ **FLOATING
C925 a_6743_9845# VGND 1.81f $ **FLOATING
C926 tdc0.w_dly_sig\[61\] VGND 2.8f $ **FLOATING
C927 a_2087_9839# VGND 0.609f $ **FLOATING
C928 a_2255_9813# VGND 0.817f $ **FLOATING
C929 a_1662_9839# VGND 0.626f $ **FLOATING
C930 a_1830_9813# VGND 0.581f $ **FLOATING
C931 a_1389_9845# VGND 1.43f $ **FLOATING
C932 tdc0.w_dly_sig\[78\] VGND 4.91f $ **FLOATING
C933 a_1223_9845# VGND 1.81f $ **FLOATING
C934 tdc0.w_dly_sig\[120\] VGND 3.38f $ **FLOATING
C935 a_17753_10383# VGND 0.23f $ **FLOATING
C936 tdc0.o_result\[1\] VGND 3.52f $ **FLOATING
C937 tdc0.o_result\[3\] VGND 1.29f $ **FLOATING
C938 a_15653_10383# VGND 0.23f $ **FLOATING
C939 a_17335_10383# VGND 0.581f $ **FLOATING
C940 a_17406_10357# VGND 0.626f $ **FLOATING
C941 a_17199_10357# VGND 1.81f $ **FLOATING
C942 a_17206_10657# VGND 1.43f $ **FLOATING
C943 a_16915_10357# VGND 0.609f $ **FLOATING
C944 a_16819_10535# VGND 0.817f $ **FLOATING
C945 a_16163_10749# VGND 0.609f $ **FLOATING
C946 a_16331_10651# VGND 0.817f $ **FLOATING
C947 a_15738_10749# VGND 0.626f $ **FLOATING
C948 a_15906_10495# VGND 0.581f $ **FLOATING
C949 a_15465_10383# VGND 1.43f $ **FLOATING
C950 a_15299_10383# VGND 1.81f $ **FLOATING
C951 _046_ VGND 1.73f $ **FLOATING
C952 _044_ VGND 3.54f $ **FLOATING
C953 _045_ VGND 3.27f $ **FLOATING
C954 _043_ VGND 1.42f $ **FLOATING
C955 _039_ VGND 4.11f $ **FLOATING
C956 _038_ VGND 5.54f $ **FLOATING
C957 _037_ VGND 0.994f $ **FLOATING
C958 a_10321_10633# VGND 0.206f $ **FLOATING
C959 a_9959_10633# VGND 0.253f $ **FLOATING
C960 _101_ VGND 5.25f $ **FLOATING
C961 _097_ VGND 2.64f $ **FLOATING
C962 a_3601_10383# VGND 0.23f $ **FLOATING
C963 a_11987_10633# VGND 0.702f $ **FLOATING
C964 a_11435_10633# VGND 0.702f $ **FLOATING
C965 a_10239_10633# VGND 0.804f $ **FLOATING
C966 tdc0.o_result\[77\] VGND 4.19f $ **FLOATING
C967 tdc0.o_result\[53\] VGND 2.96f $ **FLOATING
C968 a_9741_10357# VGND 0.55f $ **FLOATING
C969 a_6467_10633# VGND 0.702f $ **FLOATING
C970 tdc0.w_dly_sig_n\[61\] VGND 2.67f $ **FLOATING
C971 a_4111_10749# VGND 0.609f $ **FLOATING
C972 a_4279_10651# VGND 0.817f $ **FLOATING
C973 a_3686_10749# VGND 0.626f $ **FLOATING
C974 a_3854_10495# VGND 0.581f $ **FLOATING
C975 a_3413_10383# VGND 1.43f $ **FLOATING
C976 a_3247_10383# VGND 1.81f $ **FLOATING
C977 _100_ VGND 2.05f $ **FLOATING
C978 a_2593_10633# VGND 0.206f $ **FLOATING
C979 a_2511_10633# VGND 0.804f $ **FLOATING
C980 tdc0.o_result\[75\] VGND 1.02f $ **FLOATING
C981 a_13705_11305# VGND 0.23f $ **FLOATING
C982 a_11724_10927# VGND 0.14f $ **FLOATING
C983 a_11372_10927# VGND 0.171f $ **FLOATING
C984 a_10057_10927# VGND 0.253f $ **FLOATING
C985 a_11290_11247# VGND 0.482f $ **FLOATING
C986 a_18187_10901# VGND 2.1f $ **FLOATING
C987 tdc0.w_dly_sig_n\[117\] VGND 3.75f $ **FLOATING
C988 tdc0.w_dly_sig\[7\] VGND 2.91f $ **FLOATING
C989 a_13287_11305# VGND 0.581f $ **FLOATING
C990 a_13358_11204# VGND 0.626f $ **FLOATING
C991 a_13158_11049# VGND 1.43f $ **FLOATING
C992 a_13151_11145# VGND 1.81f $ **FLOATING
C993 a_12867_11159# VGND 0.609f $ **FLOATING
C994 a_12771_11159# VGND 0.817f $ **FLOATING
C995 a_11456_10927# VGND 1.37f $ **FLOATING
C996 _041_ VGND 0.958f $ **FLOATING
C997 _036_ VGND 1.69f $ **FLOATING
C998 tdc0.o_result\[5\] VGND 1.44f $ **FLOATING
C999 a_10226_11247# VGND 0.55f $ **FLOATING
C1000 _016_ VGND 5.51f $ **FLOATING
C1001 a_9503_11043# VGND 0.702f $ **FLOATING
C1002 _034_ VGND 0.832f $ **FLOATING
C1003 _035_ VGND 3.51f $ **FLOATING
C1004 a_8017_10927# VGND 0.23f $ **FLOATING
C1005 a_6545_10927# VGND 0.23f $ **FLOATING
C1006 tdc0.w_dly_sig_n\[60\] VGND 2.39f $ **FLOATING
C1007 tdc0.o_result\[55\] VGND 3.04f $ **FLOATING
C1008 a_3785_10927# VGND 0.23f $ **FLOATING
C1009 tdc0.o_result\[51\] VGND 1.15f $ **FLOATING
C1010 a_1853_10927# VGND 0.23f $ **FLOATING
C1011 a_8527_10927# VGND 0.609f $ **FLOATING
C1012 a_8695_10901# VGND 0.817f $ **FLOATING
C1013 a_8102_10927# VGND 0.626f $ **FLOATING
C1014 a_8270_10901# VGND 0.581f $ **FLOATING
C1015 a_7829_10933# VGND 1.43f $ **FLOATING
C1016 tdc0.w_dly_sig\[62\] VGND 3.76f $ **FLOATING
C1017 a_7663_10933# VGND 1.81f $ **FLOATING
C1018 a_7055_10927# VGND 0.609f $ **FLOATING
C1019 a_7223_10901# VGND 0.817f $ **FLOATING
C1020 a_6630_10927# VGND 0.626f $ **FLOATING
C1021 a_6798_10901# VGND 0.581f $ **FLOATING
C1022 a_6357_10933# VGND 1.43f $ **FLOATING
C1023 a_6191_10933# VGND 1.81f $ **FLOATING
C1024 a_4295_10927# VGND 0.609f $ **FLOATING
C1025 a_4463_10901# VGND 0.817f $ **FLOATING
C1026 a_3870_10927# VGND 0.626f $ **FLOATING
C1027 a_4038_10901# VGND 0.581f $ **FLOATING
C1028 a_3597_10933# VGND 1.43f $ **FLOATING
C1029 a_3431_10933# VGND 1.81f $ **FLOATING
C1030 a_2363_10927# VGND 0.609f $ **FLOATING
C1031 a_2531_10901# VGND 0.817f $ **FLOATING
C1032 a_1938_10927# VGND 0.626f $ **FLOATING
C1033 a_2106_10901# VGND 0.581f $ **FLOATING
C1034 a_1665_10933# VGND 1.43f $ **FLOATING
C1035 a_1499_10933# VGND 1.81f $ **FLOATING
C1036 a_11892_11471# VGND 0.482f $ **FLOATING
C1037 tdc0.w_dly_sig_n\[119\] VGND 2.53f $ **FLOATING
C1038 tdc0.w_dly_sig\[119\] VGND 4.51f $ **FLOATING
C1039 tdc0.w_dly_sig\[2\] VGND 3.23f $ **FLOATING
C1040 _356_.X VGND 0.226f $ **FLOATING
C1041 tdc0.w_dly_sig\[4\] VGND 2.98f $ **FLOATING
C1042 a_12326_11721# VGND 0.171f $ **FLOATING
C1043 a_11974_11721# VGND 0.14f $ **FLOATING
C1044 _052_ VGND 4.82f $ **FLOATING
C1045 _054_ VGND 1.07f $ **FLOATING
C1046 _055_ VGND 3.17f $ **FLOATING
C1047 _033_ VGND 1.4f $ **FLOATING
C1048 a_9677_11721# VGND 0.206f $ **FLOATING
C1049 _099_ VGND 2.04f $ **FLOATING
C1050 a_8481_11721# VGND 0.206f $ **FLOATING
C1051 tdc0.w_dly_sig\[60\] VGND 2.6f $ **FLOATING
C1052 tdc0.w_dly_sig_n\[59\] VGND 2.45f $ **FLOATING
C1053 a_1393_11471# VGND 0.23f $ **FLOATING
C1054 a_16732_11445# VGND 0.648f $ **FLOATING
C1055 tdc0.w_dly_sig_n\[4\] VGND 2.53f $ **FLOATING
C1056 tdc0.w_dly_sig_n\[5\] VGND 1.85f $ **FLOATING
C1057 tdc0.w_dly_sig_n\[6\] VGND 2.25f $ **FLOATING
C1058 tdc0.w_dly_sig\[6\] VGND 3.39f $ **FLOATING
C1059 _056_ VGND 1.12f $ **FLOATING
C1060 a_11504_11445# VGND 1.37f $ **FLOATING
C1061 a_10883_11721# VGND 0.702f $ **FLOATING
C1062 a_9595_11721# VGND 0.804f $ **FLOATING
C1063 tdc0.o_result\[61\] VGND 1.01f $ **FLOATING
C1064 a_8399_11721# VGND 0.804f $ **FLOATING
C1065 tdc0.o_result\[59\] VGND 1.12f $ **FLOATING
C1066 tdc0.w_dly_sig\[59\] VGND 4.47f $ **FLOATING
C1067 a_1903_11837# VGND 0.609f $ **FLOATING
C1068 a_2071_11739# VGND 0.817f $ **FLOATING
C1069 a_1478_11837# VGND 0.626f $ **FLOATING
C1070 a_1646_11583# VGND 0.581f $ **FLOATING
C1071 a_1205_11471# VGND 1.43f $ **FLOATING
C1072 tdc0.w_dly_sig\[73\] VGND 4.28f $ **FLOATING
C1073 a_1039_11471# VGND 1.81f $ **FLOATING
C1074 a_18581_12393# VGND 0.23f $ **FLOATING
C1075 a_16600_12015# VGND 0.14f $ **FLOATING
C1076 a_16248_12015# VGND 0.171f $ **FLOATING
C1077 a_16166_12335# VGND 0.482f $ **FLOATING
C1078 tdc0.w_dly_sig_n\[3\] VGND 2.2f $ **FLOATING
C1079 tdc0.w_dly_sig\[5\] VGND 3.93f $ **FLOATING
C1080 tdc0.w_dly_sig_n\[1\] VGND 2.67f $ **FLOATING
C1081 a_13429_12393# VGND 0.23f $ **FLOATING
C1082 tdc0.o_result\[7\] VGND 1.28f $ **FLOATING
C1083 a_11957_12393# VGND 0.23f $ **FLOATING
C1084 a_10321_12015# VGND 0.206f $ **FLOATING
C1085 a_9401_12015# VGND 0.206f $ **FLOATING
C1086 tdc0.o_result\[9\] VGND 1.98f $ **FLOATING
C1087 _078_ VGND 2.03f $ **FLOATING
C1088 a_8201_12015# VGND 0.23f $ **FLOATING
C1089 a_3329_12015# VGND 0.206f $ **FLOATING
C1090 a_2685_12015# VGND 0.206f $ **FLOATING
C1091 a_6177_12015# VGND 0.23f $ **FLOATING
C1092 tdc0.w_dly_sig_n\[58\] VGND 2.62f $ **FLOATING
C1093 tdc0.w_dly_sig_n\[57\] VGND 2.18f $ **FLOATING
C1094 tdc0.w_dly_sig\[56\] VGND 2.69f $ **FLOATING
C1095 a_1301_12015# VGND 0.23f $ **FLOATING
C1096 a_18163_12393# VGND 0.581f $ **FLOATING
C1097 a_18234_12292# VGND 0.626f $ **FLOATING
C1098 a_18034_12137# VGND 1.43f $ **FLOATING
C1099 a_18027_12233# VGND 1.81f $ **FLOATING
C1100 a_17743_12247# VGND 0.609f $ **FLOATING
C1101 a_17647_12247# VGND 0.817f $ **FLOATING
C1102 a_16332_12015# VGND 1.37f $ **FLOATING
C1103 _066_ VGND 3.48f $ **FLOATING
C1104 tdc0.w_dly_sig_n\[7\] VGND 2.4f $ **FLOATING
C1105 tdc0.w_dly_sig\[8\] VGND 2.93f $ **FLOATING
C1106 a_13011_12393# VGND 0.581f $ **FLOATING
C1107 a_13082_12292# VGND 0.626f $ **FLOATING
C1108 a_12882_12137# VGND 1.43f $ **FLOATING
C1109 a_12875_12233# VGND 1.81f $ **FLOATING
C1110 a_12591_12247# VGND 0.609f $ **FLOATING
C1111 a_12495_12247# VGND 0.817f $ **FLOATING
C1112 a_11539_12393# VGND 0.581f $ **FLOATING
C1113 a_11610_12292# VGND 0.626f $ **FLOATING
C1114 a_11410_12137# VGND 1.43f $ **FLOATING
C1115 a_11403_12233# VGND 1.81f $ **FLOATING
C1116 a_11119_12247# VGND 0.609f $ **FLOATING
C1117 a_11023_12247# VGND 0.817f $ **FLOATING
C1118 a_10239_12015# VGND 0.804f $ **FLOATING
C1119 net28 VGND 4.6f $ **FLOATING
C1120 tdc0.o_result\[79\] VGND 6.78f $ **FLOATING
C1121 a_9319_12015# VGND 0.804f $ **FLOATING
C1122 tdc0.o_result\[57\] VGND 1.49f $ **FLOATING
C1123 a_8711_12015# VGND 0.609f $ **FLOATING
C1124 a_8879_11989# VGND 0.817f $ **FLOATING
C1125 a_8286_12015# VGND 0.626f $ **FLOATING
C1126 a_8454_11989# VGND 0.581f $ **FLOATING
C1127 a_8013_12021# VGND 1.43f $ **FLOATING
C1128 tdc0.w_dly_sig\[64\] VGND 5.21f $ **FLOATING
C1129 a_7847_12021# VGND 1.81f $ **FLOATING
C1130 a_6687_12015# VGND 0.609f $ **FLOATING
C1131 a_6855_11989# VGND 0.817f $ **FLOATING
C1132 a_6262_12015# VGND 0.626f $ **FLOATING
C1133 a_6430_11989# VGND 0.581f $ **FLOATING
C1134 a_5989_12021# VGND 1.43f $ **FLOATING
C1135 tdc0.w_dly_sig\[58\] VGND 3.4f $ **FLOATING
C1136 a_5823_12021# VGND 1.81f $ **FLOATING
C1137 a_3247_12015# VGND 0.804f $ **FLOATING
C1138 tdc0.o_result\[74\] VGND 0.978f $ **FLOATING
C1139 a_2603_12015# VGND 0.804f $ **FLOATING
C1140 _026_ VGND 13.5f $ **FLOATING
C1141 tdc0.o_result\[72\] VGND 0.876f $ **FLOATING
C1142 a_1811_12015# VGND 0.609f $ **FLOATING
C1143 a_1979_11989# VGND 0.817f $ **FLOATING
C1144 a_1386_12015# VGND 0.626f $ **FLOATING
C1145 a_1554_11989# VGND 0.581f $ **FLOATING
C1146 a_1113_12021# VGND 1.43f $ **FLOATING
C1147 tdc0.w_dly_sig\[75\] VGND 5.57f $ **FLOATING
C1148 a_947_12021# VGND 1.81f $ **FLOATING
C1149 a_14510_12559# VGND 0.482f $ **FLOATING
C1150 a_17314_12559# VGND 1.98f $ **FLOATING
C1151 clknet_4_14_0_clk VGND 8.74f $ **FLOATING
C1152 a_16741_12559# VGND 0.23f $ **FLOATING
C1153 tdc0.o_result\[0\] VGND 1.3f $ **FLOATING
C1154 a_14944_12809# VGND 0.14f $ **FLOATING
C1155 a_14592_12809# VGND 0.171f $ **FLOATING
C1156 _061_ VGND 1.57f $ **FLOATING
C1157 _057_ VGND 0.823f $ **FLOATING
C1158 _060_ VGND 5.3f $ **FLOATING
C1159 _058_ VGND 1.18f $ **FLOATING
C1160 a_9493_12809# VGND 0.206f $ **FLOATING
C1161 a_8481_12809# VGND 0.206f $ **FLOATING
C1162 _071_ VGND 4.76f $ **FLOATING
C1163 _067_ VGND 3.27f $ **FLOATING
C1164 _069_ VGND 1.06f $ **FLOATING
C1165 _070_ VGND 2.92f $ **FLOATING
C1166 _087_ VGND 3.64f $ **FLOATING
C1167 _090_ VGND 2.09f $ **FLOATING
C1168 a_5717_12559# VGND 0.23f $ **FLOATING
C1169 a_16323_12559# VGND 0.581f $ **FLOATING
C1170 a_16394_12533# VGND 0.626f $ **FLOATING
C1171 a_16187_12533# VGND 1.81f $ **FLOATING
C1172 a_16194_12833# VGND 1.43f $ **FLOATING
C1173 a_15903_12533# VGND 0.609f $ **FLOATING
C1174 a_15807_12711# VGND 0.817f $ **FLOATING
C1175 a_14676_12809# VGND 1.37f $ **FLOATING
C1176 _091_ VGND 4.32f $ **FLOATING
C1177 _086_ VGND 4.58f $ **FLOATING
C1178 _005_ VGND 11.7f $ **FLOATING
C1179 tdc0.w_dly_sig_n\[8\] VGND 2.37f $ **FLOATING
C1180 tdc0.w_dly_sig\[9\] VGND 6.22f $ **FLOATING
C1181 tdc0.w_dly_sig\[10\] VGND 3.51f $ **FLOATING
C1182 a_10607_12809# VGND 0.702f $ **FLOATING
C1183 a_9411_12809# VGND 0.804f $ **FLOATING
C1184 tdc0.o_result\[63\] VGND 0.85f $ **FLOATING
C1185 a_8399_12809# VGND 0.804f $ **FLOATING
C1186 tdc0.o_result\[120\] VGND 4.74f $ **FLOATING
C1187 _013_ VGND 11f $ **FLOATING
C1188 tdc0.o_result\[56\] VGND 1.35f $ **FLOATING
C1189 a_7755_12809# VGND 0.702f $ **FLOATING
C1190 a_6835_12809# VGND 0.702f $ **FLOATING
C1191 a_6227_12925# VGND 0.609f $ **FLOATING
C1192 a_6395_12827# VGND 0.817f $ **FLOATING
C1193 a_5802_12925# VGND 0.626f $ **FLOATING
C1194 a_5970_12671# VGND 0.581f $ **FLOATING
C1195 a_5529_12559# VGND 1.43f $ **FLOATING
C1196 a_5363_12559# VGND 1.81f $ **FLOATING
C1197 tdc0.w_dly_sig\[57\] VGND 3.16f $ **FLOATING
C1198 tdc0.w_dly_sig_n\[56\] VGND 2.69f $ **FLOATING
C1199 tdc0.w_dly_sig_n\[55\] VGND 2.73f $ **FLOATING
C1200 a_3698_12559# VGND 1.98f $ **FLOATING
C1201 tdc0.w_dly_sig\[54\] VGND 3.4f $ **FLOATING
C1202 tdc0.w_dly_sig_n\[2\] VGND 2.64f $ **FLOATING
C1203 a_15545_13481# VGND 0.23f $ **FLOATING
C1204 tdc0.o_result\[2\] VGND 1.23f $ **FLOATING
C1205 a_11957_13481# VGND 0.23f $ **FLOATING
C1206 tdc0.o_result\[13\] VGND 1.89f $ **FLOATING
C1207 tdc0.o_result\[31\] VGND 1.01f $ **FLOATING
C1208 a_7561_13103# VGND 0.206f $ **FLOATING
C1209 a_5997_13103# VGND 0.206f $ **FLOATING
C1210 a_9029_13103# VGND 0.23f $ **FLOATING
C1211 _024_ VGND 3.04f $ **FLOATING
C1212 _042_ VGND 4.57f $ **FLOATING
C1213 a_4613_13103# VGND 0.23f $ **FLOATING
C1214 tdc0.o_result\[50\] VGND 1.45f $ **FLOATING
C1215 a_1485_13103# VGND 0.23f $ **FLOATING
C1216 net1 VGND 5.21f $ **FLOATING
C1217 a_16578_13103# VGND 1.98f $ **FLOATING
C1218 tdc0.w_dly_sig_n\[0\] VGND 4.16f $ **FLOATING
C1219 a_15127_13481# VGND 0.581f $ **FLOATING
C1220 a_15198_13380# VGND 0.626f $ **FLOATING
C1221 a_14998_13225# VGND 1.43f $ **FLOATING
C1222 a_14991_13321# VGND 1.81f $ **FLOATING
C1223 a_14707_13335# VGND 0.609f $ **FLOATING
C1224 a_14611_13335# VGND 0.817f $ **FLOATING
C1225 tdc0.w_dly_sig_n\[9\] VGND 2.46f $ **FLOATING
C1226 tdc0.w_dly_sig_n\[10\] VGND 2.08f $ **FLOATING
C1227 tdc0.w_dly_sig\[11\] VGND 7.7f $ **FLOATING
C1228 a_11539_13481# VGND 0.581f $ **FLOATING
C1229 a_11610_13380# VGND 0.626f $ **FLOATING
C1230 a_11410_13225# VGND 1.43f $ **FLOATING
C1231 a_11403_13321# VGND 1.81f $ **FLOATING
C1232 a_11119_13335# VGND 0.609f $ **FLOATING
C1233 a_11023_13335# VGND 0.817f $ **FLOATING
C1234 a_9539_13103# VGND 0.609f $ **FLOATING
C1235 a_9707_13077# VGND 0.817f $ **FLOATING
C1236 a_9114_13103# VGND 0.626f $ **FLOATING
C1237 a_9282_13077# VGND 0.581f $ **FLOATING
C1238 a_8841_13109# VGND 1.43f $ **FLOATING
C1239 a_8675_13109# VGND 1.81f $ **FLOATING
C1240 a_7479_13103# VGND 0.804f $ **FLOATING
C1241 a_6550_13103# VGND 1.98f $ **FLOATING
C1242 tdc0.o_result\[54\] VGND 0.929f $ **FLOATING
C1243 _022_ VGND 12.6f $ **FLOATING
C1244 a_5851_13335# VGND 0.804f $ **FLOATING
C1245 a_5123_13103# VGND 0.609f $ **FLOATING
C1246 a_5291_13077# VGND 0.817f $ **FLOATING
C1247 a_4698_13103# VGND 0.626f $ **FLOATING
C1248 a_4866_13077# VGND 0.581f $ **FLOATING
C1249 a_4425_13109# VGND 1.43f $ **FLOATING
C1250 a_4259_13109# VGND 1.81f $ **FLOATING
C1251 a_3348_13077# VGND 1.98f $ **FLOATING
C1252 a_1995_13103# VGND 0.609f $ **FLOATING
C1253 a_2163_13077# VGND 0.817f $ **FLOATING
C1254 a_1570_13103# VGND 0.626f $ **FLOATING
C1255 a_1738_13077# VGND 0.581f $ **FLOATING
C1256 a_1297_13109# VGND 1.43f $ **FLOATING
C1257 a_1131_13109# VGND 1.81f $ **FLOATING
C1258 clknet_4_4_0_clk VGND 10.1f $ **FLOATING
C1259 a_18121_13647# VGND 0.23f $ **FLOATING
C1260 tdc0.o_result\[123\] VGND 5.22f $ **FLOATING
C1261 tdc0.w_dly_sig\[3\] VGND 3.51f $ **FLOATING
C1262 a_15473_13897# VGND 0.206f $ **FLOATING
C1263 _008_ VGND 2.89f $ **FLOATING
C1264 tdc0.o_result\[36\] VGND 0.967f $ **FLOATING
C1265 a_5993_13647# VGND 0.23f $ **FLOATING
C1266 a_17703_13647# VGND 0.581f $ **FLOATING
C1267 a_17774_13621# VGND 0.626f $ **FLOATING
C1268 a_17567_13621# VGND 1.81f $ **FLOATING
C1269 a_17574_13921# VGND 1.43f $ **FLOATING
C1270 a_17283_13621# VGND 0.609f $ **FLOATING
C1271 a_17187_13799# VGND 0.817f $ **FLOATING
C1272 tdc0.w_dly_sig\[1\] VGND 5.47f $ **FLOATING
C1273 net11 VGND 5.44f $ **FLOATING
C1274 a_15327_13799# VGND 0.804f $ **FLOATING
C1275 a_14388_13621# VGND 1.98f $ **FLOATING
C1276 tdc0.w_dly_sig_n\[11\] VGND 2.33f $ **FLOATING
C1277 tdc0.w_dly_sig\[12\] VGND 5.59f $ **FLOATING
C1278 a_6503_14013# VGND 0.609f $ **FLOATING
C1279 a_6671_13915# VGND 0.817f $ **FLOATING
C1280 a_6078_14013# VGND 0.626f $ **FLOATING
C1281 a_6246_13759# VGND 0.581f $ **FLOATING
C1282 a_5805_13647# VGND 1.43f $ **FLOATING
C1283 a_5639_13647# VGND 1.81f $ **FLOATING
C1284 clknet_4_6_0_clk VGND 8.28f $ **FLOATING
C1285 tdc0.o_result\[52\] VGND 2.2f $ **FLOATING
C1286 a_4061_13647# VGND 0.23f $ **FLOATING
C1287 a_4571_14013# VGND 0.609f $ **FLOATING
C1288 a_4739_13915# VGND 0.817f $ **FLOATING
C1289 a_4146_14013# VGND 0.626f $ **FLOATING
C1290 a_4314_13759# VGND 0.581f $ **FLOATING
C1291 a_3873_13647# VGND 1.43f $ **FLOATING
C1292 a_3707_13647# VGND 1.81f $ **FLOATING
C1293 tdc0.w_dly_sig\[55\] VGND 3.86f $ **FLOATING
C1294 tdc0.w_dly_sig_n\[53\] VGND 3.17f $ **FLOATING
C1295 tdc0.w_dly_sig\[53\] VGND 3.09f $ **FLOATING
C1296 tdc0.w_dly_sig_n\[54\] VGND 2.44f $ **FLOATING
C1297 a_18397_14569# VGND 0.23f $ **FLOATING
C1298 a_16301_14191# VGND 0.206f $ **FLOATING
C1299 _089_ VGND 5.53f $ **FLOATING
C1300 tdc0.o_result\[12\] VGND 1.14f $ **FLOATING
C1301 a_13997_14191# VGND 0.23f $ **FLOATING
C1302 a_11957_14569# VGND 0.23f $ **FLOATING
C1303 tdc0.o_result\[14\] VGND 2.69f $ **FLOATING
C1304 tdc0.o_result\[29\] VGND 1.87f $ **FLOATING
C1305 a_9121_14191# VGND 0.23f $ **FLOATING
C1306 tdc0.w_dly_sig\[34\] VGND 4.63f $ **FLOATING
C1307 tdc0.o_result\[49\] VGND 3.11f $ **FLOATING
C1308 a_2497_14191# VGND 0.23f $ **FLOATING
C1309 tdc0.w_dly_sig_n\[52\] VGND 2.18f $ **FLOATING
C1310 tdc0.w_dly_sig\[52\] VGND 3.8f $ **FLOATING
C1311 tdc0.w_dly_sig\[121\] VGND 3.21f $ **FLOATING
C1312 a_17979_14569# VGND 0.581f $ **FLOATING
C1313 a_18050_14468# VGND 0.626f $ **FLOATING
C1314 a_17850_14313# VGND 1.43f $ **FLOATING
C1315 a_17843_14409# VGND 1.81f $ **FLOATING
C1316 a_17559_14423# VGND 0.609f $ **FLOATING
C1317 a_17463_14423# VGND 0.817f $ **FLOATING
C1318 tdc0.o_result\[122\] VGND 1.03f $ **FLOATING
C1319 a_16155_14423# VGND 0.804f $ **FLOATING
C1320 a_14507_14191# VGND 0.609f $ **FLOATING
C1321 a_14675_14165# VGND 0.817f $ **FLOATING
C1322 a_14082_14191# VGND 0.626f $ **FLOATING
C1323 a_14250_14165# VGND 0.581f $ **FLOATING
C1324 a_13809_14197# VGND 1.43f $ **FLOATING
C1325 a_13643_14197# VGND 1.81f $ **FLOATING
C1326 a_12548_14165# VGND 1.98f $ **FLOATING
C1327 a_11539_14569# VGND 0.581f $ **FLOATING
C1328 a_11610_14468# VGND 0.626f $ **FLOATING
C1329 a_11410_14313# VGND 1.43f $ **FLOATING
C1330 a_11403_14409# VGND 1.81f $ **FLOATING
C1331 a_11119_14423# VGND 0.609f $ **FLOATING
C1332 a_11023_14423# VGND 0.817f $ **FLOATING
C1333 a_9631_14191# VGND 0.609f $ **FLOATING
C1334 a_9799_14165# VGND 0.817f $ **FLOATING
C1335 a_9206_14191# VGND 0.626f $ **FLOATING
C1336 a_9374_14165# VGND 0.581f $ **FLOATING
C1337 a_8933_14197# VGND 1.43f $ **FLOATING
C1338 a_8767_14197# VGND 1.81f $ **FLOATING
C1339 clknet_0_clk VGND 31.8f $ **FLOATING
C1340 a_7856_14165# VGND 1.98f $ **FLOATING
C1341 tdc0.w_dly_sig\[35\] VGND 6.15f $ **FLOATING
C1342 a_3007_14191# VGND 0.609f $ **FLOATING
C1343 a_3175_14165# VGND 0.817f $ **FLOATING
C1344 a_2582_14191# VGND 0.626f $ **FLOATING
C1345 a_2750_14165# VGND 0.581f $ **FLOATING
C1346 a_2309_14197# VGND 1.43f $ **FLOATING
C1347 a_2143_14197# VGND 1.81f $ **FLOATING
C1348 tdc0.w_dly_sig_n\[121\] VGND 3.1f $ **FLOATING
C1349 tdc0.w_dly_sig_n\[120\] VGND 4.87f $ **FLOATING
C1350 a_17477_14735# VGND 0.23f $ **FLOATING
C1351 tdc0.o_result\[124\] VGND 1.28f $ **FLOATING
C1352 tdc0.o_result\[27\] VGND 3.2f $ **FLOATING
C1353 a_15377_14735# VGND 0.23f $ **FLOATING
C1354 a_17059_14735# VGND 0.581f $ **FLOATING
C1355 a_17130_14709# VGND 0.626f $ **FLOATING
C1356 a_16923_14709# VGND 1.81f $ **FLOATING
C1357 a_16930_15009# VGND 1.43f $ **FLOATING
C1358 a_16639_14709# VGND 0.609f $ **FLOATING
C1359 a_16543_14887# VGND 0.817f $ **FLOATING
C1360 a_15887_15101# VGND 0.609f $ **FLOATING
C1361 a_16055_15003# VGND 0.817f $ **FLOATING
C1362 a_15462_15101# VGND 0.626f $ **FLOATING
C1363 a_15630_14847# VGND 0.581f $ **FLOATING
C1364 a_15189_14735# VGND 1.43f $ **FLOATING
C1365 a_15023_14735# VGND 1.81f $ **FLOATING
C1366 a_14533_14735# VGND 0.23f $ **FLOATING
C1367 tdc0.o_result\[28\] VGND 2.94f $ **FLOATING
C1368 tdc0.w_dly_sig\[31\] VGND 5.27f $ **FLOATING
C1369 a_14115_14735# VGND 0.581f $ **FLOATING
C1370 a_14186_14709# VGND 0.626f $ **FLOATING
C1371 a_13979_14709# VGND 1.81f $ **FLOATING
C1372 a_13986_15009# VGND 1.43f $ **FLOATING
C1373 a_13695_14709# VGND 0.609f $ **FLOATING
C1374 a_13599_14887# VGND 0.817f $ **FLOATING
C1375 tdc0.w_dly_sig\[13\] VGND 3.67f $ **FLOATING
C1376 clknet_4_12_0_clk VGND 5.61f $ **FLOATING
C1377 a_10945_14735# VGND 0.23f $ **FLOATING
C1378 tdc0.o_result\[15\] VGND 1.94f $ **FLOATING
C1379 tdc0.w_dly_sig_n\[32\] VGND 3.16f $ **FLOATING
C1380 tdc0.o_result\[38\] VGND 1.23f $ **FLOATING
C1381 a_5441_14735# VGND 0.23f $ **FLOATING
C1382 a_10527_14735# VGND 0.581f $ **FLOATING
C1383 a_10598_14709# VGND 0.626f $ **FLOATING
C1384 a_10391_14709# VGND 1.81f $ **FLOATING
C1385 a_10398_15009# VGND 1.43f $ **FLOATING
C1386 a_10107_14709# VGND 0.609f $ **FLOATING
C1387 a_10011_14887# VGND 0.817f $ **FLOATING
C1388 tdc0.w_dly_sig_n\[31\] VGND 4.02f $ **FLOATING
C1389 tdc0.w_dly_sig\[32\] VGND 3.47f $ **FLOATING
C1390 tdc0.w_dly_sig\[33\] VGND 6.51f $ **FLOATING
C1391 tdc0.w_dly_sig_n\[34\] VGND 2.45f $ **FLOATING
C1392 tdc0.w_dly_sig_n\[33\] VGND 2.32f $ **FLOATING
C1393 tdc0.w_dly_sig_n\[35\] VGND 2.38f $ **FLOATING
C1394 a_5951_15101# VGND 0.609f $ **FLOATING
C1395 a_6119_15003# VGND 0.817f $ **FLOATING
C1396 a_5526_15101# VGND 0.626f $ **FLOATING
C1397 a_5694_14847# VGND 0.581f $ **FLOATING
C1398 a_5253_14735# VGND 1.43f $ **FLOATING
C1399 a_5087_14735# VGND 1.81f $ **FLOATING
C1400 tdc0.o_result\[46\] VGND 2.96f $ **FLOATING
C1401 a_3601_14735# VGND 0.23f $ **FLOATING
C1402 a_4111_15101# VGND 0.609f $ **FLOATING
C1403 a_4279_15003# VGND 0.817f $ **FLOATING
C1404 a_3686_15101# VGND 0.626f $ **FLOATING
C1405 a_3854_14847# VGND 0.581f $ **FLOATING
C1406 a_3413_14735# VGND 1.43f $ **FLOATING
C1407 a_3247_14735# VGND 1.81f $ **FLOATING
C1408 tdc0.w_dly_sig_n\[51\] VGND 2.93f $ **FLOATING
C1409 tdc0.o_result\[48\] VGND 2.02f $ **FLOATING
C1410 a_1577_14735# VGND 0.23f $ **FLOATING
C1411 a_2087_15101# VGND 0.609f $ **FLOATING
C1412 a_2255_15003# VGND 0.817f $ **FLOATING
C1413 a_1662_15101# VGND 0.626f $ **FLOATING
C1414 a_1830_14847# VGND 0.581f $ **FLOATING
C1415 a_1389_14735# VGND 1.43f $ **FLOATING
C1416 a_1223_14735# VGND 1.81f $ **FLOATING
C1417 tdc0.o_result\[26\] VGND 1.3f $ **FLOATING
C1418 a_11333_15279# VGND 0.206f $ **FLOATING
C1419 a_14917_15279# VGND 0.23f $ **FLOATING
C1420 tdc0.w_dly_sig_n\[30\] VGND 4.18f $ **FLOATING
C1421 tdc0.w_dly_sig\[30\] VGND 5.27f $ **FLOATING
C1422 _072_ VGND 3.41f $ **FLOATING
C1423 tdc0.o_result\[44\] VGND 4.88f $ **FLOATING
C1424 a_3877_15279# VGND 0.23f $ **FLOATING
C1425 tdc0.w_dly_sig_n\[50\] VGND 2.48f $ **FLOATING
C1426 tdc0.w_dly_sig\[51\] VGND 3.5f $ **FLOATING
C1427 tdc0.w_dly_sig\[122\] VGND 5.34f $ **FLOATING
C1428 tdc0.w_dly_sig_n\[122\] VGND 2.11f $ **FLOATING
C1429 tdc0.w_dly_sig\[123\] VGND 3.87f $ **FLOATING
C1430 tdc0.w_dly_sig_n\[123\] VGND 2.94f $ **FLOATING
C1431 a_15427_15279# VGND 0.609f $ **FLOATING
C1432 a_15595_15253# VGND 0.817f $ **FLOATING
C1433 a_15002_15279# VGND 0.626f $ **FLOATING
C1434 a_15170_15253# VGND 0.581f $ **FLOATING
C1435 a_14729_15285# VGND 1.43f $ **FLOATING
C1436 a_14563_15285# VGND 1.81f $ **FLOATING
C1437 tdc0.w_dly_sig_n\[12\] VGND 2.84f $ **FLOATING
C1438 tdc0.w_dly_sig_n\[13\] VGND 3.37f $ **FLOATING
C1439 a_11251_15279# VGND 0.804f $ **FLOATING
C1440 _012_ VGND 14.7f $ **FLOATING
C1441 tdc0.w_dly_sig\[14\] VGND 4.01f $ **FLOATING
C1442 tdc0.w_dly_sig\[36\] VGND 5.64f $ **FLOATING
C1443 tdc0.w_dly_sig_n\[36\] VGND 2.32f $ **FLOATING
C1444 tdc0.w_dly_sig\[37\] VGND 3.01f $ **FLOATING
C1445 tdc0.w_dly_sig_n\[37\] VGND 2.27f $ **FLOATING
C1446 a_4387_15279# VGND 0.609f $ **FLOATING
C1447 a_4555_15253# VGND 0.817f $ **FLOATING
C1448 a_3962_15279# VGND 0.626f $ **FLOATING
C1449 a_4130_15253# VGND 0.581f $ **FLOATING
C1450 a_3689_15285# VGND 1.43f $ **FLOATING
C1451 a_3523_15285# VGND 1.81f $ **FLOATING
C1452 tdc0.w_dly_sig\[124\] VGND 3.91f $ **FLOATING
C1453 a_15269_15823# VGND 0.23f $ **FLOATING
C1454 tdc0.o_result\[25\] VGND 2.06f $ **FLOATING
C1455 tdc0.w_dly_sig_n\[29\] VGND 2.73f $ **FLOATING
C1456 _059_ VGND 2.15f $ **FLOATING
C1457 a_10873_16073# VGND 0.206f $ **FLOATING
C1458 _040_ VGND 3.17f $ **FLOATING
C1459 a_10229_16073# VGND 0.206f $ **FLOATING
C1460 a_8753_15823# VGND 0.23f $ **FLOATING
C1461 a_14851_15823# VGND 0.581f $ **FLOATING
C1462 a_14922_15797# VGND 0.626f $ **FLOATING
C1463 a_14715_15797# VGND 1.81f $ **FLOATING
C1464 a_14722_16097# VGND 1.43f $ **FLOATING
C1465 a_14431_15797# VGND 0.609f $ **FLOATING
C1466 a_14335_15975# VGND 0.817f $ **FLOATING
C1467 a_10791_16073# VGND 0.804f $ **FLOATING
C1468 a_10147_16073# VGND 0.804f $ **FLOATING
C1469 net6 VGND 8.02f $ **FLOATING
C1470 tdc0.o_result\[37\] VGND 0.747f $ **FLOATING
C1471 a_9263_16189# VGND 0.609f $ **FLOATING
C1472 a_9431_16091# VGND 0.817f $ **FLOATING
C1473 a_8838_16189# VGND 0.626f $ **FLOATING
C1474 a_9006_15935# VGND 0.581f $ **FLOATING
C1475 a_8565_15823# VGND 1.43f $ **FLOATING
C1476 a_8399_15823# VGND 1.81f $ **FLOATING
C1477 tdc0.o_result\[41\] VGND 2.22f $ **FLOATING
C1478 a_6821_15823# VGND 0.23f $ **FLOATING
C1479 tdc0.w_dly_sig\[38\] VGND 3.15f $ **FLOATING
C1480 a_7331_16189# VGND 0.609f $ **FLOATING
C1481 a_7499_16091# VGND 0.817f $ **FLOATING
C1482 a_6906_16189# VGND 0.626f $ **FLOATING
C1483 a_7074_15935# VGND 0.581f $ **FLOATING
C1484 a_6633_15823# VGND 1.43f $ **FLOATING
C1485 a_6467_15823# VGND 1.81f $ **FLOATING
C1486 tdc0.w_dly_sig_n\[49\] VGND 2.56f $ **FLOATING
C1487 tdc0.w_dly_sig\[50\] VGND 3.27f $ **FLOATING
C1488 tdc0.w_dly_sig\[49\] VGND 2.95f $ **FLOATING
C1489 tdc0.w_dly_sig_n\[38\] VGND 2.61f $ **FLOATING
C1490 tdc0.w_dly_sig\[39\] VGND 3.07f $ **FLOATING
C1491 tt_um_hpretl_tt06_tdc_12.HI VGND 0.415f $ **FLOATING
C1492 a_18121_16745# VGND 0.23f $ **FLOATING
C1493 tdc0.o_result\[125\] VGND 3.86f $ **FLOATING
C1494 tdc0.w_dly_sig\[28\] VGND 3.89f $ **FLOATING
C1495 tdc0.w_dly_sig_n\[27\] VGND 2.88f $ **FLOATING
C1496 tdc0.w_dly_sig\[29\] VGND 4.52f $ **FLOATING
C1497 tdc0.w_dly_sig_n\[28\] VGND 2.12f $ **FLOATING
C1498 tdc0.o_result\[39\] VGND 1.48f $ **FLOATING
C1499 a_6181_16367# VGND 0.206f $ **FLOATING
C1500 a_8477_16367# VGND 0.23f $ **FLOATING
C1501 _098_ VGND 3.09f $ **FLOATING
C1502 tdc0.w_dly_sig\[47\] VGND 3.67f $ **FLOATING
C1503 tdc0.w_dly_sig_n\[48\] VGND 2.33f $ **FLOATING
C1504 a_17703_16745# VGND 0.581f $ **FLOATING
C1505 a_17774_16644# VGND 0.626f $ **FLOATING
C1506 a_17574_16489# VGND 1.43f $ **FLOATING
C1507 a_17567_16585# VGND 1.81f $ **FLOATING
C1508 a_17283_16599# VGND 0.609f $ **FLOATING
C1509 a_17187_16599# VGND 0.817f $ **FLOATING
C1510 tdc0.w_dly_sig\[125\] VGND 3.28f $ **FLOATING
C1511 tdc0.w_dly_sig\[27\] VGND 3.01f $ **FLOATING
C1512 tdc0.w_dly_sig_n\[14\] VGND 2.32f $ **FLOATING
C1513 tdc0.w_dly_sig\[15\] VGND 3.93f $ **FLOATING
C1514 a_8987_16367# VGND 0.609f $ **FLOATING
C1515 a_9155_16341# VGND 0.817f $ **FLOATING
C1516 a_8562_16367# VGND 0.626f $ **FLOATING
C1517 a_8730_16341# VGND 0.581f $ **FLOATING
C1518 a_8289_16373# VGND 1.43f $ **FLOATING
C1519 a_8123_16373# VGND 1.81f $ **FLOATING
C1520 a_6099_16367# VGND 0.804f $ **FLOATING
C1521 tdc0.w_dly_sig\[40\] VGND 4.12f $ **FLOATING
C1522 tdc0.w_dly_sig_n\[39\] VGND 2.2f $ **FLOATING
C1523 tdc0.w_dly_sig_n\[40\] VGND 2.3f $ **FLOATING
C1524 tdc0.w_dly_sig_n\[47\] VGND 2.24f $ **FLOATING
C1525 tdc0.w_dly_sig_n\[26\] VGND 2.33f $ **FLOATING
C1526 _068_ VGND 2.43f $ **FLOATING
C1527 a_7653_17161# VGND 0.206f $ **FLOATING
C1528 a_5901_16911# VGND 0.23f $ **FLOATING
C1529 tdc0.w_dly_sig_n\[127\] VGND 2.35f $ **FLOATING
C1530 tdc0.w_dly_sig_n\[125\] VGND 3.14f $ **FLOATING
C1531 tdc0.w_dly_sig_n\[124\] VGND 2.64f $ **FLOATING
C1532 tdc0.w_dly_sig\[126\] VGND 3.2f $ **FLOATING
C1533 tdc0.w_dly_sig_n\[126\] VGND 2.34f $ **FLOATING
C1534 tdc0.w_dly_sig\[26\] VGND 3.05f $ **FLOATING
C1535 tdc0.w_dly_sig_n\[15\] VGND 2.51f $ **FLOATING
C1536 tdc0.w_dly_sig_n\[16\] VGND 2.05f $ **FLOATING
C1537 tdc0.w_dly_sig\[16\] VGND 3.48f $ **FLOATING
C1538 a_9227_16911# VGND 0.524f $ **FLOATING
C1539 a_7571_17161# VGND 0.804f $ **FLOATING
C1540 tdc0.o_result\[40\] VGND 0.864f $ **FLOATING
C1541 a_6411_17277# VGND 0.609f $ **FLOATING
C1542 a_6579_17179# VGND 0.817f $ **FLOATING
C1543 a_5986_17277# VGND 0.626f $ **FLOATING
C1544 a_6154_17023# VGND 0.581f $ **FLOATING
C1545 a_5713_16911# VGND 1.43f $ **FLOATING
C1546 a_5547_16911# VGND 1.81f $ **FLOATING
C1547 tdc0.w_dly_sig\[45\] VGND 3.23f $ **FLOATING
C1548 tt_um_hpretl_tt06_tdc_14.HI VGND 0.415f $ **FLOATING
C1549 a_1945_16911# VGND 0.23f $ **FLOATING
C1550 tdc0.w_dly_sig\[41\] VGND 3.21f $ **FLOATING
C1551 tdc0.w_dly_sig_n\[41\] VGND 2.1f $ **FLOATING
C1552 tdc0.w_dly_sig\[42\] VGND 3.83f $ **FLOATING
C1553 tdc0.w_dly_sig_n\[42\] VGND 2.41f $ **FLOATING
C1554 a_2455_17277# VGND 0.609f $ **FLOATING
C1555 a_2623_17179# VGND 0.817f $ **FLOATING
C1556 a_2030_17277# VGND 0.626f $ **FLOATING
C1557 a_2198_17023# VGND 0.581f $ **FLOATING
C1558 a_1757_16911# VGND 1.43f $ **FLOATING
C1559 a_1591_16911# VGND 1.81f $ **FLOATING
C1560 tdc0.w_dly_sig\[129\] VGND 1.5f $ **FLOATING
C1561 a_18121_17833# VGND 0.23f $ **FLOATING
C1562 a_16301_17455# VGND 0.206f $ **FLOATING
C1563 tdc0.o_result\[127\] VGND 4.07f $ **FLOATING
C1564 tdc0.w_dly_sig_n\[128\] VGND 1.43f $ **FLOATING
C1565 _047_ VGND 5.9f $ **FLOATING
C1566 tdc0.o_result\[24\] VGND 5.5f $ **FLOATING
C1567 a_14917_17455# VGND 0.23f $ **FLOATING
C1568 tdc0.w_dly_sig_n\[25\] VGND 2.64f $ **FLOATING
C1569 a_12877_17833# VGND 0.23f $ **FLOATING
C1570 a_11057_17455# VGND 0.206f $ **FLOATING
C1571 a_9953_17455# VGND 0.206f $ **FLOATING
C1572 tdc0.o_result\[20\] VGND 4.89f $ **FLOATING
C1573 _053_ VGND 3.25f $ **FLOATING
C1574 _032_ VGND 3.18f $ **FLOATING
C1575 tdc0.o_result\[17\] VGND 3.35f $ **FLOATING
C1576 a_8661_17455# VGND 0.23f $ **FLOATING
C1577 a_7817_17833# VGND 0.23f $ **FLOATING
C1578 a_6273_17455# VGND 0.206f $ **FLOATING
C1579 tdc0.o_result\[16\] VGND 1.28f $ **FLOATING
C1580 _088_ VGND 2.68f $ **FLOATING
C1581 a_4521_17455# VGND 0.23f $ **FLOATING
C1582 tdc0.w_dly_sig_n\[43\] VGND 2.67f $ **FLOATING
C1583 a_2773_17455# VGND 0.23f $ **FLOATING
C1584 tdc0.w_dly_sig_n\[46\] VGND 2.36f $ **FLOATING
C1585 tdc0.w_dly_sig\[48\] VGND 3.24f $ **FLOATING
C1586 a_17703_17833# VGND 0.581f $ **FLOATING
C1587 a_17774_17732# VGND 0.626f $ **FLOATING
C1588 a_17574_17577# VGND 1.43f $ **FLOATING
C1589 a_17567_17673# VGND 1.81f $ **FLOATING
C1590 a_17283_17687# VGND 0.609f $ **FLOATING
C1591 a_17187_17687# VGND 0.817f $ **FLOATING
C1592 tdc0.w_dly_sig\[128\] VGND 3.06f $ **FLOATING
C1593 _007_ VGND 12.8f $ **FLOATING
C1594 a_16155_17687# VGND 0.804f $ **FLOATING
C1595 a_15427_17455# VGND 0.609f $ **FLOATING
C1596 a_15595_17429# VGND 0.817f $ **FLOATING
C1597 a_15002_17455# VGND 0.626f $ **FLOATING
C1598 a_15170_17429# VGND 0.581f $ **FLOATING
C1599 a_14729_17461# VGND 1.43f $ **FLOATING
C1600 a_14563_17461# VGND 1.81f $ **FLOATING
C1601 tdc0.w_dly_sig_n\[23\] VGND 2.29f $ **FLOATING
C1602 a_12459_17833# VGND 0.581f $ **FLOATING
C1603 a_12530_17732# VGND 0.626f $ **FLOATING
C1604 a_12330_17577# VGND 1.43f $ **FLOATING
C1605 a_12323_17673# VGND 1.81f $ **FLOATING
C1606 a_12039_17687# VGND 0.609f $ **FLOATING
C1607 a_11943_17687# VGND 0.817f $ **FLOATING
C1608 a_10975_17455# VGND 0.804f $ **FLOATING
C1609 tdc0.o_result\[47\] VGND 4.64f $ **FLOATING
C1610 tdc0.o_result\[45\] VGND 3.47f $ **FLOATING
C1611 net9 VGND 4.48f $ **FLOATING
C1612 a_9807_17687# VGND 0.804f $ **FLOATING
C1613 a_9171_17455# VGND 0.609f $ **FLOATING
C1614 a_9339_17429# VGND 0.817f $ **FLOATING
C1615 a_8746_17455# VGND 0.626f $ **FLOATING
C1616 a_8914_17429# VGND 0.581f $ **FLOATING
C1617 a_8473_17461# VGND 1.43f $ **FLOATING
C1618 a_8307_17461# VGND 1.81f $ **FLOATING
C1619 tdc0.w_dly_sig\[17\] VGND 4.66f $ **FLOATING
C1620 a_7399_17833# VGND 0.581f $ **FLOATING
C1621 a_7470_17732# VGND 0.626f $ **FLOATING
C1622 a_7270_17577# VGND 1.43f $ **FLOATING
C1623 a_7263_17673# VGND 1.81f $ **FLOATING
C1624 a_6979_17687# VGND 0.609f $ **FLOATING
C1625 a_6883_17687# VGND 0.817f $ **FLOATING
C1626 a_6191_17455# VGND 0.804f $ **FLOATING
C1627 net10 VGND 9.63f $ **FLOATING
C1628 _029_ VGND 14.7f $ **FLOATING
C1629 tdc0.o_result\[42\] VGND 0.864f $ **FLOATING
C1630 a_5031_17455# VGND 0.609f $ **FLOATING
C1631 a_5199_17429# VGND 0.817f $ **FLOATING
C1632 a_4606_17455# VGND 0.626f $ **FLOATING
C1633 a_4774_17429# VGND 0.581f $ **FLOATING
C1634 a_4333_17461# VGND 1.43f $ **FLOATING
C1635 a_4167_17461# VGND 1.81f $ **FLOATING
C1636 tdc0.w_dly_sig\[43\] VGND 2.84f $ **FLOATING
C1637 a_3283_17455# VGND 0.609f $ **FLOATING
C1638 a_3451_17429# VGND 0.817f $ **FLOATING
C1639 a_2858_17455# VGND 0.626f $ **FLOATING
C1640 a_3026_17429# VGND 0.581f $ **FLOATING
C1641 a_2585_17461# VGND 1.43f $ **FLOATING
C1642 a_2419_17461# VGND 1.81f $ **FLOATING
C1643 tdc0.w_dly_sig_n\[44\] VGND 2.73f $ **FLOATING
C1644 tt_um_hpretl_tt06_tdc_22.HI VGND 0.415f $ **FLOATING
C1645 a_17661_17999# VGND 0.23f $ **FLOATING
C1646 tdc0.o_result\[126\] VGND 1.05f $ **FLOATING
C1647 tdc0.o_result\[22\] VGND 0.811f $ **FLOATING
C1648 a_15561_17999# VGND 0.23f $ **FLOATING
C1649 tdc0.w_dly_sig\[127\] VGND 3.78f $ **FLOATING
C1650 a_17243_17999# VGND 0.581f $ **FLOATING
C1651 a_17314_17973# VGND 0.626f $ **FLOATING
C1652 a_17107_17973# VGND 1.81f $ **FLOATING
C1653 a_17114_18273# VGND 1.43f $ **FLOATING
C1654 a_16823_17973# VGND 0.609f $ **FLOATING
C1655 a_16727_18151# VGND 0.817f $ **FLOATING
C1656 a_16071_18365# VGND 0.609f $ **FLOATING
C1657 a_16239_18267# VGND 0.817f $ **FLOATING
C1658 a_15646_18365# VGND 0.626f $ **FLOATING
C1659 a_15814_18111# VGND 0.581f $ **FLOATING
C1660 a_15373_17999# VGND 1.43f $ **FLOATING
C1661 a_15207_17999# VGND 1.81f $ **FLOATING
C1662 clknet_4_15_0_clk VGND 11.4f $ **FLOATING
C1663 clknet_4_13_0_clk VGND 7.33f $ **FLOATING
C1664 a_14717_17999# VGND 0.23f $ **FLOATING
C1665 tdc0.o_result\[23\] VGND 1.97f $ **FLOATING
C1666 tdc0.o_result\[21\] VGND 0.865f $ **FLOATING
C1667 a_9213_17999# VGND 0.23f $ **FLOATING
C1668 a_14299_17999# VGND 0.581f $ **FLOATING
C1669 a_14370_17973# VGND 0.626f $ **FLOATING
C1670 a_14163_17973# VGND 1.81f $ **FLOATING
C1671 a_14170_18273# VGND 1.43f $ **FLOATING
C1672 a_13879_17973# VGND 0.609f $ **FLOATING
C1673 a_13783_18151# VGND 0.817f $ **FLOATING
C1674 tdc0.w_dly_sig_n\[19\] VGND 1.99f $ **FLOATING
C1675 tdc0.w_dly_sig_n\[18\] VGND 2.34f $ **FLOATING
C1676 tdc0.w_dly_sig_n\[17\] VGND 2.38f $ **FLOATING
C1677 tdc0.w_dly_sig\[18\] VGND 3.83f $ **FLOATING
C1678 a_9723_18365# VGND 0.609f $ **FLOATING
C1679 a_9891_18267# VGND 0.817f $ **FLOATING
C1680 a_9298_18365# VGND 0.626f $ **FLOATING
C1681 a_9466_18111# VGND 0.581f $ **FLOATING
C1682 a_9025_17999# VGND 1.43f $ **FLOATING
C1683 a_8859_17999# VGND 1.81f $ **FLOATING
C1684 clknet_4_7_0_clk VGND 8.9f $ **FLOATING
C1685 a_7173_17999# VGND 0.23f $ **FLOATING
C1686 tdc0.o_result\[18\] VGND 0.911f $ **FLOATING
C1687 tdc0.o_result\[19\] VGND 1.33f $ **FLOATING
C1688 a_5073_17999# VGND 0.23f $ **FLOATING
C1689 tdc0.w_dly_sig\[19\] VGND 4.56f $ **FLOATING
C1690 a_6755_17999# VGND 0.581f $ **FLOATING
C1691 a_6826_17973# VGND 0.626f $ **FLOATING
C1692 a_6619_17973# VGND 1.81f $ **FLOATING
C1693 a_6626_18273# VGND 1.43f $ **FLOATING
C1694 a_6335_17973# VGND 0.609f $ **FLOATING
C1695 a_6239_18151# VGND 0.817f $ **FLOATING
C1696 a_5583_18365# VGND 0.609f $ **FLOATING
C1697 a_5751_18267# VGND 0.817f $ **FLOATING
C1698 a_5158_18365# VGND 0.626f $ **FLOATING
C1699 a_5326_18111# VGND 0.581f $ **FLOATING
C1700 a_4885_17999# VGND 1.43f $ **FLOATING
C1701 a_4719_17999# VGND 1.81f $ **FLOATING
C1702 tdc0.o_result\[43\] VGND 1.89f $ **FLOATING
C1703 a_3601_17999# VGND 0.23f $ **FLOATING
C1704 a_4111_18365# VGND 0.609f $ **FLOATING
C1705 a_4279_18267# VGND 0.817f $ **FLOATING
C1706 a_3686_18365# VGND 0.626f $ **FLOATING
C1707 a_3854_18111# VGND 0.581f $ **FLOATING
C1708 a_3413_17999# VGND 1.43f $ **FLOATING
C1709 a_3247_17999# VGND 1.81f $ **FLOATING
C1710 clknet_4_5_0_clk VGND 13.5f $ **FLOATING
C1711 tdc0.w_dly_sig\[46\] VGND 3.04f $ **FLOATING
C1712 tt_um_hpretl_tt06_tdc_24.HI VGND 0.415f $ **FLOATING
C1713 tdc0.w_dly_sig\[44\] VGND 3.69f $ **FLOATING
C1714 tdc0.w_dly_sig_n\[45\] VGND 2.87f $ **FLOATING
C1715 tt_um_hpretl_tt06_tdc_16.HI VGND 0.415f $ **FLOATING
C1716 tt_um_hpretl_tt06_tdc_25.HI VGND 0.415f $ **FLOATING
C1717 tdc0.w_dly_sig\[25\] VGND 3.6f $ **FLOATING
C1718 tdc0.w_dly_sig\[24\] VGND 4.08f $ **FLOATING
C1719 tdc0.w_dly_sig\[23\] VGND 4.6f $ **FLOATING
C1720 tdc0.w_dly_sig_n\[24\] VGND 2.76f $ **FLOATING
C1721 tdc0.w_dly_sig_n\[22\] VGND 2.59f $ **FLOATING
C1722 tdc0.w_dly_sig\[22\] VGND 4.2f $ **FLOATING
C1723 tdc0.w_dly_sig\[21\] VGND 3.27f $ **FLOATING
C1724 tdc0.w_dly_sig_n\[21\] VGND 2.25f $ **FLOATING
C1725 tdc0.w_dly_sig_n\[20\] VGND 2.49f $ **FLOATING
C1726 tdc0.w_dly_sig\[20\] VGND 5.79f $ **FLOATING
C1727 tt_um_hpretl_tt06_tdc_26.HI VGND 0.415f $ **FLOATING
C1728 tt_um_hpretl_tt06_tdc_13.HI VGND 0.415f $ **FLOATING
C1729 tt_um_hpretl_tt06_tdc_20.HI VGND 0.415f $ **FLOATING
.ends
