magic
tech sky130A
magscale 1 2
timestamp 1710673697
<< viali >>
rect 20637 17697 20671 17731
rect 20729 17493 20763 17527
rect 12817 17289 12851 17323
rect 20269 17289 20303 17323
rect 21373 17289 21407 17323
rect 21925 17289 21959 17323
rect 11621 17221 11655 17255
rect 13093 17221 13127 17255
rect 21097 17221 21131 17255
rect 12173 17153 12207 17187
rect 11069 17085 11103 17119
rect 11161 17095 11195 17129
rect 11437 17085 11471 17119
rect 11713 17085 11747 17119
rect 11805 17085 11839 17119
rect 12081 17085 12115 17119
rect 12633 17085 12667 17119
rect 12725 17085 12759 17119
rect 13001 17085 13035 17119
rect 13737 17085 13771 17119
rect 13829 17085 13863 17119
rect 14841 17085 14875 17119
rect 20361 17085 20395 17119
rect 20637 17087 20671 17121
rect 20729 17085 20763 17119
rect 21005 17085 21039 17119
rect 21465 17085 21499 17119
rect 21741 17085 21775 17119
rect 22017 17085 22051 17119
rect 22109 17085 22143 17119
rect 22385 17085 22419 17119
rect 22477 17085 22511 17119
rect 22661 17085 22695 17119
rect 23121 17085 23155 17119
rect 13645 17017 13679 17051
rect 20545 17017 20579 17051
rect 11345 16949 11379 16983
rect 11897 16949 11931 16983
rect 12541 16949 12575 16983
rect 13921 16949 13955 16983
rect 14933 16949 14967 16983
rect 20821 16949 20855 16983
rect 21649 16949 21683 16983
rect 22201 16949 22235 16983
rect 22753 16949 22787 16983
rect 23029 16949 23063 16983
rect 10701 16745 10735 16779
rect 13829 16745 13863 16779
rect 22477 16745 22511 16779
rect 22753 16745 22787 16779
rect 23029 16745 23063 16779
rect 23581 16745 23615 16779
rect 10425 16677 10459 16711
rect 11897 16677 11931 16711
rect 15025 16677 15059 16711
rect 15853 16677 15887 16711
rect 18889 16677 18923 16711
rect 20637 16677 20671 16711
rect 22201 16677 22235 16711
rect 23305 16677 23339 16711
rect 10149 16609 10183 16643
rect 10517 16609 10551 16643
rect 10609 16609 10643 16643
rect 10977 16609 11011 16643
rect 11069 16609 11103 16643
rect 11253 16609 11287 16643
rect 11345 16609 11379 16643
rect 11529 16609 11563 16643
rect 11989 16609 12023 16643
rect 12265 16609 12299 16643
rect 12357 16609 12391 16643
rect 12725 16609 12759 16643
rect 13185 16609 13219 16643
rect 13461 16609 13495 16643
rect 13737 16609 13771 16643
rect 14013 16609 14047 16643
rect 14105 16609 14139 16643
rect 14289 16609 14323 16643
rect 14749 16609 14783 16643
rect 14841 16609 14875 16643
rect 14933 16609 14967 16643
rect 15209 16609 15243 16643
rect 15669 16609 15703 16643
rect 15945 16609 15979 16643
rect 16221 16609 16255 16643
rect 16313 16609 16347 16643
rect 18981 16609 19015 16643
rect 19257 16609 19291 16643
rect 19349 16609 19383 16643
rect 19625 16609 19659 16643
rect 20085 16609 20119 16643
rect 20453 16609 20487 16643
rect 20729 16609 20763 16643
rect 21005 16609 21039 16643
rect 21465 16609 21499 16643
rect 21557 16609 21591 16643
rect 21925 16609 21959 16643
rect 22017 16609 22051 16643
rect 22293 16609 22327 16643
rect 22569 16609 22603 16643
rect 22845 16609 22879 16643
rect 23121 16609 23155 16643
rect 23213 16609 23247 16643
rect 23673 16609 23707 16643
rect 10057 16541 10091 16575
rect 20361 16541 20395 16575
rect 11621 16473 11655 16507
rect 14381 16473 14415 16507
rect 15577 16473 15611 16507
rect 19165 16473 19199 16507
rect 12173 16405 12207 16439
rect 12449 16405 12483 16439
rect 12817 16405 12851 16439
rect 13093 16405 13127 16439
rect 13369 16405 13403 16439
rect 15301 16405 15335 16439
rect 19441 16405 19475 16439
rect 19717 16405 19751 16439
rect 19993 16405 20027 16439
rect 20913 16405 20947 16439
rect 21373 16405 21407 16439
rect 21649 16405 21683 16439
rect 10977 16201 11011 16235
rect 11805 16201 11839 16235
rect 13001 16201 13035 16235
rect 14013 16201 14047 16235
rect 15117 16201 15151 16235
rect 19901 16201 19935 16235
rect 21005 16201 21039 16235
rect 21281 16201 21315 16235
rect 22109 16201 22143 16235
rect 23213 16201 23247 16235
rect 24501 16201 24535 16235
rect 10425 16133 10459 16167
rect 18153 16133 18187 16167
rect 23489 16065 23523 16099
rect 9689 15997 9723 16031
rect 9781 15997 9815 16031
rect 10241 15997 10275 16031
rect 10341 15991 10375 16025
rect 10609 15997 10643 16031
rect 10885 15997 10919 16031
rect 11161 15997 11195 16031
rect 11621 15997 11655 16031
rect 11713 15997 11747 16031
rect 11989 15997 12023 16031
rect 12081 15997 12115 16031
rect 12265 15997 12299 16031
rect 12633 15997 12667 16031
rect 12817 15997 12851 16031
rect 13093 15997 13127 16031
rect 13369 15997 13403 16031
rect 13645 15997 13679 16031
rect 13737 15997 13771 16031
rect 13921 15997 13955 16031
rect 14381 15997 14415 16031
rect 14473 15997 14507 16031
rect 14565 15997 14599 16031
rect 14749 15997 14783 16031
rect 15209 15997 15243 16031
rect 15577 15997 15611 16031
rect 15761 15997 15795 16031
rect 15945 15997 15979 16031
rect 16221 15997 16255 16031
rect 16313 15997 16347 16031
rect 16581 15997 16615 16031
rect 17233 15997 17267 16031
rect 17417 15997 17451 16031
rect 17509 15997 17543 16031
rect 18245 15999 18279 16033
rect 18337 15997 18371 16031
rect 18889 15997 18923 16031
rect 18981 15997 19015 16031
rect 19441 15997 19475 16031
rect 19717 15997 19751 16031
rect 19809 15997 19843 16031
rect 19993 15997 20027 16031
rect 20269 15997 20303 16031
rect 20545 15997 20579 16031
rect 20637 15997 20671 16031
rect 20913 15997 20947 16031
rect 21097 15997 21131 16031
rect 21373 15997 21407 16031
rect 21465 15997 21499 16031
rect 21925 15997 21959 16031
rect 22017 15997 22051 16031
rect 22201 15997 22235 16031
rect 22293 15997 22327 16031
rect 22569 15997 22603 16031
rect 23029 15997 23063 16031
rect 23305 15997 23339 16031
rect 23581 15997 23615 16031
rect 23857 15997 23891 16031
rect 24133 15997 24167 16031
rect 24593 15997 24627 16031
rect 9597 15929 9631 15963
rect 13277 15929 13311 15963
rect 14289 15929 14323 15963
rect 16405 15929 16439 15963
rect 18797 15929 18831 15963
rect 19625 15929 19659 15963
rect 20453 15929 20487 15963
rect 23949 15929 23983 15963
rect 9873 15861 9907 15895
rect 10149 15861 10183 15895
rect 10701 15861 10735 15895
rect 11253 15861 11287 15895
rect 11529 15861 11563 15895
rect 12357 15861 12391 15895
rect 12725 15861 12759 15895
rect 14841 15861 14875 15895
rect 15485 15861 15519 15895
rect 15945 15861 15979 15895
rect 16129 15861 16163 15895
rect 16681 15861 16715 15895
rect 17141 15861 17175 15895
rect 18429 15861 18463 15895
rect 19073 15861 19107 15895
rect 19349 15861 19383 15895
rect 20177 15861 20211 15895
rect 20729 15861 20763 15895
rect 21557 15861 21591 15895
rect 21833 15861 21867 15895
rect 22385 15861 22419 15895
rect 22661 15861 22695 15895
rect 22937 15861 22971 15895
rect 24225 15861 24259 15895
rect 8769 15657 8803 15691
rect 9873 15657 9907 15691
rect 11713 15657 11747 15691
rect 13553 15657 13587 15691
rect 13737 15657 13771 15691
rect 14105 15657 14139 15691
rect 15117 15657 15151 15691
rect 15301 15657 15335 15691
rect 16773 15657 16807 15691
rect 19165 15657 19199 15691
rect 20361 15657 20395 15691
rect 23029 15657 23063 15691
rect 24409 15657 24443 15691
rect 24961 15657 24995 15691
rect 9597 15589 9631 15623
rect 12817 15589 12851 15623
rect 19809 15589 19843 15623
rect 24133 15589 24167 15623
rect 8677 15521 8711 15555
rect 8953 15521 8987 15555
rect 9413 15521 9447 15555
rect 9505 15521 9539 15555
rect 9781 15521 9815 15555
rect 10057 15521 10091 15555
rect 10149 15521 10183 15555
rect 10333 15521 10367 15555
rect 10517 15521 10551 15555
rect 10793 15521 10827 15555
rect 11253 15521 11287 15555
rect 11345 15521 11379 15555
rect 11437 15521 11471 15555
rect 11805 15521 11839 15555
rect 12081 15521 12115 15555
rect 12173 15521 12207 15555
rect 12449 15521 12483 15555
rect 12725 15521 12759 15555
rect 13185 15521 13219 15555
rect 13461 15521 13495 15555
rect 13737 15521 13771 15555
rect 13921 15521 13955 15555
rect 14197 15521 14231 15555
rect 14381 15521 14415 15555
rect 14473 15521 14507 15555
rect 14565 15521 14599 15555
rect 15025 15521 15059 15555
rect 15301 15521 15335 15555
rect 15485 15521 15519 15555
rect 15577 15521 15611 15555
rect 16313 15521 16347 15555
rect 16405 15521 16439 15555
rect 16681 15519 16715 15553
rect 16957 15521 16991 15555
rect 17417 15521 17451 15555
rect 17601 15521 17635 15555
rect 17693 15521 17727 15555
rect 17785 15521 17819 15555
rect 18245 15521 18279 15555
rect 18337 15521 18371 15555
rect 18797 15521 18831 15555
rect 18981 15521 19015 15555
rect 19073 15521 19107 15555
rect 19165 15521 19199 15555
rect 19349 15521 19383 15555
rect 19625 15521 19659 15555
rect 19717 15521 19751 15555
rect 19993 15521 20027 15555
rect 20453 15521 20487 15555
rect 20545 15521 20579 15555
rect 20821 15521 20855 15555
rect 21281 15521 21315 15555
rect 21557 15521 21591 15555
rect 21925 15521 21959 15555
rect 22017 15521 22051 15555
rect 22293 15521 22327 15555
rect 22385 15521 22419 15555
rect 22569 15521 22603 15555
rect 22661 15521 22695 15555
rect 23121 15521 23155 15555
rect 23397 15521 23431 15555
rect 23581 15521 23615 15555
rect 23673 15521 23707 15555
rect 23949 15521 23983 15555
rect 24225 15521 24259 15555
rect 24317 15521 24351 15555
rect 24593 15521 24627 15555
rect 24869 15521 24903 15555
rect 10425 15453 10459 15487
rect 11161 15453 11195 15487
rect 11989 15453 12023 15487
rect 15669 15453 15703 15487
rect 17049 15453 17083 15487
rect 17877 15453 17911 15487
rect 19533 15453 19567 15487
rect 24685 15453 24719 15487
rect 9321 15385 9355 15419
rect 10701 15385 10735 15419
rect 16221 15385 16255 15419
rect 18429 15385 18463 15419
rect 20085 15385 20119 15419
rect 22201 15385 22235 15419
rect 22477 15385 22511 15419
rect 9045 15317 9079 15351
rect 12265 15317 12299 15351
rect 12541 15317 12575 15351
rect 13277 15317 13311 15351
rect 14657 15317 14691 15351
rect 16497 15317 16531 15351
rect 17325 15317 17359 15351
rect 18153 15317 18187 15351
rect 18705 15317 18739 15351
rect 20637 15317 20671 15351
rect 20913 15317 20947 15351
rect 21373 15317 21407 15351
rect 21649 15317 21683 15351
rect 22753 15317 22787 15351
rect 23305 15317 23339 15351
rect 23857 15317 23891 15351
rect 9045 15113 9079 15147
rect 10149 15113 10183 15147
rect 10701 15113 10735 15147
rect 13645 15113 13679 15147
rect 16589 15113 16623 15147
rect 18429 15113 18463 15147
rect 20085 15113 20119 15147
rect 23489 15113 23523 15147
rect 23949 15113 23983 15147
rect 12633 15045 12667 15079
rect 18153 15045 18187 15079
rect 23213 15045 23247 15079
rect 24777 15045 24811 15079
rect 25053 15045 25087 15079
rect 25329 15045 25363 15079
rect 9597 14977 9631 15011
rect 10885 14977 10919 15011
rect 12909 14977 12943 15011
rect 18705 14977 18739 15011
rect 21741 14977 21775 15011
rect 21833 14977 21867 15011
rect 7941 14909 7975 14943
rect 8033 14909 8067 14943
rect 8401 14909 8435 14943
rect 8677 14909 8711 14943
rect 8861 14909 8895 14943
rect 9137 14909 9171 14943
rect 9413 14909 9447 14943
rect 9689 14909 9723 14943
rect 9965 14909 9999 14943
rect 10057 14909 10091 14943
rect 10517 14909 10551 14943
rect 10793 14909 10827 14943
rect 12541 14909 12575 14943
rect 13001 14909 13035 14943
rect 13093 14909 13127 14943
rect 15025 14909 15059 14943
rect 15209 14909 15243 14943
rect 16773 14909 16807 14943
rect 18337 14909 18371 14943
rect 18972 14909 19006 14943
rect 21485 14909 21519 14943
rect 23397 14909 23431 14943
rect 23581 14909 23615 14943
rect 23857 14909 23891 14943
rect 24317 14909 24351 14943
rect 24501 14909 24535 14943
rect 24593 14909 24627 14943
rect 24685 14909 24719 14943
rect 24961 14909 24995 14943
rect 25237 14909 25271 14943
rect 25513 14909 25547 14943
rect 7849 14841 7883 14875
rect 8125 14841 8159 14875
rect 9873 14841 9907 14875
rect 11130 14841 11164 14875
rect 14780 14841 14814 14875
rect 15476 14841 15510 14875
rect 17040 14841 17074 14875
rect 22100 14841 22134 14875
rect 8493 14773 8527 14807
rect 8677 14773 8711 14807
rect 9321 14773 9355 14807
rect 10425 14773 10459 14807
rect 12265 14773 12299 14807
rect 13185 14773 13219 14807
rect 20361 14773 20395 14807
rect 24225 14773 24259 14807
rect 25605 14773 25639 14807
rect 7941 14569 7975 14603
rect 9045 14569 9079 14603
rect 10609 14569 10643 14603
rect 13369 14569 13403 14603
rect 15761 14569 15795 14603
rect 16773 14569 16807 14603
rect 17693 14569 17727 14603
rect 18981 14569 19015 14603
rect 24041 14569 24075 14603
rect 25421 14569 25455 14603
rect 25697 14569 25731 14603
rect 7665 14501 7699 14535
rect 11253 14501 11287 14535
rect 13001 14501 13035 14535
rect 19809 14501 19843 14535
rect 21925 14501 21959 14535
rect 22201 14501 22235 14535
rect 22652 14501 22686 14535
rect 7481 14433 7515 14467
rect 7757 14433 7791 14467
rect 7849 14433 7883 14467
rect 8033 14433 8067 14467
rect 8125 14433 8159 14467
rect 8585 14433 8619 14467
rect 8677 14433 8711 14467
rect 9137 14433 9171 14467
rect 9485 14433 9519 14467
rect 11161 14433 11195 14467
rect 13461 14433 13495 14467
rect 13737 14433 13771 14467
rect 13829 14433 13863 14467
rect 14289 14433 14323 14467
rect 14648 14433 14682 14467
rect 16313 14433 16347 14467
rect 16405 14433 16439 14467
rect 16865 14433 16899 14467
rect 16957 14433 16991 14467
rect 17233 14433 17267 14467
rect 17509 14433 17543 14467
rect 17693 14433 17727 14467
rect 17969 14433 18003 14467
rect 18061 14433 18095 14467
rect 18521 14433 18555 14467
rect 18797 14433 18831 14467
rect 18889 14433 18923 14467
rect 19165 14433 19199 14467
rect 19349 14433 19383 14467
rect 19441 14433 19475 14467
rect 19901 14433 19935 14467
rect 19993 14433 20027 14467
rect 20453 14433 20487 14467
rect 20729 14423 20763 14457
rect 21005 14433 21039 14467
rect 21465 14433 21499 14467
rect 21557 14433 21591 14467
rect 22017 14433 22051 14467
rect 22293 14433 22327 14467
rect 22385 14433 22419 14467
rect 24133 14433 24167 14467
rect 24225 14433 24259 14467
rect 24685 14433 24719 14467
rect 24961 14431 24995 14465
rect 25061 14433 25095 14467
rect 25513 14433 25547 14467
rect 25789 14433 25823 14467
rect 25881 14433 25915 14467
rect 9229 14365 9263 14399
rect 13645 14365 13679 14399
rect 14381 14365 14415 14399
rect 16497 14365 16531 14399
rect 17877 14365 17911 14399
rect 25973 14365 26007 14399
rect 7389 14297 7423 14331
rect 14197 14297 14231 14331
rect 17049 14297 17083 14331
rect 24317 14297 24351 14331
rect 8217 14229 8251 14263
rect 8493 14229 8527 14263
rect 8769 14229 8803 14263
rect 11069 14229 11103 14263
rect 13921 14229 13955 14263
rect 16221 14229 16255 14263
rect 17325 14229 17359 14263
rect 18153 14229 18187 14263
rect 18429 14229 18463 14263
rect 18705 14229 18739 14263
rect 19257 14229 19291 14263
rect 19533 14229 19567 14263
rect 20085 14229 20119 14263
rect 20361 14229 20395 14263
rect 20637 14229 20671 14263
rect 20913 14229 20947 14263
rect 21373 14229 21407 14263
rect 21649 14229 21683 14263
rect 23765 14229 23799 14263
rect 24593 14229 24627 14263
rect 24869 14229 24903 14263
rect 25145 14229 25179 14263
rect 7021 14025 7055 14059
rect 8125 14025 8159 14059
rect 10057 14025 10091 14059
rect 12173 14025 12207 14059
rect 12449 14025 12483 14059
rect 17877 14025 17911 14059
rect 18153 14025 18187 14059
rect 20637 14025 20671 14059
rect 20913 14025 20947 14059
rect 21465 14025 21499 14059
rect 25053 14025 25087 14059
rect 25329 14025 25363 14059
rect 25605 14025 25639 14059
rect 26157 14025 26191 14059
rect 26433 14025 26467 14059
rect 7297 13957 7331 13991
rect 10517 13957 10551 13991
rect 11345 13957 11379 13991
rect 11621 13957 11655 13991
rect 13001 13957 13035 13991
rect 13277 13957 13311 13991
rect 13829 13957 13863 13991
rect 15393 13957 15427 13991
rect 19993 13957 20027 13991
rect 21189 13957 21223 13991
rect 23581 13957 23615 13991
rect 24225 13957 24259 13991
rect 25881 13957 25915 13991
rect 7573 13889 7607 13923
rect 8677 13889 8711 13923
rect 12725 13889 12759 13923
rect 16037 13889 16071 13923
rect 16589 13889 16623 13923
rect 17601 13889 17635 13923
rect 18429 13889 18463 13923
rect 7113 13821 7147 13855
rect 7205 13821 7239 13855
rect 7397 13815 7431 13849
rect 7665 13821 7699 13855
rect 7941 13821 7975 13855
rect 8033 13821 8067 13855
rect 8401 13821 8435 13855
rect 10609 13821 10643 13855
rect 10701 13821 10735 13855
rect 10793 13821 10827 13855
rect 10977 13821 11011 13855
rect 11437 13821 11471 13855
rect 11713 13821 11747 13855
rect 11989 13821 12023 13855
rect 12081 13821 12115 13855
rect 12541 13821 12575 13855
rect 12817 13821 12851 13855
rect 13093 13821 13127 13855
rect 13369 13821 13403 13855
rect 15209 13821 15243 13855
rect 15485 13821 15519 13855
rect 15853 13821 15887 13855
rect 15945 13821 15979 13855
rect 16221 13821 16255 13855
rect 16313 13821 16347 13855
rect 16497 13821 16531 13855
rect 17141 13821 17175 13855
rect 17233 13821 17267 13855
rect 17693 13821 17727 13855
rect 17969 13821 18003 13855
rect 18245 13821 18279 13855
rect 18337 13821 18371 13855
rect 18705 13821 18739 13855
rect 20729 13821 20763 13855
rect 20821 13821 20855 13855
rect 21281 13821 21315 13855
rect 21373 13821 21407 13855
rect 21833 13821 21867 13855
rect 21925 13821 21959 13855
rect 22201 13821 22235 13855
rect 22468 13821 22502 13855
rect 24041 13821 24075 13855
rect 24133 13821 24167 13855
rect 24593 13821 24627 13855
rect 24869 13821 24903 13855
rect 25145 13821 25179 13855
rect 25421 13821 25455 13855
rect 25697 13821 25731 13855
rect 25789 13821 25823 13855
rect 26065 13821 26099 13855
rect 26341 13821 26375 13855
rect 26617 13821 26651 13855
rect 8922 13753 8956 13787
rect 11069 13753 11103 13787
rect 14942 13753 14976 13787
rect 23949 13753 23983 13787
rect 7849 13685 7883 13719
rect 8493 13685 8527 13719
rect 11897 13685 11931 13719
rect 15761 13685 15795 13719
rect 17049 13685 17083 13719
rect 17325 13685 17359 13719
rect 21741 13685 21775 13719
rect 22017 13685 22051 13719
rect 24501 13685 24535 13719
rect 24777 13685 24811 13719
rect 26709 13685 26743 13719
rect 9597 13481 9631 13515
rect 10149 13481 10183 13515
rect 10425 13481 10459 13515
rect 13369 13481 13403 13515
rect 13737 13481 13771 13515
rect 14013 13481 14047 13515
rect 17509 13481 17543 13515
rect 19073 13481 19107 13515
rect 20637 13481 20671 13515
rect 21741 13481 21775 13515
rect 25329 13481 25363 13515
rect 25697 13481 25731 13515
rect 25973 13481 26007 13515
rect 11253 13413 11287 13447
rect 12256 13413 12290 13447
rect 15945 13413 15979 13447
rect 19524 13413 19558 13447
rect 7481 13345 7515 13379
rect 7573 13345 7607 13379
rect 7757 13345 7791 13379
rect 8033 13345 8067 13379
rect 8125 13345 8159 13379
rect 8217 13345 8251 13379
rect 8401 13345 8435 13379
rect 8861 13345 8895 13379
rect 9137 13335 9171 13369
rect 9229 13345 9263 13379
rect 9505 13345 9539 13379
rect 9781 13345 9815 13379
rect 9965 13345 9999 13379
rect 10057 13345 10091 13379
rect 10333 13345 10367 13379
rect 10609 13345 10643 13379
rect 11161 13345 11195 13379
rect 11621 13345 11655 13379
rect 11713 13345 11747 13379
rect 13829 13345 13863 13379
rect 13921 13345 13955 13379
rect 16385 13345 16419 13379
rect 17693 13345 17727 13379
rect 17960 13345 17994 13379
rect 19257 13345 19291 13379
rect 21005 13345 21039 13379
rect 21557 13345 21591 13379
rect 21649 13345 21683 13379
rect 22109 13345 22143 13379
rect 22468 13345 22502 13379
rect 23765 13345 23799 13379
rect 24032 13345 24066 13379
rect 25329 13345 25363 13379
rect 25513 13345 25547 13379
rect 25605 13345 25639 13379
rect 25881 13345 25915 13379
rect 26433 13345 26467 13379
rect 7665 13277 7699 13311
rect 9321 13277 9355 13311
rect 11989 13277 12023 13311
rect 14197 13277 14231 13311
rect 16129 13277 16163 13311
rect 22201 13277 22235 13311
rect 10701 13209 10735 13243
rect 22017 13209 22051 13243
rect 7389 13141 7423 13175
rect 7941 13141 7975 13175
rect 8493 13141 8527 13175
rect 8769 13141 8803 13175
rect 9045 13141 9079 13175
rect 9873 13141 9907 13175
rect 11529 13141 11563 13175
rect 11805 13141 11839 13175
rect 20913 13141 20947 13175
rect 21465 13141 21499 13175
rect 23581 13141 23615 13175
rect 25145 13141 25179 13175
rect 26525 13141 26559 13175
rect 7573 12937 7607 12971
rect 8953 12937 8987 12971
rect 10793 12937 10827 12971
rect 13001 12937 13035 12971
rect 15025 12937 15059 12971
rect 18429 12937 18463 12971
rect 20085 12937 20119 12971
rect 24501 12937 24535 12971
rect 24777 12937 24811 12971
rect 7895 12869 7929 12903
rect 10517 12869 10551 12903
rect 16497 12869 16531 12903
rect 24225 12801 24259 12835
rect 25605 12801 25639 12835
rect 26157 12801 26191 12835
rect 26433 12801 26467 12835
rect 7665 12733 7699 12767
rect 7824 12727 7858 12761
rect 8033 12733 8067 12767
rect 8217 12733 8251 12767
rect 8585 12733 8619 12767
rect 10333 12733 10367 12767
rect 10425 12733 10459 12767
rect 10885 12733 10919 12767
rect 12725 12733 12759 12767
rect 12909 12733 12943 12767
rect 13185 12733 13219 12767
rect 13645 12733 13679 12767
rect 15209 12733 15243 12767
rect 17049 12733 17083 12767
rect 18705 12733 18739 12767
rect 20453 12733 20487 12767
rect 20637 12733 20671 12767
rect 20729 12733 20763 12767
rect 21005 12733 21039 12767
rect 21281 12733 21315 12767
rect 21557 12733 21591 12767
rect 21833 12733 21867 12767
rect 23857 12733 23891 12767
rect 23949 12733 23983 12767
rect 24133 12733 24167 12767
rect 24317 12733 24351 12767
rect 24409 12733 24443 12767
rect 24685 12733 24719 12767
rect 24869 12733 24903 12767
rect 24961 12733 24995 12767
rect 25421 12733 25455 12767
rect 25697 12733 25731 12767
rect 25881 12733 25915 12767
rect 25973 12733 26007 12767
rect 26249 12733 26283 12767
rect 26341 12733 26375 12767
rect 26617 12733 26651 12767
rect 10066 12665 10100 12699
rect 10977 12665 11011 12699
rect 13890 12665 13924 12699
rect 17294 12665 17328 12699
rect 18972 12665 19006 12699
rect 20361 12665 20395 12699
rect 21741 12665 21775 12699
rect 21925 12665 21959 12699
rect 23673 12665 23707 12699
rect 25329 12665 25363 12699
rect 26709 12665 26743 12699
rect 8217 12597 8251 12631
rect 8677 12597 8711 12631
rect 13277 12597 13311 12631
rect 20913 12597 20947 12631
rect 21189 12597 21223 12631
rect 21465 12597 21499 12631
rect 25053 12597 25087 12631
rect 8493 12393 8527 12427
rect 8769 12393 8803 12427
rect 9275 12393 9309 12427
rect 9597 12393 9631 12427
rect 10241 12393 10275 12427
rect 11161 12393 11195 12427
rect 11437 12393 11471 12427
rect 11989 12393 12023 12427
rect 12541 12393 12575 12427
rect 12817 12393 12851 12427
rect 15025 12393 15059 12427
rect 15209 12393 15243 12427
rect 15577 12393 15611 12427
rect 16773 12393 16807 12427
rect 18889 12393 18923 12427
rect 20913 12393 20947 12427
rect 24501 12393 24535 12427
rect 8217 12325 8251 12359
rect 21281 12325 21315 12359
rect 23388 12325 23422 12359
rect 25881 12325 25915 12359
rect 26157 12325 26191 12359
rect 7849 12257 7883 12291
rect 8125 12257 8159 12291
rect 8585 12257 8619 12291
rect 8861 12257 8895 12291
rect 9137 12257 9171 12291
rect 9378 12257 9412 12291
rect 9689 12257 9723 12291
rect 9781 12257 9815 12291
rect 9873 12257 9907 12291
rect 10057 12257 10091 12291
rect 10241 12257 10275 12291
rect 10333 12257 10367 12291
rect 10425 12257 10459 12291
rect 10609 12257 10643 12291
rect 11069 12257 11103 12291
rect 11529 12257 11563 12291
rect 11621 12257 11655 12291
rect 11897 12257 11931 12291
rect 12081 12257 12115 12291
rect 12357 12257 12391 12291
rect 12449 12257 12483 12291
rect 12717 12255 12751 12289
rect 13001 12257 13035 12291
rect 13277 12257 13311 12291
rect 13461 12257 13495 12291
rect 13553 12257 13587 12291
rect 13645 12257 13679 12291
rect 14013 12257 14047 12291
rect 14289 12247 14323 12281
rect 14381 12257 14415 12291
rect 14473 12257 14507 12291
rect 14657 12257 14691 12291
rect 14933 12257 14967 12291
rect 15209 12257 15243 12291
rect 15393 12257 15427 12291
rect 15669 12257 15703 12291
rect 15761 12257 15795 12291
rect 15853 12257 15887 12291
rect 16129 12257 16163 12291
rect 16589 12257 16623 12291
rect 16681 12257 16715 12291
rect 17141 12257 17175 12291
rect 17233 12257 17267 12291
rect 17601 12257 17635 12291
rect 19441 12257 19475 12291
rect 19717 12257 19751 12291
rect 20177 12257 20211 12291
rect 20637 12257 20671 12291
rect 20729 12257 20763 12291
rect 20913 12257 20947 12291
rect 24685 12257 24719 12291
rect 24777 12257 24811 12291
rect 25145 12257 25179 12291
rect 25329 12257 25363 12291
rect 25421 12257 25455 12291
rect 25513 12257 25547 12291
rect 25973 12257 26007 12291
rect 26249 12257 26283 12291
rect 23121 12189 23155 12223
rect 12265 12121 12299 12155
rect 14197 12121 14231 12155
rect 17049 12121 17083 12155
rect 19809 12121 19843 12155
rect 25053 12121 25087 12155
rect 7941 12053 7975 12087
rect 9045 12053 9079 12087
rect 10701 12053 10735 12087
rect 11713 12053 11747 12087
rect 13093 12053 13127 12087
rect 13369 12053 13403 12087
rect 13921 12053 13955 12087
rect 14749 12053 14783 12087
rect 16221 12053 16255 12087
rect 16497 12053 16531 12087
rect 17325 12053 17359 12087
rect 19533 12053 19567 12087
rect 20085 12053 20119 12087
rect 20545 12053 20579 12087
rect 22569 12053 22603 12087
rect 25605 12053 25639 12087
rect 7619 11849 7653 11883
rect 11437 11849 11471 11883
rect 11713 11849 11747 11883
rect 13737 11849 13771 11883
rect 14013 11849 14047 11883
rect 14289 11849 14323 11883
rect 15393 11849 15427 11883
rect 16313 11849 16347 11883
rect 18429 11849 18463 11883
rect 20269 11849 20303 11883
rect 20545 11849 20579 11883
rect 20821 11849 20855 11883
rect 21097 11849 21131 11883
rect 24501 11849 24535 11883
rect 24777 11849 24811 11883
rect 8447 11781 8481 11815
rect 9045 11781 9079 11815
rect 14565 11781 14599 11815
rect 16589 11781 16623 11815
rect 21649 11781 21683 11815
rect 25881 11781 25915 11815
rect 8723 11713 8757 11747
rect 13093 11713 13127 11747
rect 15669 11713 15703 11747
rect 16865 11713 16899 11747
rect 18705 11713 18739 11747
rect 21925 11713 21959 11747
rect 7548 11645 7582 11679
rect 7792 11645 7826 11679
rect 8100 11645 8134 11679
rect 8518 11645 8552 11679
rect 8826 11645 8860 11679
rect 8953 11645 8987 11679
rect 9264 11653 9298 11687
rect 9689 11645 9723 11679
rect 9965 11645 9999 11679
rect 10057 11645 10091 11679
rect 13185 11645 13219 11679
rect 13277 11645 13311 11679
rect 13645 11645 13679 11679
rect 13829 11645 13863 11679
rect 13921 11645 13955 11679
rect 14197 11645 14231 11679
rect 14473 11645 14507 11679
rect 14933 11645 14967 11679
rect 15025 11645 15059 11679
rect 15485 11647 15519 11681
rect 15577 11645 15611 11679
rect 16037 11645 16071 11679
rect 16405 11645 16439 11679
rect 16681 11645 16715 11679
rect 17141 11645 17175 11679
rect 18981 11645 19015 11679
rect 20637 11645 20671 11679
rect 20913 11645 20947 11679
rect 21189 11645 21223 11679
rect 21465 11645 21499 11679
rect 21741 11645 21775 11679
rect 21833 11645 21867 11679
rect 22201 11645 22235 11679
rect 22468 11645 22502 11679
rect 24041 11655 24075 11689
rect 24317 11645 24351 11679
rect 24593 11645 24627 11679
rect 24685 11645 24719 11679
rect 24869 11645 24903 11679
rect 25145 11645 25179 11679
rect 25421 11645 25455 11679
rect 25697 11645 25731 11679
rect 25789 11645 25823 11679
rect 26065 11645 26099 11679
rect 7895 11577 7929 11611
rect 10302 11577 10336 11611
rect 12826 11577 12860 11611
rect 15945 11577 15979 11611
rect 21373 11577 21407 11611
rect 23949 11577 23983 11611
rect 25605 11577 25639 11611
rect 26157 11577 26191 11611
rect 8171 11509 8205 11543
rect 9367 11509 9401 11543
rect 9597 11509 9631 11543
rect 9873 11509 9907 11543
rect 14841 11509 14875 11543
rect 15117 11509 15151 11543
rect 23581 11509 23615 11543
rect 24225 11509 24259 11543
rect 25053 11509 25087 11543
rect 25329 11509 25363 11543
rect 11621 11305 11655 11339
rect 14565 11305 14599 11339
rect 15669 11305 15703 11339
rect 18245 11305 18279 11339
rect 19441 11305 19475 11339
rect 19717 11305 19751 11339
rect 10425 11237 10459 11271
rect 20361 11237 20395 11271
rect 21005 11237 21039 11271
rect 23305 11237 23339 11271
rect 8125 11169 8159 11203
rect 8401 11169 8435 11203
rect 8861 11169 8895 11203
rect 9137 11169 9171 11203
rect 9321 11169 9355 11203
rect 9413 11169 9447 11203
rect 9689 11169 9723 11203
rect 9965 11169 9999 11203
rect 10241 11169 10275 11203
rect 10333 11169 10367 11203
rect 10609 11169 10643 11203
rect 10977 11169 11011 11203
rect 11437 11169 11471 11203
rect 11529 11169 11563 11203
rect 11989 11169 12023 11203
rect 12265 11169 12299 11203
rect 12357 11169 12391 11203
rect 12449 11169 12483 11203
rect 12633 11169 12667 11203
rect 12909 11169 12943 11203
rect 13185 11169 13219 11203
rect 13441 11169 13475 11203
rect 15117 11169 15151 11203
rect 15393 11169 15427 11203
rect 15485 11169 15519 11203
rect 15669 11169 15703 11203
rect 15945 11169 15979 11203
rect 16129 11169 16163 11203
rect 17969 11169 18003 11203
rect 18245 11169 18279 11203
rect 18429 11169 18463 11203
rect 18705 11169 18739 11203
rect 18797 11169 18831 11203
rect 19165 11169 19199 11203
rect 19257 11169 19291 11203
rect 19349 11169 19383 11203
rect 19809 11169 19843 11203
rect 19993 11169 20027 11203
rect 20177 11169 20211 11203
rect 20269 11169 20303 11203
rect 20545 11169 20579 11203
rect 20913 11169 20947 11203
rect 21465 11169 21499 11203
rect 21649 11169 21683 11203
rect 23397 11169 23431 11203
rect 23673 11169 23707 11203
rect 23765 11169 23799 11203
rect 23949 11169 23983 11203
rect 24409 11169 24443 11203
rect 24501 11169 24535 11203
rect 24777 11169 24811 11203
rect 25237 11169 25271 11203
rect 25329 11169 25363 11203
rect 9045 11101 9079 11135
rect 20637 11101 20671 11135
rect 21925 11101 21959 11135
rect 8217 11033 8251 11067
rect 8493 11033 8527 11067
rect 9873 11033 9907 11067
rect 11345 11033 11379 11067
rect 12173 11033 12207 11067
rect 12725 11033 12759 11067
rect 15025 11033 15059 11067
rect 17601 11033 17635 11067
rect 20085 11033 20119 11067
rect 8769 10965 8803 10999
rect 9597 10965 9631 10999
rect 10149 10965 10183 10999
rect 10701 10965 10735 10999
rect 11069 10965 11103 10999
rect 11897 10965 11931 10999
rect 13001 10965 13035 10999
rect 15301 10965 15335 10999
rect 15853 10965 15887 10999
rect 18061 10965 18095 10999
rect 18613 10965 18647 10999
rect 18889 10965 18923 10999
rect 21373 10965 21407 10999
rect 23489 10965 23523 10999
rect 24041 10965 24075 10999
rect 24317 10965 24351 10999
rect 24593 10965 24627 10999
rect 24869 10965 24903 10999
rect 25145 10965 25179 10999
rect 25421 10965 25455 10999
rect 7573 10761 7607 10795
rect 8493 10761 8527 10795
rect 9597 10761 9631 10795
rect 13277 10761 13311 10795
rect 16037 10761 16071 10795
rect 16865 10761 16899 10795
rect 19349 10761 19383 10795
rect 21925 10761 21959 10795
rect 24225 10761 24259 10795
rect 24501 10761 24535 10795
rect 24777 10761 24811 10795
rect 25329 10761 25363 10795
rect 15301 10693 15335 10727
rect 18429 10693 18463 10727
rect 20269 10693 20303 10727
rect 23581 10693 23615 10727
rect 17049 10625 17083 10659
rect 19625 10625 19659 10659
rect 21373 10625 21407 10659
rect 23949 10625 23983 10659
rect 7481 10557 7515 10591
rect 7941 10557 7975 10591
rect 8217 10557 8251 10591
rect 8585 10557 8619 10591
rect 8677 10557 8711 10591
rect 9137 10557 9171 10591
rect 9413 10557 9447 10591
rect 9689 10557 9723 10591
rect 9965 10557 9999 10591
rect 10057 10557 10091 10591
rect 11805 10557 11839 10591
rect 11897 10557 11931 10591
rect 13829 10557 13863 10591
rect 13921 10557 13955 10591
rect 15853 10557 15887 10591
rect 16129 10557 16163 10591
rect 16405 10557 16439 10591
rect 16589 10557 16623 10591
rect 16681 10557 16715 10591
rect 16957 10557 16991 10591
rect 18705 10557 18739 10591
rect 18981 10557 19015 10591
rect 19257 10557 19291 10591
rect 19717 10557 19751 10591
rect 19809 10557 19843 10591
rect 20361 10557 20395 10591
rect 20453 10557 20487 10591
rect 20637 10557 20671 10591
rect 20729 10557 20763 10591
rect 21189 10557 21223 10591
rect 21465 10557 21499 10591
rect 21741 10557 21775 10591
rect 21833 10557 21867 10591
rect 22201 10557 22235 10591
rect 23857 10557 23891 10591
rect 24317 10557 24351 10591
rect 24409 10557 24443 10591
rect 24685 10557 24719 10591
rect 25145 10557 25179 10591
rect 25421 10557 25455 10591
rect 25605 10557 25639 10591
rect 25697 10557 25731 10591
rect 11538 10489 11572 10523
rect 12142 10489 12176 10523
rect 14166 10489 14200 10523
rect 17316 10489 17350 10523
rect 19073 10489 19107 10523
rect 20545 10489 20579 10523
rect 21097 10489 21131 10523
rect 22468 10489 22502 10523
rect 25053 10489 25087 10523
rect 7849 10421 7883 10455
rect 8125 10421 8159 10455
rect 8769 10421 8803 10455
rect 9045 10421 9079 10455
rect 9321 10421 9355 10455
rect 9873 10421 9907 10455
rect 10149 10421 10183 10455
rect 10425 10421 10459 10455
rect 13737 10421 13771 10455
rect 15761 10421 15795 10455
rect 16313 10421 16347 10455
rect 18797 10421 18831 10455
rect 19901 10421 19935 10455
rect 20821 10421 20855 10455
rect 21649 10421 21683 10455
rect 8033 10217 8067 10251
rect 8861 10217 8895 10251
rect 9137 10217 9171 10251
rect 12541 10217 12575 10251
rect 13369 10217 13403 10251
rect 13645 10217 13679 10251
rect 13921 10217 13955 10251
rect 15577 10217 15611 10251
rect 16773 10217 16807 10251
rect 18613 10217 18647 10251
rect 20729 10217 20763 10251
rect 22017 10217 22051 10251
rect 23857 10217 23891 10251
rect 11437 10149 11471 10183
rect 19064 10149 19098 10183
rect 20913 10149 20947 10183
rect 7021 10081 7055 10115
rect 7297 10081 7331 10115
rect 7389 10081 7423 10115
rect 7573 10081 7607 10115
rect 7849 10081 7883 10115
rect 7941 10081 7975 10115
rect 8125 10081 8159 10115
rect 8401 10081 8435 10115
rect 8677 10081 8711 10115
rect 8769 10081 8803 10115
rect 8953 10081 8987 10115
rect 10250 10081 10284 10115
rect 10793 10081 10827 10115
rect 11253 10081 11287 10115
rect 11529 10081 11563 10115
rect 11805 10081 11839 10115
rect 12081 10081 12115 10115
rect 12173 10081 12207 10115
rect 12449 10081 12483 10115
rect 12909 10081 12943 10115
rect 13185 10081 13219 10115
rect 13277 10081 13311 10115
rect 13737 10081 13771 10115
rect 14013 10081 14047 10115
rect 14105 10081 14139 10115
rect 14381 10081 14415 10115
rect 14841 10081 14875 10115
rect 14933 10081 14967 10115
rect 15209 10081 15243 10115
rect 15669 10081 15703 10115
rect 15761 10081 15795 10115
rect 16313 10081 16347 10115
rect 16405 10081 16439 10115
rect 16681 10081 16715 10115
rect 17141 10081 17175 10115
rect 17500 10081 17534 10115
rect 18797 10081 18831 10115
rect 20545 10081 20579 10115
rect 20729 10081 20763 10115
rect 21005 10081 21039 10115
rect 21373 10081 21407 10115
rect 21465 10081 21499 10115
rect 21649 10081 21683 10115
rect 22109 10081 22143 10115
rect 22385 10081 22419 10115
rect 22744 10081 22778 10115
rect 24041 10081 24075 10115
rect 24317 10081 24351 10115
rect 24593 10081 24627 10115
rect 24869 10081 24903 10115
rect 25145 10081 25179 10115
rect 25329 10081 25363 10115
rect 25605 10081 25639 10115
rect 25789 10081 25823 10115
rect 25881 10081 25915 10115
rect 25973 10081 26007 10115
rect 10517 10013 10551 10047
rect 14197 10013 14231 10047
rect 15853 10013 15887 10047
rect 17233 10013 17267 10047
rect 22293 10013 22327 10047
rect 22477 10013 22511 10047
rect 7205 9945 7239 9979
rect 12817 9945 12851 9979
rect 17049 9945 17083 9979
rect 21741 9945 21775 9979
rect 24961 9945 24995 9979
rect 6929 9877 6963 9911
rect 7481 9877 7515 9911
rect 7757 9877 7791 9911
rect 8309 9877 8343 9911
rect 8585 9877 8619 9911
rect 10701 9877 10735 9911
rect 11161 9877 11195 9911
rect 11713 9877 11747 9911
rect 11989 9877 12023 9911
rect 12265 9877 12299 9911
rect 13093 9877 13127 9911
rect 14473 9877 14507 9911
rect 14749 9877 14783 9911
rect 15025 9877 15059 9911
rect 15301 9877 15335 9911
rect 16221 9877 16255 9911
rect 16497 9877 16531 9911
rect 20177 9877 20211 9911
rect 24133 9877 24167 9911
rect 24409 9877 24443 9911
rect 24685 9877 24719 9911
rect 25237 9877 25271 9911
rect 25513 9877 25547 9911
rect 26065 9877 26099 9911
rect 7297 9673 7331 9707
rect 7849 9673 7883 9707
rect 13277 9673 13311 9707
rect 13921 9673 13955 9707
rect 14197 9673 14231 9707
rect 15301 9673 15335 9707
rect 24501 9673 24535 9707
rect 25053 9673 25087 9707
rect 25605 9673 25639 9707
rect 26709 9673 26743 9707
rect 6193 9605 6227 9639
rect 7021 9605 7055 9639
rect 8677 9605 8711 9639
rect 10793 9605 10827 9639
rect 11069 9605 11103 9639
rect 11897 9605 11931 9639
rect 14749 9605 14783 9639
rect 15853 9605 15887 9639
rect 17509 9605 17543 9639
rect 17969 9605 18003 9639
rect 20913 9605 20947 9639
rect 23397 9605 23431 9639
rect 24777 9605 24811 9639
rect 12725 9537 12759 9571
rect 15577 9537 15611 9571
rect 18705 9537 18739 9571
rect 6285 9469 6319 9503
rect 6469 9469 6503 9503
rect 6561 9469 6595 9503
rect 6837 9469 6871 9503
rect 7113 9469 7147 9503
rect 7205 9469 7239 9503
rect 7481 9469 7515 9503
rect 7949 9469 7983 9503
rect 8225 9479 8259 9513
rect 10057 9469 10091 9503
rect 10333 9469 10367 9503
rect 10425 9469 10459 9503
rect 10885 9469 10919 9503
rect 10977 9469 11011 9503
rect 11161 9469 11195 9503
rect 11437 9469 11471 9503
rect 11529 9469 11563 9503
rect 11713 9469 11747 9503
rect 11989 9469 12023 9503
rect 12265 9469 12299 9503
rect 12357 9469 12391 9503
rect 12541 9469 12575 9503
rect 12817 9469 12851 9503
rect 13093 9469 13127 9503
rect 13369 9469 13403 9503
rect 13553 9469 13587 9503
rect 13737 9469 13771 9503
rect 14013 9469 14047 9503
rect 14105 9469 14139 9503
rect 14565 9469 14599 9503
rect 14657 9469 14691 9503
rect 14933 9469 14967 9503
rect 15393 9469 15427 9503
rect 15669 9469 15703 9503
rect 15945 9469 15979 9503
rect 18061 9469 18095 9503
rect 18153 9469 18187 9503
rect 18961 9469 18995 9503
rect 20361 9469 20395 9503
rect 20453 9469 20487 9503
rect 20545 9469 20579 9503
rect 20637 9469 20671 9503
rect 20821 9469 20855 9503
rect 21373 9469 21407 9503
rect 21649 9469 21683 9503
rect 21925 9469 21959 9503
rect 22017 9469 22051 9503
rect 22284 9469 22318 9503
rect 23857 9469 23891 9503
rect 24133 9469 24167 9503
rect 24409 9469 24443 9503
rect 24685 9469 24719 9503
rect 24961 9469 24995 9503
rect 25237 9469 25271 9503
rect 25329 9469 25363 9503
rect 25513 9469 25547 9503
rect 25789 9469 25823 9503
rect 25881 9469 25915 9503
rect 26065 9469 26099 9503
rect 26341 9469 26375 9503
rect 26801 9469 26835 9503
rect 26893 9469 26927 9503
rect 8125 9401 8159 9435
rect 9790 9401 9824 9435
rect 12173 9401 12207 9435
rect 12449 9401 12483 9435
rect 13001 9401 13035 9435
rect 13645 9401 13679 9435
rect 14473 9401 14507 9435
rect 16037 9401 16071 9435
rect 21833 9401 21867 9435
rect 6745 9333 6779 9367
rect 7573 9333 7607 9367
rect 10241 9333 10275 9367
rect 10517 9333 10551 9367
rect 11345 9333 11379 9367
rect 11713 9333 11747 9367
rect 15025 9333 15059 9367
rect 18245 9333 18279 9367
rect 20085 9333 20119 9367
rect 21281 9333 21315 9367
rect 21557 9333 21591 9367
rect 23949 9333 23983 9367
rect 24225 9333 24259 9367
rect 26157 9333 26191 9367
rect 26433 9333 26467 9367
rect 26985 9333 27019 9367
rect 6653 9129 6687 9163
rect 7941 9129 7975 9163
rect 9321 9129 9355 9163
rect 10425 9129 10459 9163
rect 10701 9129 10735 9163
rect 13185 9129 13219 9163
rect 15025 9129 15059 9163
rect 15761 9129 15795 9163
rect 18061 9129 18095 9163
rect 21097 9129 21131 9163
rect 21925 9129 21959 9163
rect 25973 9129 26007 9163
rect 9873 9061 9907 9095
rect 12909 9061 12943 9095
rect 17877 9061 17911 9095
rect 21649 9061 21683 9095
rect 22385 9061 22419 9095
rect 6469 8993 6503 9027
rect 6653 8993 6687 9027
rect 6745 8993 6779 9027
rect 7205 8993 7239 9027
rect 7481 8993 7515 9027
rect 7573 8993 7607 9027
rect 7849 8993 7883 9027
rect 8125 8993 8159 9027
rect 8401 8993 8435 9027
rect 8677 8993 8711 9027
rect 8953 8993 8987 9027
rect 9413 8993 9447 9027
rect 9505 8993 9539 9027
rect 9965 8993 9999 9027
rect 10241 8993 10275 9027
rect 10517 8993 10551 9027
rect 10609 8993 10643 9027
rect 12725 8993 12759 9027
rect 13001 8993 13035 9027
rect 13277 8993 13311 9027
rect 13625 8993 13659 9027
rect 15117 8993 15151 9027
rect 15301 8993 15335 9027
rect 15393 8993 15427 9027
rect 15669 8993 15703 9027
rect 15761 8993 15795 9027
rect 15945 8993 15979 9027
rect 18153 8993 18187 9027
rect 18245 8993 18279 9027
rect 18521 8993 18555 9027
rect 20453 8993 20487 9027
rect 20545 8993 20579 9027
rect 20913 8993 20947 9027
rect 21097 8993 21131 9027
rect 21281 8993 21315 9027
rect 21557 8993 21591 9027
rect 21833 8993 21867 9027
rect 22109 8993 22143 9027
rect 24492 8993 24526 9027
rect 25789 8993 25823 9027
rect 25973 8993 26007 9027
rect 26065 8993 26099 9027
rect 26525 8993 26559 9027
rect 26617 8993 26651 9027
rect 7113 8925 7147 8959
rect 7389 8925 7423 8959
rect 13369 8925 13403 8959
rect 16129 8925 16163 8959
rect 18797 8925 18831 8959
rect 21373 8925 21407 8959
rect 24225 8925 24259 8959
rect 6837 8857 6871 8891
rect 7665 8857 7699 8891
rect 11253 8857 11287 8891
rect 8217 8789 8251 8823
rect 8493 8789 8527 8823
rect 8769 8789 8803 8823
rect 9045 8789 9079 8823
rect 9597 8789 9631 8823
rect 10149 8789 10183 8823
rect 14749 8789 14783 8823
rect 15577 8789 15611 8823
rect 18337 8789 18371 8823
rect 20085 8789 20119 8823
rect 20361 8789 20395 8823
rect 20637 8789 20671 8823
rect 22201 8789 22235 8823
rect 23857 8789 23891 8823
rect 25605 8789 25639 8823
rect 26157 8789 26191 8823
rect 8125 8585 8159 8619
rect 8585 8585 8619 8619
rect 10885 8585 10919 8619
rect 11161 8585 11195 8619
rect 14381 8585 14415 8619
rect 17785 8585 17819 8619
rect 19349 8585 19383 8619
rect 20177 8585 20211 8619
rect 21281 8585 21315 8619
rect 24225 8585 24259 8619
rect 25329 8585 25363 8619
rect 7297 8517 7331 8551
rect 8861 8517 8895 8551
rect 13829 8517 13863 8551
rect 14105 8517 14139 8551
rect 15945 8517 15979 8551
rect 22845 8517 22879 8551
rect 23397 8517 23431 8551
rect 26709 8517 26743 8551
rect 7573 8449 7607 8483
rect 10241 8449 10275 8483
rect 11621 8449 11655 8483
rect 14565 8449 14599 8483
rect 18061 8449 18095 8483
rect 19901 8449 19935 8483
rect 21465 8449 21499 8483
rect 23949 8449 23983 8483
rect 6745 8381 6779 8415
rect 6837 8381 6871 8415
rect 7021 8381 7055 8415
rect 7113 8381 7147 8415
rect 7389 8381 7423 8415
rect 7481 8381 7515 8415
rect 7757 8381 7791 8415
rect 8033 8381 8067 8415
rect 8493 8381 8527 8415
rect 10517 8381 10551 8415
rect 10793 8381 10827 8415
rect 11069 8381 11103 8415
rect 11345 8381 11379 8415
rect 13185 8381 13219 8415
rect 13737 8381 13771 8415
rect 14013 8381 14047 8415
rect 14473 8381 14507 8415
rect 16129 8381 16163 8415
rect 17877 8381 17911 8415
rect 17969 8381 18003 8415
rect 18429 8381 18463 8415
rect 18705 8381 18739 8415
rect 18981 8381 19015 8415
rect 19441 8381 19475 8415
rect 19533 8381 19567 8415
rect 19625 8381 19659 8415
rect 19809 8381 19843 8415
rect 20269 8381 20303 8415
rect 20545 8381 20579 8415
rect 20645 8381 20679 8415
rect 20913 8381 20947 8415
rect 21097 8381 21131 8415
rect 21189 8381 21223 8415
rect 23029 8381 23063 8415
rect 23213 8381 23247 8415
rect 23305 8381 23339 8415
rect 23857 8381 23891 8415
rect 24133 8381 24167 8415
rect 24409 8381 24443 8415
rect 24869 8381 24903 8415
rect 25145 8381 25179 8415
rect 25421 8381 25455 8415
rect 25697 8381 25731 8415
rect 25789 8381 25823 8415
rect 26065 8381 26099 8415
rect 26341 8381 26375 8415
rect 26433 8381 26467 8415
rect 26617 8381 26651 8415
rect 7849 8313 7883 8347
rect 9974 8313 10008 8347
rect 11437 8313 11471 8347
rect 11866 8313 11900 8347
rect 14832 8313 14866 8347
rect 16374 8313 16408 8347
rect 18337 8313 18371 8347
rect 18797 8313 18831 8347
rect 19073 8313 19107 8347
rect 20453 8313 20487 8347
rect 21005 8313 21039 8347
rect 21732 8313 21766 8347
rect 24501 8313 24535 8347
rect 10609 8245 10643 8279
rect 13001 8245 13035 8279
rect 13277 8245 13311 8279
rect 17509 8245 17543 8279
rect 20729 8245 20763 8279
rect 23029 8245 23063 8279
rect 24777 8245 24811 8279
rect 25053 8245 25087 8279
rect 25605 8245 25639 8279
rect 25881 8245 25915 8279
rect 26157 8245 26191 8279
rect 9045 8041 9079 8075
rect 10425 8041 10459 8075
rect 20913 8041 20947 8075
rect 10977 7973 11011 8007
rect 12725 7973 12759 8007
rect 13522 7973 13556 8007
rect 15301 7973 15335 8007
rect 18337 7973 18371 8007
rect 20085 7973 20119 8007
rect 21281 7973 21315 8007
rect 22845 7973 22879 8007
rect 23388 7973 23422 8007
rect 7205 7905 7239 7939
rect 7389 7905 7423 7939
rect 7481 7905 7515 7939
rect 7757 7905 7791 7939
rect 8033 7905 8067 7939
rect 8309 7905 8343 7939
rect 8401 7905 8435 7939
rect 8677 7905 8711 7939
rect 8953 7905 8987 7939
rect 9413 7905 9447 7939
rect 9689 7905 9723 7939
rect 9965 7905 9999 7939
rect 10241 7905 10275 7939
rect 10333 7905 10367 7939
rect 10609 7905 10643 7939
rect 13001 7905 13035 7939
rect 13277 7905 13311 7939
rect 14933 7905 14967 7939
rect 15401 7903 15435 7937
rect 15577 7905 15611 7939
rect 15669 7905 15703 7939
rect 15761 7905 15795 7939
rect 16221 7905 16255 7939
rect 16497 7905 16531 7939
rect 16773 7905 16807 7939
rect 17040 7905 17074 7939
rect 20177 7905 20211 7939
rect 20453 7905 20487 7939
rect 21005 7905 21039 7939
rect 23110 7905 23144 7939
rect 24685 7905 24719 7939
rect 24961 7905 24995 7939
rect 25237 7905 25271 7939
rect 25697 7905 25731 7939
rect 25789 7895 25823 7929
rect 26065 7905 26099 7939
rect 7941 7837 7975 7871
rect 8769 7837 8803 7871
rect 13093 7837 13127 7871
rect 24777 7837 24811 7871
rect 25329 7837 25363 7871
rect 8493 7769 8527 7803
rect 10149 7769 10183 7803
rect 20545 7769 20579 7803
rect 7113 7701 7147 7735
rect 7665 7701 7699 7735
rect 8217 7701 8251 7735
rect 9321 7701 9355 7735
rect 9597 7701 9631 7735
rect 9873 7701 9907 7735
rect 10701 7701 10735 7735
rect 14657 7701 14691 7735
rect 15025 7701 15059 7735
rect 15853 7701 15887 7735
rect 16313 7701 16347 7735
rect 16589 7701 16623 7735
rect 18153 7701 18187 7735
rect 20269 7701 20303 7735
rect 24501 7701 24535 7735
rect 25053 7701 25087 7735
rect 25605 7701 25639 7735
rect 25881 7701 25915 7735
rect 26157 7701 26191 7735
rect 7021 7497 7055 7531
rect 8861 7497 8895 7531
rect 9137 7497 9171 7531
rect 10701 7497 10735 7531
rect 14381 7497 14415 7531
rect 15485 7497 15519 7531
rect 15761 7497 15795 7531
rect 24501 7497 24535 7531
rect 24777 7497 24811 7531
rect 25605 7497 25639 7531
rect 6239 7429 6273 7463
rect 7297 7429 7331 7463
rect 19349 7429 19383 7463
rect 23581 7429 23615 7463
rect 25053 7429 25087 7463
rect 10057 7361 10091 7395
rect 16589 7361 16623 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 18797 7361 18831 7395
rect 19625 7361 19659 7395
rect 21925 7361 21959 7395
rect 6168 7293 6202 7327
rect 6423 7293 6457 7327
rect 6526 7293 6560 7327
rect 6720 7293 6754 7327
rect 7113 7293 7147 7327
rect 7205 7293 7239 7327
rect 7657 7293 7691 7327
rect 7757 7293 7791 7327
rect 7941 7293 7975 7327
rect 8217 7293 8251 7327
rect 8677 7293 8711 7327
rect 8953 7295 8987 7329
rect 9045 7293 9079 7327
rect 9229 7293 9263 7327
rect 9321 7293 9355 7327
rect 9413 7293 9447 7327
rect 9781 7293 9815 7327
rect 10333 7293 10367 7327
rect 10609 7293 10643 7327
rect 10885 7293 10919 7327
rect 11069 7293 11103 7327
rect 11345 7293 11379 7327
rect 11621 7293 11655 7327
rect 12918 7293 12952 7327
rect 13185 7293 13219 7327
rect 13737 7293 13771 7327
rect 14013 7293 14047 7327
rect 14289 7293 14323 7327
rect 14565 7293 14599 7327
rect 14749 7293 14783 7327
rect 15025 7293 15059 7327
rect 15301 7293 15335 7327
rect 15577 7293 15611 7327
rect 15853 7293 15887 7327
rect 16037 7293 16071 7327
rect 16129 7293 16163 7327
rect 16221 7293 16255 7327
rect 16405 7293 16439 7327
rect 16673 7293 16707 7327
rect 16957 7293 16991 7327
rect 18705 7293 18739 7327
rect 19165 7293 19199 7327
rect 19257 7293 19291 7327
rect 19533 7293 19567 7327
rect 19993 7293 20027 7327
rect 20269 7295 20303 7329
rect 20361 7293 20395 7327
rect 20637 7293 20671 7327
rect 20729 7293 20763 7327
rect 20913 7293 20947 7327
rect 21189 7293 21223 7327
rect 21281 7293 21315 7327
rect 21465 7293 21499 7327
rect 22192 7293 22226 7327
rect 23673 7293 23707 7327
rect 23857 7293 23891 7327
rect 24041 7293 24075 7327
rect 24317 7293 24351 7327
rect 24593 7293 24627 7327
rect 24685 7293 24719 7327
rect 24961 7293 24995 7327
rect 25421 7293 25455 7327
rect 25513 7293 25547 7327
rect 7849 7225 7883 7259
rect 13829 7225 13863 7259
rect 16313 7225 16347 7259
rect 17316 7225 17350 7259
rect 23949 7225 23983 7259
rect 6791 7157 6825 7191
rect 7573 7157 7607 7191
rect 8125 7157 8159 7191
rect 8585 7157 8619 7191
rect 9689 7157 9723 7191
rect 11069 7157 11103 7191
rect 11253 7157 11287 7191
rect 11529 7157 11563 7191
rect 11805 7157 11839 7191
rect 14105 7157 14139 7191
rect 14749 7157 14783 7191
rect 14933 7157 14967 7191
rect 15209 7157 15243 7191
rect 18429 7157 18463 7191
rect 19073 7157 19107 7191
rect 19901 7157 19935 7191
rect 20177 7157 20211 7191
rect 20453 7157 20487 7191
rect 21005 7157 21039 7191
rect 21557 7157 21591 7191
rect 23305 7157 23339 7191
rect 24225 7157 24259 7191
rect 25329 7157 25363 7191
rect 7343 6953 7377 6987
rect 8217 6953 8251 6987
rect 9229 6953 9263 6987
rect 10425 6953 10459 6987
rect 12265 6953 12299 6987
rect 15853 6953 15887 6987
rect 16589 6953 16623 6987
rect 19533 6953 19567 6987
rect 24869 6953 24903 6987
rect 11161 6885 11195 6919
rect 11713 6885 11747 6919
rect 6260 6817 6294 6851
rect 6536 6817 6570 6851
rect 6812 6817 6846 6851
rect 7056 6817 7090 6851
rect 7446 6817 7480 6851
rect 7573 6817 7607 6851
rect 7849 6817 7883 6851
rect 8125 6817 8159 6851
rect 8493 6817 8527 6851
rect 8585 6817 8619 6851
rect 8677 6807 8711 6841
rect 8861 6817 8895 6851
rect 9321 6817 9355 6851
rect 9505 6817 9539 6851
rect 9597 6817 9631 6851
rect 10517 6817 10551 6851
rect 10609 6817 10643 6851
rect 10701 6817 10735 6851
rect 11253 6817 11287 6851
rect 11345 6807 11379 6841
rect 11437 6817 11471 6851
rect 11621 6817 11655 6851
rect 11897 6817 11931 6851
rect 12357 6817 12391 6851
rect 12705 6817 12739 6851
rect 14464 6817 14498 6851
rect 15945 6817 15979 6851
rect 16405 6817 16439 6851
rect 16681 6817 16715 6851
rect 16957 6817 16991 6851
rect 18981 6817 19015 6851
rect 19073 6817 19107 6851
rect 19349 6817 19383 6851
rect 19533 6817 19567 6851
rect 19809 6817 19843 6851
rect 20085 6817 20119 6851
rect 20177 6817 20211 6851
rect 20453 6817 20487 6851
rect 20637 6817 20671 6851
rect 20913 6817 20947 6851
rect 21281 6817 21315 6851
rect 21548 6817 21582 6851
rect 23029 6817 23063 6851
rect 23121 6817 23155 6851
rect 23581 6817 23615 6851
rect 23673 6817 23707 6851
rect 23949 6817 23983 6851
rect 24225 6817 24259 6851
rect 24317 6817 24351 6851
rect 24501 6817 24535 6851
rect 24685 6817 24719 6851
rect 24777 6817 24811 6851
rect 8769 6749 8803 6783
rect 10149 6749 10183 6783
rect 12449 6749 12483 6783
rect 14197 6749 14231 6783
rect 16313 6749 16347 6783
rect 19165 6749 19199 6783
rect 7941 6681 7975 6715
rect 9781 6681 9815 6715
rect 18245 6681 18279 6715
rect 19993 6681 20027 6715
rect 24041 6681 24075 6715
rect 6331 6613 6365 6647
rect 6607 6613 6641 6647
rect 6883 6613 6917 6647
rect 7159 6613 7193 6647
rect 7757 6613 7791 6647
rect 9689 6613 9723 6647
rect 11989 6613 12023 6647
rect 13829 6613 13863 6647
rect 15577 6613 15611 6647
rect 18889 6613 18923 6647
rect 19717 6613 19751 6647
rect 20269 6613 20303 6647
rect 20545 6613 20579 6647
rect 20821 6613 20855 6647
rect 22661 6613 22695 6647
rect 22937 6613 22971 6647
rect 23213 6613 23247 6647
rect 23489 6613 23523 6647
rect 23765 6613 23799 6647
rect 24593 6613 24627 6647
rect 8079 6409 8113 6443
rect 8539 6409 8573 6443
rect 10517 6409 10551 6443
rect 12725 6409 12759 6443
rect 17785 6409 17819 6443
rect 19073 6409 19107 6443
rect 21189 6409 21223 6443
rect 21741 6409 21775 6443
rect 22569 6409 22603 6443
rect 22845 6409 22879 6443
rect 23949 6409 23983 6443
rect 9689 6341 9723 6375
rect 13001 6341 13035 6375
rect 13277 6341 13311 6375
rect 17509 6341 17543 6375
rect 18337 6341 18371 6375
rect 24225 6341 24259 6375
rect 10149 6273 10183 6307
rect 10333 6273 10367 6307
rect 11069 6273 11103 6307
rect 7354 6205 7388 6239
rect 7527 6205 7561 6239
rect 7630 6205 7664 6239
rect 7874 6205 7908 6239
rect 8150 6205 8184 6239
rect 8436 6205 8470 6239
rect 8677 6205 8711 6239
rect 8861 6205 8895 6239
rect 9413 6205 9447 6239
rect 9505 6205 9539 6239
rect 10057 6205 10091 6239
rect 10609 6205 10643 6239
rect 10793 6205 10827 6239
rect 12817 6205 12851 6239
rect 13093 6205 13127 6239
rect 13185 6205 13219 6239
rect 13829 6205 13863 6239
rect 15669 6205 15703 6239
rect 15853 6205 15887 6239
rect 16129 6205 16163 6239
rect 17877 6205 17911 6239
rect 18061 6205 18095 6239
rect 18153 6205 18187 6239
rect 18429 6205 18463 6239
rect 18889 6205 18923 6239
rect 18981 6205 19015 6239
rect 19441 6205 19475 6239
rect 19533 6205 19567 6239
rect 21097 6205 21131 6239
rect 21557 6205 21591 6239
rect 21649 6205 21683 6239
rect 22109 6205 22143 6239
rect 22201 6205 22235 6239
rect 22661 6205 22695 6239
rect 22753 6205 22787 6239
rect 23213 6205 23247 6239
rect 23305 6205 23339 6239
rect 23489 6205 23523 6239
rect 23857 6215 23891 6249
rect 24317 6205 24351 6239
rect 8953 6137 8987 6171
rect 9137 6137 9171 6171
rect 9689 6137 9723 6171
rect 10333 6137 10367 6171
rect 10885 6137 10919 6171
rect 11336 6137 11370 6171
rect 13737 6137 13771 6171
rect 13921 6137 13955 6171
rect 15945 6137 15979 6171
rect 16374 6137 16408 6171
rect 18797 6137 18831 6171
rect 19800 6137 19834 6171
rect 7251 6069 7285 6103
rect 7803 6069 7837 6103
rect 8769 6069 8803 6103
rect 9321 6069 9355 6103
rect 12449 6069 12483 6103
rect 19349 6069 19383 6103
rect 20913 6069 20947 6103
rect 21465 6069 21499 6103
rect 22017 6069 22051 6103
rect 22293 6069 22327 6103
rect 23121 6069 23155 6103
rect 23305 6069 23339 6103
rect 7803 5865 7837 5899
rect 8585 5865 8619 5899
rect 9137 5865 9171 5899
rect 10793 5865 10827 5899
rect 14381 5865 14415 5899
rect 19349 5865 19383 5899
rect 22753 5865 22787 5899
rect 12550 5797 12584 5831
rect 14718 5797 14752 5831
rect 21373 5797 21407 5831
rect 23029 5797 23063 5831
rect 7700 5729 7734 5763
rect 8058 5729 8092 5763
rect 8401 5729 8435 5763
rect 8493 5729 8527 5763
rect 8886 5729 8920 5763
rect 9229 5729 9263 5763
rect 9680 5729 9714 5763
rect 11069 5729 11103 5763
rect 13268 5729 13302 5763
rect 14473 5729 14507 5763
rect 16385 5729 16419 5763
rect 17693 5729 17727 5763
rect 17960 5729 17994 5763
rect 19257 5729 19291 5763
rect 19533 5729 19567 5763
rect 19993 5729 20027 5763
rect 20177 5729 20211 5763
rect 20269 5729 20303 5763
rect 20545 5729 20579 5763
rect 20637 5729 20671 5763
rect 20821 5729 20855 5763
rect 21097 5729 21131 5763
rect 21465 5729 21499 5763
rect 21649 5729 21683 5763
rect 21741 5729 21775 5763
rect 22017 5729 22051 5763
rect 22293 5729 22327 5763
rect 22385 5729 22419 5763
rect 22477 5729 22511 5763
rect 22661 5729 22695 5763
rect 23121 5729 23155 5763
rect 23397 5729 23431 5763
rect 9413 5661 9447 5695
rect 11161 5661 11195 5695
rect 12817 5661 12851 5695
rect 13001 5661 13035 5695
rect 16129 5661 16163 5695
rect 19625 5661 19659 5695
rect 21005 5661 21039 5695
rect 7987 5593 8021 5627
rect 8309 5593 8343 5627
rect 19073 5593 19107 5627
rect 23305 5593 23339 5627
rect 8815 5525 8849 5559
rect 11437 5525 11471 5559
rect 15853 5525 15887 5559
rect 17509 5525 17543 5559
rect 19901 5525 19935 5559
rect 20453 5525 20487 5559
rect 20729 5525 20763 5559
rect 21925 5525 21959 5559
rect 22201 5525 22235 5559
rect 10149 5321 10183 5355
rect 12541 5321 12575 5355
rect 13093 5321 13127 5355
rect 15301 5321 15335 5355
rect 16313 5321 16347 5355
rect 16681 5321 16715 5355
rect 19257 5321 19291 5355
rect 19533 5321 19567 5355
rect 21465 5321 21499 5355
rect 21741 5321 21775 5355
rect 22293 5321 22327 5355
rect 10701 5253 10735 5287
rect 18797 5253 18831 5287
rect 19809 5253 19843 5287
rect 10885 5185 10919 5219
rect 13737 5185 13771 5219
rect 17049 5185 17083 5219
rect 8033 5117 8067 5151
rect 8401 5117 8435 5151
rect 10517 5117 10551 5151
rect 10609 5117 10643 5151
rect 10793 5117 10827 5151
rect 12449 5117 12483 5151
rect 12725 5117 12759 5151
rect 13829 5117 13863 5151
rect 13921 5117 13955 5151
rect 14013 5117 14047 5151
rect 14473 5117 14507 5151
rect 14565 5117 14599 5151
rect 14933 5117 14967 5151
rect 15209 5117 15243 5151
rect 15577 5117 15611 5151
rect 15853 5117 15887 5151
rect 16129 5117 16163 5151
rect 17316 5117 17350 5151
rect 18889 5117 18923 5151
rect 19157 5117 19191 5151
rect 19625 5117 19659 5151
rect 19901 5117 19935 5151
rect 19993 5117 20027 5151
rect 20453 5117 20487 5151
rect 20545 5117 20579 5151
rect 21005 5117 21039 5151
rect 21281 5117 21315 5151
rect 21557 5117 21591 5151
rect 21649 5117 21683 5151
rect 22109 5117 22143 5151
rect 22201 5117 22235 5151
rect 8646 5049 8680 5083
rect 11130 5049 11164 5083
rect 13093 5049 13127 5083
rect 14841 5049 14875 5083
rect 15669 5049 15703 5083
rect 16865 5049 16899 5083
rect 20361 5049 20395 5083
rect 22017 5049 22051 5083
rect 8217 4981 8251 5015
rect 9781 4981 9815 5015
rect 9965 4981 9999 5015
rect 10149 4981 10183 5015
rect 12265 4981 12299 5015
rect 13277 4981 13311 5015
rect 13553 4981 13587 5015
rect 14289 4981 14323 5015
rect 14657 4981 14691 5015
rect 15025 4981 15059 5015
rect 15945 4981 15979 5015
rect 16497 4981 16531 5015
rect 16665 4981 16699 5015
rect 18429 4981 18463 5015
rect 20085 4981 20119 5015
rect 20637 4981 20671 5015
rect 20913 4981 20947 5015
rect 21189 4981 21223 5015
rect 9873 4777 9907 4811
rect 10701 4777 10735 4811
rect 11805 4777 11839 4811
rect 13185 4777 13219 4811
rect 13461 4777 13495 4811
rect 16129 4777 16163 4811
rect 16589 4777 16623 4811
rect 9689 4709 9723 4743
rect 10241 4709 10275 4743
rect 9229 4641 9263 4675
rect 9505 4641 9539 4675
rect 9965 4641 9999 4675
rect 10149 4641 10183 4675
rect 10333 4641 10367 4675
rect 10793 4641 10827 4675
rect 11345 4641 11379 4675
rect 11437 4641 11471 4675
rect 11713 4641 11747 4675
rect 12081 4641 12115 4675
rect 12909 4641 12943 4675
rect 13093 4641 13127 4675
rect 13645 4641 13679 4675
rect 14013 4641 14047 4675
rect 14105 4641 14139 4675
rect 14289 4641 14323 4675
rect 14657 4641 14691 4675
rect 14749 4641 14783 4675
rect 15393 4641 15427 4675
rect 15669 4641 15703 4675
rect 15853 4641 15887 4675
rect 15945 4641 15979 4675
rect 16129 4641 16163 4675
rect 16313 4641 16347 4675
rect 16497 4641 16531 4675
rect 16957 4641 16991 4675
rect 17213 4641 17247 4675
rect 19901 4641 19935 4675
rect 20453 4641 20487 4675
rect 20729 4641 20763 4675
rect 20821 4641 20855 4675
rect 21005 4641 21039 4675
rect 11253 4573 11287 4607
rect 12357 4573 12391 4607
rect 12817 4573 12851 4607
rect 20637 4573 20671 4607
rect 10517 4505 10551 4539
rect 12265 4505 12299 4539
rect 15577 4505 15611 4539
rect 15945 4505 15979 4539
rect 20361 4505 20395 4539
rect 20913 4505 20947 4539
rect 9321 4437 9355 4471
rect 11529 4437 11563 4471
rect 12173 4437 12207 4471
rect 14289 4437 14323 4471
rect 18337 4437 18371 4471
rect 19993 4437 20027 4471
rect 9689 4233 9723 4267
rect 15301 4233 15335 4267
rect 10057 4165 10091 4199
rect 11253 4165 11287 4199
rect 15669 4097 15703 4131
rect 8953 4029 8987 4063
rect 10333 4029 10367 4063
rect 10609 4029 10643 4063
rect 10977 4029 11011 4063
rect 11253 4029 11287 4063
rect 11621 4029 11655 4063
rect 11877 4029 11911 4063
rect 13921 4029 13955 4063
rect 14188 4029 14222 4063
rect 15936 3961 15970 3995
rect 8769 3893 8803 3927
rect 9505 3893 9539 3927
rect 9689 3893 9723 3927
rect 10149 3893 10183 3927
rect 10517 3893 10551 3927
rect 11069 3893 11103 3927
rect 13001 3893 13035 3927
rect 17049 3893 17083 3927
rect 9873 3689 9907 3723
rect 10041 3689 10075 3723
rect 12633 3689 12667 3723
rect 14473 3689 14507 3723
rect 16129 3689 16163 3723
rect 8668 3621 8702 3655
rect 10241 3621 10275 3655
rect 12182 3621 12216 3655
rect 15393 3621 15427 3655
rect 17202 3621 17236 3655
rect 8401 3553 8435 3587
rect 12449 3553 12483 3587
rect 13746 3553 13780 3587
rect 14013 3553 14047 3587
rect 14197 3553 14231 3587
rect 15033 3553 15067 3587
rect 16313 3553 16347 3587
rect 16405 3553 16439 3587
rect 16957 3553 16991 3587
rect 14473 3485 14507 3519
rect 14933 3485 14967 3519
rect 14289 3417 14323 3451
rect 15761 3417 15795 3451
rect 16497 3417 16531 3451
rect 9781 3349 9815 3383
rect 10057 3349 10091 3383
rect 11069 3349 11103 3383
rect 15853 3349 15887 3383
rect 18337 3349 18371 3383
rect 8033 969 8067 1003
rect 7849 765 7883 799
<< metal1 >>
rect 552 19066 31531 19088
rect 552 19014 8102 19066
rect 8154 19014 8166 19066
rect 8218 19014 8230 19066
rect 8282 19014 8294 19066
rect 8346 19014 8358 19066
rect 8410 19014 15807 19066
rect 15859 19014 15871 19066
rect 15923 19014 15935 19066
rect 15987 19014 15999 19066
rect 16051 19014 16063 19066
rect 16115 19014 23512 19066
rect 23564 19014 23576 19066
rect 23628 19014 23640 19066
rect 23692 19014 23704 19066
rect 23756 19014 23768 19066
rect 23820 19014 31217 19066
rect 31269 19014 31281 19066
rect 31333 19014 31345 19066
rect 31397 19014 31409 19066
rect 31461 19014 31473 19066
rect 31525 19014 31531 19066
rect 552 18992 31531 19014
rect 552 18522 31372 18544
rect 552 18470 4250 18522
rect 4302 18470 4314 18522
rect 4366 18470 4378 18522
rect 4430 18470 4442 18522
rect 4494 18470 4506 18522
rect 4558 18470 11955 18522
rect 12007 18470 12019 18522
rect 12071 18470 12083 18522
rect 12135 18470 12147 18522
rect 12199 18470 12211 18522
rect 12263 18470 19660 18522
rect 19712 18470 19724 18522
rect 19776 18470 19788 18522
rect 19840 18470 19852 18522
rect 19904 18470 19916 18522
rect 19968 18470 27365 18522
rect 27417 18470 27429 18522
rect 27481 18470 27493 18522
rect 27545 18470 27557 18522
rect 27609 18470 27621 18522
rect 27673 18470 31372 18522
rect 552 18448 31372 18470
rect 552 17978 31531 18000
rect 552 17926 8102 17978
rect 8154 17926 8166 17978
rect 8218 17926 8230 17978
rect 8282 17926 8294 17978
rect 8346 17926 8358 17978
rect 8410 17926 15807 17978
rect 15859 17926 15871 17978
rect 15923 17926 15935 17978
rect 15987 17926 15999 17978
rect 16051 17926 16063 17978
rect 16115 17926 23512 17978
rect 23564 17926 23576 17978
rect 23628 17926 23640 17978
rect 23692 17926 23704 17978
rect 23756 17926 23768 17978
rect 23820 17926 31217 17978
rect 31269 17926 31281 17978
rect 31333 17926 31345 17978
rect 31397 17926 31409 17978
rect 31461 17926 31473 17978
rect 31525 17926 31531 17978
rect 552 17904 31531 17926
rect 20625 17731 20683 17737
rect 20625 17697 20637 17731
rect 20671 17728 20683 17731
rect 20671 17700 21036 17728
rect 20671 17697 20683 17700
rect 20625 17691 20683 17697
rect 21008 17604 21036 17700
rect 20990 17552 20996 17604
rect 21048 17552 21054 17604
rect 20717 17527 20775 17533
rect 20717 17493 20729 17527
rect 20763 17524 20775 17527
rect 21174 17524 21180 17536
rect 20763 17496 21180 17524
rect 20763 17493 20775 17496
rect 20717 17487 20775 17493
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 552 17434 31372 17456
rect 552 17382 4250 17434
rect 4302 17382 4314 17434
rect 4366 17382 4378 17434
rect 4430 17382 4442 17434
rect 4494 17382 4506 17434
rect 4558 17382 11955 17434
rect 12007 17382 12019 17434
rect 12071 17382 12083 17434
rect 12135 17382 12147 17434
rect 12199 17382 12211 17434
rect 12263 17382 19660 17434
rect 19712 17382 19724 17434
rect 19776 17382 19788 17434
rect 19840 17382 19852 17434
rect 19904 17382 19916 17434
rect 19968 17382 27365 17434
rect 27417 17382 27429 17434
rect 27481 17382 27493 17434
rect 27545 17382 27557 17434
rect 27609 17382 27621 17434
rect 27673 17382 31372 17434
rect 552 17360 31372 17382
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 12805 17323 12863 17329
rect 12805 17320 12817 17323
rect 11388 17292 12817 17320
rect 11388 17280 11394 17292
rect 12805 17289 12817 17292
rect 12851 17289 12863 17323
rect 12805 17283 12863 17289
rect 20257 17323 20315 17329
rect 20257 17289 20269 17323
rect 20303 17320 20315 17323
rect 21266 17320 21272 17332
rect 20303 17292 21272 17320
rect 20303 17289 20315 17292
rect 20257 17283 20315 17289
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 21361 17323 21419 17329
rect 21361 17289 21373 17323
rect 21407 17320 21419 17323
rect 21818 17320 21824 17332
rect 21407 17292 21824 17320
rect 21407 17289 21419 17292
rect 21361 17283 21419 17289
rect 21818 17280 21824 17292
rect 21876 17280 21882 17332
rect 21913 17323 21971 17329
rect 21913 17289 21925 17323
rect 21959 17320 21971 17323
rect 23290 17320 23296 17332
rect 21959 17292 23296 17320
rect 21959 17289 21971 17292
rect 21913 17283 21971 17289
rect 23290 17280 23296 17292
rect 23348 17280 23354 17332
rect 11609 17255 11667 17261
rect 11609 17252 11621 17255
rect 11256 17224 11621 17252
rect 11149 17129 11207 17135
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 11057 17119 11115 17125
rect 11057 17116 11069 17119
rect 9824 17088 11069 17116
rect 9824 17076 9830 17088
rect 11057 17085 11069 17088
rect 11103 17085 11115 17119
rect 11149 17095 11161 17129
rect 11195 17095 11207 17129
rect 11149 17089 11207 17095
rect 11256 17116 11284 17224
rect 11609 17221 11621 17224
rect 11655 17221 11667 17255
rect 11609 17215 11667 17221
rect 12342 17212 12348 17264
rect 12400 17252 12406 17264
rect 13081 17255 13139 17261
rect 13081 17252 13093 17255
rect 12400 17224 13093 17252
rect 12400 17212 12406 17224
rect 13081 17221 13093 17224
rect 13127 17221 13139 17255
rect 21085 17255 21143 17261
rect 13081 17215 13139 17221
rect 19260 17224 20944 17252
rect 12161 17187 12219 17193
rect 11532 17156 12112 17184
rect 11532 17128 11560 17156
rect 12084 17128 12112 17156
rect 12161 17153 12173 17187
rect 12207 17184 12219 17187
rect 12207 17156 12756 17184
rect 12207 17153 12219 17156
rect 12161 17147 12219 17153
rect 11425 17119 11483 17125
rect 11425 17116 11437 17119
rect 11057 17079 11115 17085
rect 11164 17060 11192 17089
rect 11256 17088 11437 17116
rect 11425 17085 11437 17088
rect 11471 17085 11483 17119
rect 11425 17079 11483 17085
rect 11514 17076 11520 17128
rect 11572 17116 11578 17128
rect 11701 17119 11759 17125
rect 11701 17116 11713 17119
rect 11572 17088 11713 17116
rect 11572 17076 11578 17088
rect 11701 17085 11713 17088
rect 11747 17085 11759 17119
rect 11701 17079 11759 17085
rect 11793 17119 11851 17125
rect 11793 17085 11805 17119
rect 11839 17085 11851 17119
rect 11793 17079 11851 17085
rect 8662 17008 8668 17060
rect 8720 17048 8726 17060
rect 8720 17020 11100 17048
rect 8720 17008 8726 17020
rect 11072 16980 11100 17020
rect 11146 17008 11152 17060
rect 11204 17008 11210 17060
rect 11238 17008 11244 17060
rect 11296 17048 11302 17060
rect 11808 17048 11836 17079
rect 11882 17076 11888 17128
rect 11940 17076 11946 17128
rect 12066 17076 12072 17128
rect 12124 17076 12130 17128
rect 12618 17076 12624 17128
rect 12676 17076 12682 17128
rect 12728 17125 12756 17156
rect 12713 17119 12771 17125
rect 12713 17085 12725 17119
rect 12759 17085 12771 17119
rect 12713 17079 12771 17085
rect 12986 17076 12992 17128
rect 13044 17076 13050 17128
rect 13725 17119 13783 17125
rect 13725 17085 13737 17119
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 11296 17020 11836 17048
rect 11900 17048 11928 17076
rect 13633 17051 13691 17057
rect 13633 17048 13645 17051
rect 11900 17020 13645 17048
rect 11296 17008 11302 17020
rect 13633 17017 13645 17020
rect 13679 17017 13691 17051
rect 13633 17011 13691 17017
rect 13740 16992 13768 17079
rect 13814 17076 13820 17128
rect 13872 17076 13878 17128
rect 13998 17076 14004 17128
rect 14056 17116 14062 17128
rect 14829 17119 14887 17125
rect 14829 17116 14841 17119
rect 14056 17088 14841 17116
rect 14056 17076 14062 17088
rect 14829 17085 14841 17088
rect 14875 17085 14887 17119
rect 14829 17079 14887 17085
rect 19260 16992 19288 17224
rect 19518 17144 19524 17196
rect 19576 17184 19582 17196
rect 19576 17156 20760 17184
rect 19576 17144 19582 17156
rect 20346 17076 20352 17128
rect 20404 17076 20410 17128
rect 20625 17121 20683 17127
rect 20732 17125 20760 17156
rect 20625 17087 20637 17121
rect 20671 17087 20683 17121
rect 20625 17081 20683 17087
rect 20717 17119 20775 17125
rect 20717 17085 20729 17119
rect 20763 17085 20775 17119
rect 20916 17116 20944 17224
rect 21085 17221 21097 17255
rect 21131 17252 21143 17255
rect 22094 17252 22100 17264
rect 21131 17224 22100 17252
rect 21131 17221 21143 17224
rect 21085 17215 21143 17221
rect 22094 17212 22100 17224
rect 22152 17212 22158 17264
rect 22278 17212 22284 17264
rect 22336 17252 22342 17264
rect 23934 17252 23940 17264
rect 22336 17224 23940 17252
rect 22336 17212 22342 17224
rect 23934 17212 23940 17224
rect 23992 17212 23998 17264
rect 22738 17184 22744 17196
rect 21376 17156 21680 17184
rect 20990 17116 20996 17128
rect 20916 17088 20996 17116
rect 20438 17008 20444 17060
rect 20496 17048 20502 17060
rect 20533 17051 20591 17057
rect 20533 17048 20545 17051
rect 20496 17020 20545 17048
rect 20496 17008 20502 17020
rect 20533 17017 20545 17020
rect 20579 17017 20591 17051
rect 20640 17048 20668 17081
rect 20717 17079 20775 17085
rect 20990 17076 20996 17088
rect 21048 17116 21054 17128
rect 21376 17116 21404 17156
rect 21652 17128 21680 17156
rect 21744 17156 22744 17184
rect 21048 17088 21404 17116
rect 21048 17076 21054 17088
rect 21450 17076 21456 17128
rect 21508 17076 21514 17128
rect 21634 17076 21640 17128
rect 21692 17076 21698 17128
rect 21744 17125 21772 17156
rect 22738 17144 22744 17156
rect 22796 17144 22802 17196
rect 21729 17119 21787 17125
rect 21729 17085 21741 17119
rect 21775 17085 21787 17119
rect 21729 17079 21787 17085
rect 22002 17076 22008 17128
rect 22060 17076 22066 17128
rect 22097 17119 22155 17125
rect 22097 17085 22109 17119
rect 22143 17085 22155 17119
rect 22097 17079 22155 17085
rect 21082 17048 21088 17060
rect 20640 17020 21088 17048
rect 20533 17011 20591 17017
rect 21082 17008 21088 17020
rect 21140 17048 21146 17060
rect 22103 17048 22131 17079
rect 22370 17076 22376 17128
rect 22428 17076 22434 17128
rect 22465 17119 22523 17125
rect 22465 17085 22477 17119
rect 22511 17116 22523 17119
rect 22649 17119 22707 17125
rect 22649 17116 22661 17119
rect 22511 17088 22661 17116
rect 22511 17085 22523 17088
rect 22465 17079 22523 17085
rect 22649 17085 22661 17088
rect 22695 17085 22707 17119
rect 22649 17079 22707 17085
rect 23109 17119 23167 17125
rect 23109 17085 23121 17119
rect 23155 17116 23167 17119
rect 24946 17116 24952 17128
rect 23155 17088 24952 17116
rect 23155 17085 23167 17088
rect 23109 17079 23167 17085
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 25130 17048 25136 17060
rect 21140 17020 22131 17048
rect 22940 17020 25136 17048
rect 21140 17008 21146 17020
rect 21928 16992 21956 17020
rect 11333 16983 11391 16989
rect 11333 16980 11345 16983
rect 11072 16952 11345 16980
rect 11333 16949 11345 16952
rect 11379 16949 11391 16983
rect 11333 16943 11391 16949
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 11885 16983 11943 16989
rect 11885 16980 11897 16983
rect 11572 16952 11897 16980
rect 11572 16940 11578 16952
rect 11885 16949 11897 16952
rect 11931 16949 11943 16983
rect 11885 16943 11943 16949
rect 12526 16940 12532 16992
rect 12584 16940 12590 16992
rect 13722 16940 13728 16992
rect 13780 16940 13786 16992
rect 13906 16940 13912 16992
rect 13964 16940 13970 16992
rect 14918 16940 14924 16992
rect 14976 16940 14982 16992
rect 19242 16940 19248 16992
rect 19300 16940 19306 16992
rect 20806 16940 20812 16992
rect 20864 16940 20870 16992
rect 21634 16940 21640 16992
rect 21692 16940 21698 16992
rect 21910 16940 21916 16992
rect 21968 16940 21974 16992
rect 22189 16983 22247 16989
rect 22189 16949 22201 16983
rect 22235 16980 22247 16983
rect 22646 16980 22652 16992
rect 22235 16952 22652 16980
rect 22235 16949 22247 16952
rect 22189 16943 22247 16949
rect 22646 16940 22652 16952
rect 22704 16940 22710 16992
rect 22741 16983 22799 16989
rect 22741 16949 22753 16983
rect 22787 16980 22799 16983
rect 22940 16980 22968 17020
rect 25130 17008 25136 17020
rect 25188 17008 25194 17060
rect 22787 16952 22968 16980
rect 22787 16949 22799 16952
rect 22741 16943 22799 16949
rect 23014 16940 23020 16992
rect 23072 16940 23078 16992
rect 552 16890 31531 16912
rect 552 16838 8102 16890
rect 8154 16838 8166 16890
rect 8218 16838 8230 16890
rect 8282 16838 8294 16890
rect 8346 16838 8358 16890
rect 8410 16838 15807 16890
rect 15859 16838 15871 16890
rect 15923 16838 15935 16890
rect 15987 16838 15999 16890
rect 16051 16838 16063 16890
rect 16115 16838 23512 16890
rect 23564 16838 23576 16890
rect 23628 16838 23640 16890
rect 23692 16838 23704 16890
rect 23756 16838 23768 16890
rect 23820 16838 31217 16890
rect 31269 16838 31281 16890
rect 31333 16838 31345 16890
rect 31397 16838 31409 16890
rect 31461 16838 31473 16890
rect 31525 16838 31531 16890
rect 552 16816 31531 16838
rect 7926 16736 7932 16788
rect 7984 16776 7990 16788
rect 10689 16779 10747 16785
rect 10689 16776 10701 16779
rect 7984 16748 10701 16776
rect 7984 16736 7990 16748
rect 10689 16745 10701 16748
rect 10735 16745 10747 16779
rect 10689 16739 10747 16745
rect 10796 16748 12020 16776
rect 8754 16668 8760 16720
rect 8812 16708 8818 16720
rect 10413 16711 10471 16717
rect 10413 16708 10425 16711
rect 8812 16680 10425 16708
rect 8812 16668 8818 16680
rect 10413 16677 10425 16680
rect 10459 16677 10471 16711
rect 10796 16708 10824 16748
rect 10413 16671 10471 16677
rect 10520 16680 10824 16708
rect 10520 16649 10548 16680
rect 10704 16652 10732 16680
rect 10870 16668 10876 16720
rect 10928 16708 10934 16720
rect 11885 16711 11943 16717
rect 11885 16708 11897 16711
rect 10928 16680 11897 16708
rect 10928 16668 10934 16680
rect 11885 16677 11897 16680
rect 11931 16677 11943 16711
rect 11885 16671 11943 16677
rect 11992 16708 12020 16748
rect 12618 16736 12624 16788
rect 12676 16776 12682 16788
rect 12676 16748 13216 16776
rect 12676 16736 12682 16748
rect 13188 16708 13216 16748
rect 13814 16736 13820 16788
rect 13872 16736 13878 16788
rect 13998 16736 14004 16788
rect 14056 16736 14062 16788
rect 14918 16736 14924 16788
rect 14976 16776 14982 16788
rect 21358 16776 21364 16788
rect 14976 16748 15240 16776
rect 14976 16736 14982 16748
rect 14016 16708 14044 16736
rect 15013 16711 15071 16717
rect 15013 16708 15025 16711
rect 11992 16680 12756 16708
rect 10137 16643 10195 16649
rect 10137 16609 10149 16643
rect 10183 16609 10195 16643
rect 10137 16603 10195 16609
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16609 10563 16643
rect 10505 16603 10563 16609
rect 10597 16643 10655 16649
rect 10597 16609 10609 16643
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 10042 16532 10048 16584
rect 10100 16532 10106 16584
rect 10152 16572 10180 16603
rect 10612 16572 10640 16603
rect 10686 16600 10692 16652
rect 10744 16600 10750 16652
rect 10962 16600 10968 16652
rect 11020 16600 11026 16652
rect 11054 16600 11060 16652
rect 11112 16600 11118 16652
rect 11238 16600 11244 16652
rect 11296 16600 11302 16652
rect 11330 16600 11336 16652
rect 11388 16600 11394 16652
rect 11992 16649 12020 16680
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16609 11575 16643
rect 11517 16603 11575 16609
rect 11977 16643 12035 16649
rect 11977 16609 11989 16643
rect 12023 16609 12035 16643
rect 11977 16603 12035 16609
rect 11532 16572 11560 16603
rect 12066 16600 12072 16652
rect 12124 16640 12130 16652
rect 12253 16643 12311 16649
rect 12253 16640 12265 16643
rect 12124 16612 12265 16640
rect 12124 16600 12130 16612
rect 12253 16609 12265 16612
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 12342 16600 12348 16652
rect 12400 16600 12406 16652
rect 12434 16600 12440 16652
rect 12492 16600 12498 16652
rect 12728 16649 12756 16680
rect 13188 16680 14044 16708
rect 14844 16680 15025 16708
rect 13188 16649 13216 16680
rect 12713 16643 12771 16649
rect 12713 16609 12725 16643
rect 12759 16609 12771 16643
rect 12713 16603 12771 16609
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16609 13231 16643
rect 13449 16643 13507 16649
rect 13449 16640 13461 16643
rect 13173 16603 13231 16609
rect 13372 16612 13461 16640
rect 10152 16544 10640 16572
rect 10704 16544 11560 16572
rect 10520 16516 10548 16544
rect 10502 16464 10508 16516
rect 10560 16464 10566 16516
rect 10594 16464 10600 16516
rect 10652 16504 10658 16516
rect 10704 16504 10732 16544
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 12452 16572 12480 16600
rect 13372 16572 13400 16612
rect 13449 16609 13461 16612
rect 13495 16640 13507 16643
rect 13722 16640 13728 16652
rect 13495 16612 13728 16640
rect 13495 16609 13507 16612
rect 13449 16603 13507 16609
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 14001 16643 14059 16649
rect 14001 16609 14013 16643
rect 14047 16609 14059 16643
rect 14001 16603 14059 16609
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16640 14151 16643
rect 14277 16643 14335 16649
rect 14277 16640 14289 16643
rect 14139 16612 14289 16640
rect 14139 16609 14151 16612
rect 14093 16603 14151 16609
rect 14277 16609 14289 16612
rect 14323 16609 14335 16643
rect 14277 16603 14335 16609
rect 14016 16572 14044 16603
rect 14642 16600 14648 16652
rect 14700 16640 14706 16652
rect 14844 16649 14872 16680
rect 15013 16677 15025 16680
rect 15059 16677 15071 16711
rect 15013 16671 15071 16677
rect 14737 16643 14795 16649
rect 14737 16640 14749 16643
rect 14700 16612 14749 16640
rect 14700 16600 14706 16612
rect 14737 16609 14749 16612
rect 14783 16609 14795 16643
rect 14737 16603 14795 16609
rect 14829 16643 14887 16649
rect 14829 16609 14841 16643
rect 14875 16609 14887 16643
rect 14829 16603 14887 16609
rect 14918 16600 14924 16652
rect 14976 16600 14982 16652
rect 15212 16649 15240 16748
rect 20364 16748 21364 16776
rect 15562 16668 15568 16720
rect 15620 16708 15626 16720
rect 15841 16711 15899 16717
rect 15841 16708 15853 16711
rect 15620 16680 15853 16708
rect 15620 16668 15626 16680
rect 15841 16677 15853 16680
rect 15887 16677 15899 16711
rect 15841 16671 15899 16677
rect 18877 16711 18935 16717
rect 18877 16677 18889 16711
rect 18923 16708 18935 16711
rect 20254 16708 20260 16720
rect 18923 16680 20260 16708
rect 18923 16677 18935 16680
rect 18877 16671 18935 16677
rect 20254 16668 20260 16680
rect 20312 16668 20318 16720
rect 15197 16643 15255 16649
rect 15197 16609 15209 16643
rect 15243 16609 15255 16643
rect 15197 16603 15255 16609
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16640 15715 16643
rect 15746 16640 15752 16652
rect 15703 16612 15752 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16209 16643 16267 16649
rect 16209 16640 16221 16643
rect 15979 16612 16221 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16209 16609 16221 16612
rect 16255 16609 16267 16643
rect 16209 16603 16267 16609
rect 16301 16643 16359 16649
rect 16301 16609 16313 16643
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 18969 16643 19027 16649
rect 18969 16609 18981 16643
rect 19015 16640 19027 16643
rect 19015 16612 19196 16640
rect 19015 16609 19027 16612
rect 18969 16603 19027 16609
rect 16114 16572 16120 16584
rect 11756 16544 12480 16572
rect 13188 16544 13400 16572
rect 13464 16544 16120 16572
rect 11756 16532 11762 16544
rect 10652 16476 10732 16504
rect 10652 16464 10658 16476
rect 10962 16464 10968 16516
rect 11020 16504 11026 16516
rect 11609 16507 11667 16513
rect 11609 16504 11621 16507
rect 11020 16476 11621 16504
rect 11020 16464 11026 16476
rect 11609 16473 11621 16476
rect 11655 16473 11667 16507
rect 11609 16467 11667 16473
rect 13188 16448 13216 16544
rect 13464 16448 13492 16544
rect 16114 16532 16120 16544
rect 16172 16572 16178 16584
rect 16316 16572 16344 16603
rect 16850 16572 16856 16584
rect 16172 16544 16856 16572
rect 16172 16532 16178 16544
rect 16850 16532 16856 16544
rect 16908 16532 16914 16584
rect 19168 16572 19196 16612
rect 19242 16600 19248 16652
rect 19300 16600 19306 16652
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 19518 16640 19524 16652
rect 19392 16612 19524 16640
rect 19392 16600 19398 16612
rect 19518 16600 19524 16612
rect 19576 16600 19582 16652
rect 19613 16643 19671 16649
rect 19613 16609 19625 16643
rect 19659 16609 19671 16643
rect 19613 16603 19671 16609
rect 20073 16643 20131 16649
rect 20073 16609 20085 16643
rect 20119 16640 20131 16643
rect 20364 16640 20392 16748
rect 21358 16736 21364 16748
rect 21416 16736 21422 16788
rect 21450 16736 21456 16788
rect 21508 16776 21514 16788
rect 22465 16779 22523 16785
rect 22465 16776 22477 16779
rect 21508 16748 22477 16776
rect 21508 16736 21514 16748
rect 22465 16745 22477 16748
rect 22511 16745 22523 16779
rect 22465 16739 22523 16745
rect 22646 16736 22652 16788
rect 22704 16736 22710 16788
rect 22738 16736 22744 16788
rect 22796 16736 22802 16788
rect 22830 16736 22836 16788
rect 22888 16776 22894 16788
rect 23017 16779 23075 16785
rect 23017 16776 23029 16779
rect 22888 16748 23029 16776
rect 22888 16736 22894 16748
rect 23017 16745 23029 16748
rect 23063 16745 23075 16779
rect 23017 16739 23075 16745
rect 23106 16736 23112 16788
rect 23164 16776 23170 16788
rect 23569 16779 23627 16785
rect 23569 16776 23581 16779
rect 23164 16748 23581 16776
rect 23164 16736 23170 16748
rect 23569 16745 23581 16748
rect 23615 16745 23627 16779
rect 23569 16739 23627 16745
rect 20625 16711 20683 16717
rect 20625 16677 20637 16711
rect 20671 16708 20683 16711
rect 20898 16708 20904 16720
rect 20671 16680 20904 16708
rect 20671 16677 20683 16680
rect 20625 16671 20683 16677
rect 20898 16668 20904 16680
rect 20956 16668 20962 16720
rect 21082 16708 21088 16720
rect 21008 16680 21088 16708
rect 21008 16649 21036 16680
rect 21082 16668 21088 16680
rect 21140 16668 21146 16720
rect 21266 16668 21272 16720
rect 21324 16708 21330 16720
rect 22189 16711 22247 16717
rect 22189 16708 22201 16711
rect 21324 16680 22201 16708
rect 21324 16668 21330 16680
rect 22189 16677 22201 16680
rect 22235 16677 22247 16711
rect 22664 16708 22692 16736
rect 22664 16680 23244 16708
rect 22189 16671 22247 16677
rect 20119 16612 20392 16640
rect 20441 16643 20499 16649
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 20441 16609 20453 16643
rect 20487 16640 20499 16643
rect 20717 16643 20775 16649
rect 20487 16612 20576 16640
rect 20487 16609 20499 16612
rect 20441 16603 20499 16609
rect 19628 16572 19656 16603
rect 19168 16544 20208 16572
rect 13722 16464 13728 16516
rect 13780 16504 13786 16516
rect 14369 16507 14427 16513
rect 14369 16504 14381 16507
rect 13780 16476 14381 16504
rect 13780 16464 13786 16476
rect 14369 16473 14381 16476
rect 14415 16504 14427 16507
rect 14458 16504 14464 16516
rect 14415 16476 14464 16504
rect 14415 16473 14427 16476
rect 14369 16467 14427 16473
rect 14458 16464 14464 16476
rect 14516 16464 14522 16516
rect 15010 16464 15016 16516
rect 15068 16504 15074 16516
rect 15565 16507 15623 16513
rect 15565 16504 15577 16507
rect 15068 16476 15577 16504
rect 15068 16464 15074 16476
rect 15565 16473 15577 16476
rect 15611 16473 15623 16507
rect 15565 16467 15623 16473
rect 19153 16507 19211 16513
rect 19153 16473 19165 16507
rect 19199 16504 19211 16507
rect 19199 16476 20116 16504
rect 19199 16473 19211 16476
rect 19153 16467 19211 16473
rect 11422 16396 11428 16448
rect 11480 16436 11486 16448
rect 12161 16439 12219 16445
rect 12161 16436 12173 16439
rect 11480 16408 12173 16436
rect 11480 16396 11486 16408
rect 12161 16405 12173 16408
rect 12207 16405 12219 16439
rect 12161 16399 12219 16405
rect 12434 16396 12440 16448
rect 12492 16396 12498 16448
rect 12802 16396 12808 16448
rect 12860 16396 12866 16448
rect 13078 16396 13084 16448
rect 13136 16396 13142 16448
rect 13170 16396 13176 16448
rect 13228 16396 13234 16448
rect 13354 16396 13360 16448
rect 13412 16396 13418 16448
rect 13446 16396 13452 16448
rect 13504 16396 13510 16448
rect 14476 16436 14504 16464
rect 20088 16448 20116 16476
rect 14918 16436 14924 16448
rect 14476 16408 14924 16436
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 15194 16396 15200 16448
rect 15252 16436 15258 16448
rect 15289 16439 15347 16445
rect 15289 16436 15301 16439
rect 15252 16408 15301 16436
rect 15252 16396 15258 16408
rect 15289 16405 15301 16408
rect 15335 16405 15347 16439
rect 15289 16399 15347 16405
rect 19426 16396 19432 16448
rect 19484 16396 19490 16448
rect 19518 16396 19524 16448
rect 19576 16436 19582 16448
rect 19705 16439 19763 16445
rect 19705 16436 19717 16439
rect 19576 16408 19717 16436
rect 19576 16396 19582 16408
rect 19705 16405 19717 16408
rect 19751 16405 19763 16439
rect 19705 16399 19763 16405
rect 19978 16396 19984 16448
rect 20036 16396 20042 16448
rect 20070 16396 20076 16448
rect 20128 16396 20134 16448
rect 20180 16436 20208 16544
rect 20346 16532 20352 16584
rect 20404 16532 20410 16584
rect 20548 16504 20576 16612
rect 20717 16609 20729 16643
rect 20763 16640 20775 16643
rect 20993 16643 21051 16649
rect 20763 16612 20944 16640
rect 20763 16609 20775 16612
rect 20717 16603 20775 16609
rect 20916 16504 20944 16612
rect 20993 16609 21005 16643
rect 21039 16609 21051 16643
rect 20993 16603 21051 16609
rect 21450 16600 21456 16652
rect 21508 16600 21514 16652
rect 21545 16643 21603 16649
rect 21545 16609 21557 16643
rect 21591 16609 21603 16643
rect 21545 16603 21603 16609
rect 21266 16532 21272 16584
rect 21324 16572 21330 16584
rect 21560 16572 21588 16603
rect 21726 16600 21732 16652
rect 21784 16640 21790 16652
rect 21913 16643 21971 16649
rect 21913 16640 21925 16643
rect 21784 16612 21925 16640
rect 21784 16600 21790 16612
rect 21913 16609 21925 16612
rect 21959 16609 21971 16643
rect 21913 16603 21971 16609
rect 22002 16600 22008 16652
rect 22060 16600 22066 16652
rect 22278 16600 22284 16652
rect 22336 16600 22342 16652
rect 23216 16649 23244 16680
rect 23290 16668 23296 16720
rect 23348 16668 23354 16720
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16609 22615 16643
rect 22557 16603 22615 16609
rect 22833 16643 22891 16649
rect 22833 16609 22845 16643
rect 22879 16640 22891 16643
rect 23109 16643 23167 16649
rect 22879 16612 23060 16640
rect 22879 16609 22891 16612
rect 22833 16603 22891 16609
rect 21324 16544 21588 16572
rect 22572 16572 22600 16603
rect 22738 16572 22744 16584
rect 22572 16544 22744 16572
rect 21324 16532 21330 16544
rect 22738 16532 22744 16544
rect 22796 16532 22802 16584
rect 23032 16504 23060 16612
rect 23109 16609 23121 16643
rect 23155 16609 23167 16643
rect 23109 16603 23167 16609
rect 23201 16643 23259 16649
rect 23201 16609 23213 16643
rect 23247 16609 23259 16643
rect 23201 16603 23259 16609
rect 23124 16572 23152 16603
rect 23658 16600 23664 16652
rect 23716 16600 23722 16652
rect 23750 16572 23756 16584
rect 23124 16544 23756 16572
rect 23750 16532 23756 16544
rect 23808 16532 23814 16584
rect 24302 16504 24308 16516
rect 20548 16476 20752 16504
rect 20916 16476 24308 16504
rect 20530 16436 20536 16448
rect 20180 16408 20536 16436
rect 20530 16396 20536 16408
rect 20588 16396 20594 16448
rect 20724 16436 20752 16476
rect 24302 16464 24308 16476
rect 24360 16464 24366 16516
rect 20901 16439 20959 16445
rect 20901 16436 20913 16439
rect 20724 16408 20913 16436
rect 20901 16405 20913 16408
rect 20947 16405 20959 16439
rect 20901 16399 20959 16405
rect 21174 16396 21180 16448
rect 21232 16436 21238 16448
rect 21361 16439 21419 16445
rect 21361 16436 21373 16439
rect 21232 16408 21373 16436
rect 21232 16396 21238 16408
rect 21361 16405 21373 16408
rect 21407 16405 21419 16439
rect 21361 16399 21419 16405
rect 21637 16439 21695 16445
rect 21637 16405 21649 16439
rect 21683 16436 21695 16439
rect 22462 16436 22468 16448
rect 21683 16408 22468 16436
rect 21683 16405 21695 16408
rect 21637 16399 21695 16405
rect 22462 16396 22468 16408
rect 22520 16396 22526 16448
rect 23566 16396 23572 16448
rect 23624 16436 23630 16448
rect 24578 16436 24584 16448
rect 23624 16408 24584 16436
rect 23624 16396 23630 16408
rect 24578 16396 24584 16408
rect 24636 16396 24642 16448
rect 552 16346 31372 16368
rect 552 16294 4250 16346
rect 4302 16294 4314 16346
rect 4366 16294 4378 16346
rect 4430 16294 4442 16346
rect 4494 16294 4506 16346
rect 4558 16294 11955 16346
rect 12007 16294 12019 16346
rect 12071 16294 12083 16346
rect 12135 16294 12147 16346
rect 12199 16294 12211 16346
rect 12263 16294 19660 16346
rect 19712 16294 19724 16346
rect 19776 16294 19788 16346
rect 19840 16294 19852 16346
rect 19904 16294 19916 16346
rect 19968 16294 27365 16346
rect 27417 16294 27429 16346
rect 27481 16294 27493 16346
rect 27545 16294 27557 16346
rect 27609 16294 27621 16346
rect 27673 16294 31372 16346
rect 552 16272 31372 16294
rect 7466 16192 7472 16244
rect 7524 16232 7530 16244
rect 7524 16204 10548 16232
rect 7524 16192 7530 16204
rect 9766 16124 9772 16176
rect 9824 16124 9830 16176
rect 9858 16124 9864 16176
rect 9916 16164 9922 16176
rect 10413 16167 10471 16173
rect 10413 16164 10425 16167
rect 9916 16136 10425 16164
rect 9916 16124 9922 16136
rect 10413 16133 10425 16136
rect 10459 16133 10471 16167
rect 10520 16164 10548 16204
rect 10962 16192 10968 16244
rect 11020 16192 11026 16244
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11793 16235 11851 16241
rect 11112 16204 11284 16232
rect 11112 16192 11118 16204
rect 11256 16164 11284 16204
rect 11793 16201 11805 16235
rect 11839 16232 11851 16235
rect 12342 16232 12348 16244
rect 11839 16204 12348 16232
rect 11839 16201 11851 16204
rect 11793 16195 11851 16201
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 12618 16192 12624 16244
rect 12676 16192 12682 16244
rect 12989 16235 13047 16241
rect 12989 16201 13001 16235
rect 13035 16232 13047 16235
rect 13906 16232 13912 16244
rect 13035 16204 13912 16232
rect 13035 16201 13047 16204
rect 12989 16195 13047 16201
rect 13906 16192 13912 16204
rect 13964 16192 13970 16244
rect 13998 16192 14004 16244
rect 14056 16192 14062 16244
rect 14550 16192 14556 16244
rect 14608 16232 14614 16244
rect 15105 16235 15163 16241
rect 15105 16232 15117 16235
rect 14608 16204 15117 16232
rect 14608 16192 14614 16204
rect 15105 16201 15117 16204
rect 15151 16201 15163 16235
rect 15105 16195 15163 16201
rect 15746 16192 15752 16244
rect 15804 16232 15810 16244
rect 18230 16232 18236 16244
rect 15804 16204 18236 16232
rect 15804 16192 15810 16204
rect 10520 16136 11192 16164
rect 11256 16136 11836 16164
rect 10413 16127 10471 16133
rect 9784 16096 9812 16124
rect 9692 16068 9812 16096
rect 10244 16068 10732 16096
rect 9692 16037 9720 16068
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 9766 15988 9772 16040
rect 9824 15988 9830 16040
rect 10134 16028 10140 16040
rect 10069 16000 10140 16028
rect 9585 15963 9643 15969
rect 9585 15929 9597 15963
rect 9631 15960 9643 15963
rect 10069 15960 10097 16000
rect 10134 15988 10140 16000
rect 10192 15988 10198 16040
rect 10244 16037 10272 16068
rect 10704 16040 10732 16068
rect 10229 16031 10287 16037
rect 10229 15997 10241 16031
rect 10275 15997 10287 16031
rect 10229 15991 10287 15997
rect 10329 16025 10387 16031
rect 10329 15991 10341 16025
rect 10375 15991 10387 16025
rect 10329 15985 10387 15991
rect 10502 15988 10508 16040
rect 10560 16028 10566 16040
rect 10597 16031 10655 16037
rect 10597 16028 10609 16031
rect 10560 16000 10609 16028
rect 10560 15988 10566 16000
rect 10597 15997 10609 16000
rect 10643 15997 10655 16031
rect 10597 15991 10655 15997
rect 9631 15932 10097 15960
rect 9631 15929 9643 15932
rect 9585 15923 9643 15929
rect 10336 15904 10364 15985
rect 10612 15960 10640 15991
rect 10686 15988 10692 16040
rect 10744 15988 10750 16040
rect 10873 16031 10931 16037
rect 10873 15997 10885 16031
rect 10919 16030 10931 16031
rect 10962 16030 10968 16040
rect 10919 16002 10968 16030
rect 10919 15997 10931 16002
rect 10873 15991 10931 15997
rect 10962 15988 10968 16002
rect 11020 15988 11026 16040
rect 11164 16037 11192 16136
rect 11514 16056 11520 16108
rect 11572 16096 11578 16108
rect 11808 16096 11836 16136
rect 11882 16124 11888 16176
rect 11940 16164 11946 16176
rect 12636 16164 12664 16192
rect 11940 16136 12664 16164
rect 11940 16124 11946 16136
rect 14826 16124 14832 16176
rect 14884 16164 14890 16176
rect 16298 16164 16304 16176
rect 14884 16136 16304 16164
rect 14884 16124 14890 16136
rect 16298 16124 16304 16136
rect 16356 16124 16362 16176
rect 12434 16096 12440 16108
rect 11572 16068 11744 16096
rect 11808 16068 12440 16096
rect 11572 16056 11578 16068
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 15997 11207 16031
rect 11149 15991 11207 15997
rect 11238 15988 11244 16040
rect 11296 16028 11302 16040
rect 11716 16037 11744 16068
rect 11992 16037 12020 16068
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 15580 16068 16344 16096
rect 11609 16031 11667 16037
rect 11609 16028 11621 16031
rect 11296 16000 11621 16028
rect 11296 15988 11302 16000
rect 11609 15997 11621 16000
rect 11655 15997 11667 16031
rect 11609 15991 11667 15997
rect 11701 16031 11759 16037
rect 11701 15997 11713 16031
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 12069 16031 12127 16037
rect 12069 15997 12081 16031
rect 12115 16028 12127 16031
rect 12253 16031 12311 16037
rect 12253 16028 12265 16031
rect 12115 16000 12265 16028
rect 12115 15997 12127 16000
rect 12069 15991 12127 15997
rect 12253 15997 12265 16000
rect 12299 15997 12311 16031
rect 12253 15991 12311 15997
rect 11624 15960 11652 15991
rect 12618 15988 12624 16040
rect 12676 15988 12682 16040
rect 12802 15988 12808 16040
rect 12860 15988 12866 16040
rect 13078 15988 13084 16040
rect 13136 15988 13142 16040
rect 13354 15988 13360 16040
rect 13412 15988 13418 16040
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 15997 13691 16031
rect 13633 15991 13691 15997
rect 13725 16031 13783 16037
rect 13725 15997 13737 16031
rect 13771 16028 13783 16031
rect 13909 16031 13967 16037
rect 13909 16028 13921 16031
rect 13771 16000 13921 16028
rect 13771 15997 13783 16000
rect 13725 15991 13783 15997
rect 13909 15997 13921 16000
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 14369 16031 14427 16037
rect 14369 15997 14381 16031
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 13265 15963 13323 15969
rect 13265 15960 13277 15963
rect 10612 15932 11008 15960
rect 11624 15932 13277 15960
rect 10980 15904 11008 15932
rect 13265 15929 13277 15932
rect 13311 15929 13323 15963
rect 13265 15923 13323 15929
rect 8018 15852 8024 15904
rect 8076 15892 8082 15904
rect 9861 15895 9919 15901
rect 9861 15892 9873 15895
rect 8076 15864 9873 15892
rect 8076 15852 8082 15864
rect 9861 15861 9873 15864
rect 9907 15861 9919 15895
rect 9861 15855 9919 15861
rect 10134 15852 10140 15904
rect 10192 15852 10198 15904
rect 10318 15852 10324 15904
rect 10376 15852 10382 15904
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 10689 15895 10747 15901
rect 10689 15892 10701 15895
rect 10560 15864 10701 15892
rect 10560 15852 10566 15864
rect 10689 15861 10701 15864
rect 10735 15861 10747 15895
rect 10689 15855 10747 15861
rect 10962 15852 10968 15904
rect 11020 15852 11026 15904
rect 11146 15852 11152 15904
rect 11204 15892 11210 15904
rect 11241 15895 11299 15901
rect 11241 15892 11253 15895
rect 11204 15864 11253 15892
rect 11204 15852 11210 15864
rect 11241 15861 11253 15864
rect 11287 15861 11299 15895
rect 11241 15855 11299 15861
rect 11514 15852 11520 15904
rect 11572 15852 11578 15904
rect 12342 15852 12348 15904
rect 12400 15852 12406 15904
rect 12710 15852 12716 15904
rect 12768 15852 12774 15904
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 13648 15892 13676 15991
rect 13814 15920 13820 15972
rect 13872 15960 13878 15972
rect 14277 15963 14335 15969
rect 14277 15960 14289 15963
rect 13872 15932 14289 15960
rect 13872 15920 13878 15932
rect 14277 15929 14289 15932
rect 14323 15929 14335 15963
rect 14277 15923 14335 15929
rect 14384 15960 14412 15991
rect 14458 15988 14464 16040
rect 14516 15988 14522 16040
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 16028 14611 16031
rect 14737 16031 14795 16037
rect 14737 16028 14749 16031
rect 14599 16000 14749 16028
rect 14599 15997 14611 16000
rect 14553 15991 14611 15997
rect 14737 15997 14749 16000
rect 14783 15997 14795 16031
rect 14737 15991 14795 15997
rect 15197 16031 15255 16037
rect 15197 15997 15209 16031
rect 15243 15997 15255 16031
rect 15197 15991 15255 15997
rect 15212 15960 15240 15991
rect 15286 15988 15292 16040
rect 15344 16028 15350 16040
rect 15580 16037 15608 16068
rect 15565 16031 15623 16037
rect 15565 16028 15577 16031
rect 15344 16000 15577 16028
rect 15344 15988 15350 16000
rect 15565 15997 15577 16000
rect 15611 15997 15623 16031
rect 15565 15991 15623 15997
rect 15654 15988 15660 16040
rect 15712 16028 15718 16040
rect 15749 16031 15807 16037
rect 15749 16028 15761 16031
rect 15712 16000 15761 16028
rect 15712 15988 15718 16000
rect 15749 15997 15761 16000
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 15933 16031 15991 16037
rect 15933 15997 15945 16031
rect 15979 15997 15991 16031
rect 15933 15991 15991 15997
rect 14384 15932 15240 15960
rect 15948 15960 15976 15991
rect 16114 15988 16120 16040
rect 16172 16028 16178 16040
rect 16316 16037 16344 16068
rect 16209 16031 16267 16037
rect 16209 16028 16221 16031
rect 16172 16000 16221 16028
rect 16172 15988 16178 16000
rect 16209 15997 16221 16000
rect 16255 15997 16267 16031
rect 16209 15991 16267 15997
rect 16301 16031 16359 16037
rect 16301 15997 16313 16031
rect 16347 15997 16359 16031
rect 16500 16028 16528 16204
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 19518 16192 19524 16244
rect 19576 16232 19582 16244
rect 19889 16235 19947 16241
rect 19889 16232 19901 16235
rect 19576 16204 19901 16232
rect 19576 16192 19582 16204
rect 19889 16201 19901 16204
rect 19935 16201 19947 16235
rect 19889 16195 19947 16201
rect 20254 16192 20260 16244
rect 20312 16192 20318 16244
rect 20806 16192 20812 16244
rect 20864 16192 20870 16244
rect 20898 16192 20904 16244
rect 20956 16232 20962 16244
rect 20993 16235 21051 16241
rect 20993 16232 21005 16235
rect 20956 16204 21005 16232
rect 20956 16192 20962 16204
rect 20993 16201 21005 16204
rect 21039 16201 21051 16235
rect 20993 16195 21051 16201
rect 21269 16235 21327 16241
rect 21269 16201 21281 16235
rect 21315 16232 21327 16235
rect 21358 16232 21364 16244
rect 21315 16204 21364 16232
rect 21315 16201 21327 16204
rect 21269 16195 21327 16201
rect 21358 16192 21364 16204
rect 21416 16192 21422 16244
rect 22094 16192 22100 16244
rect 22152 16192 22158 16244
rect 22462 16192 22468 16244
rect 22520 16232 22526 16244
rect 23201 16235 23259 16241
rect 22520 16204 22968 16232
rect 22520 16192 22526 16204
rect 18141 16167 18199 16173
rect 18141 16133 18153 16167
rect 18187 16164 18199 16167
rect 19794 16164 19800 16176
rect 18187 16136 19800 16164
rect 18187 16133 18199 16136
rect 18141 16127 18199 16133
rect 19794 16124 19800 16136
rect 19852 16124 19858 16176
rect 18782 16056 18788 16108
rect 18840 16056 18846 16108
rect 19610 16056 19616 16108
rect 19668 16096 19674 16108
rect 20272 16096 20300 16192
rect 20824 16096 20852 16192
rect 22940 16164 22968 16204
rect 23201 16201 23213 16235
rect 23247 16232 23259 16235
rect 23290 16232 23296 16244
rect 23247 16204 23296 16232
rect 23247 16201 23259 16204
rect 23201 16195 23259 16201
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 23658 16192 23664 16244
rect 23716 16232 23722 16244
rect 24489 16235 24547 16241
rect 24489 16232 24501 16235
rect 23716 16204 24501 16232
rect 23716 16192 23722 16204
rect 24489 16201 24501 16204
rect 24535 16201 24547 16235
rect 24489 16195 24547 16201
rect 23382 16164 23388 16176
rect 22940 16136 23388 16164
rect 23382 16124 23388 16136
rect 23440 16124 23446 16176
rect 24302 16164 24308 16176
rect 23860 16136 24308 16164
rect 22370 16096 22376 16108
rect 19668 16068 19840 16096
rect 20272 16068 20668 16096
rect 20824 16068 22048 16096
rect 19668 16056 19674 16068
rect 16569 16031 16627 16037
rect 16569 16028 16581 16031
rect 16500 16000 16581 16028
rect 16301 15991 16359 15997
rect 16569 15997 16581 16000
rect 16615 15997 16627 16031
rect 16569 15991 16627 15997
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 16028 17279 16031
rect 17405 16031 17463 16037
rect 17405 16028 17417 16031
rect 17267 16000 17417 16028
rect 17267 15997 17279 16000
rect 17221 15991 17279 15997
rect 17405 15997 17417 16000
rect 17451 15997 17463 16031
rect 17405 15991 17463 15997
rect 17497 16031 17555 16037
rect 17497 15997 17509 16031
rect 17543 16028 17555 16031
rect 17954 16028 17960 16040
rect 17543 16000 17960 16028
rect 17543 15997 17555 16000
rect 17497 15991 17555 15997
rect 17954 15988 17960 16000
rect 18012 15988 18018 16040
rect 18233 16033 18291 16039
rect 18233 15999 18245 16033
rect 18279 15999 18291 16033
rect 18233 15993 18291 15999
rect 16393 15963 16451 15969
rect 16393 15960 16405 15963
rect 15948 15932 16405 15960
rect 14384 15892 14412 15932
rect 14752 15904 14780 15932
rect 16393 15929 16405 15932
rect 16439 15929 16451 15963
rect 18248 15960 18276 15993
rect 18322 15988 18328 16040
rect 18380 15988 18386 16040
rect 18800 16028 18828 16056
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 18800 16000 18889 16028
rect 18877 15997 18889 16000
rect 18923 15997 18935 16031
rect 18877 15991 18935 15997
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 16028 19027 16031
rect 19015 16000 19196 16028
rect 19015 15997 19027 16000
rect 18969 15991 19027 15997
rect 18785 15963 18843 15969
rect 18785 15960 18797 15963
rect 18248 15932 18797 15960
rect 16393 15923 16451 15929
rect 18785 15929 18797 15932
rect 18831 15929 18843 15963
rect 18785 15923 18843 15929
rect 19168 15904 19196 16000
rect 19426 15988 19432 16040
rect 19484 15988 19490 16040
rect 19812 16037 19840 16068
rect 19705 16031 19763 16037
rect 19705 16028 19717 16031
rect 19536 16000 19717 16028
rect 12860 15864 14412 15892
rect 12860 15852 12866 15864
rect 14734 15852 14740 15904
rect 14792 15852 14798 15904
rect 14826 15852 14832 15904
rect 14884 15852 14890 15904
rect 15470 15852 15476 15904
rect 15528 15852 15534 15904
rect 15933 15895 15991 15901
rect 15933 15861 15945 15895
rect 15979 15892 15991 15895
rect 16117 15895 16175 15901
rect 16117 15892 16129 15895
rect 15979 15864 16129 15892
rect 15979 15861 15991 15864
rect 15933 15855 15991 15861
rect 16117 15861 16129 15864
rect 16163 15861 16175 15895
rect 16117 15855 16175 15861
rect 16666 15852 16672 15904
rect 16724 15852 16730 15904
rect 17126 15852 17132 15904
rect 17184 15852 17190 15904
rect 18414 15852 18420 15904
rect 18472 15852 18478 15904
rect 19058 15852 19064 15904
rect 19116 15852 19122 15904
rect 19150 15852 19156 15904
rect 19208 15852 19214 15904
rect 19337 15895 19395 15901
rect 19337 15861 19349 15895
rect 19383 15892 19395 15895
rect 19426 15892 19432 15904
rect 19383 15864 19432 15892
rect 19383 15861 19395 15864
rect 19337 15855 19395 15861
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 19536 15892 19564 16000
rect 19705 15997 19717 16000
rect 19751 15997 19763 16031
rect 19705 15991 19763 15997
rect 19797 16031 19855 16037
rect 19797 15997 19809 16031
rect 19843 15997 19855 16031
rect 19797 15991 19855 15997
rect 19978 15988 19984 16040
rect 20036 15988 20042 16040
rect 20257 16031 20315 16037
rect 20257 15997 20269 16031
rect 20303 16028 20315 16031
rect 20346 16028 20352 16040
rect 20303 16000 20352 16028
rect 20303 15997 20315 16000
rect 20257 15991 20315 15997
rect 20346 15988 20352 16000
rect 20404 15988 20410 16040
rect 20640 16037 20668 16068
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 20625 16031 20683 16037
rect 20625 15997 20637 16031
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 19613 15963 19671 15969
rect 19613 15929 19625 15963
rect 19659 15960 19671 15963
rect 20441 15963 20499 15969
rect 20441 15960 20453 15963
rect 19659 15932 20453 15960
rect 19659 15929 19671 15932
rect 19613 15923 19671 15929
rect 20441 15929 20453 15932
rect 20487 15929 20499 15963
rect 20548 15960 20576 15991
rect 20898 15988 20904 16040
rect 20956 15988 20962 16040
rect 21085 16031 21143 16037
rect 21085 15997 21097 16031
rect 21131 16028 21143 16031
rect 21174 16028 21180 16040
rect 21131 16000 21180 16028
rect 21131 15997 21143 16000
rect 21085 15991 21143 15997
rect 21174 15988 21180 16000
rect 21232 15988 21238 16040
rect 21358 15988 21364 16040
rect 21416 15988 21422 16040
rect 22020 16037 22048 16068
rect 22112 16068 22376 16096
rect 21453 16031 21511 16037
rect 21453 15997 21465 16031
rect 21499 15997 21511 16031
rect 21453 15991 21511 15997
rect 21913 16031 21971 16037
rect 21913 15997 21925 16031
rect 21959 15997 21971 16031
rect 21913 15991 21971 15997
rect 22005 16031 22063 16037
rect 22005 15997 22017 16031
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 21468 15960 21496 15991
rect 20548 15932 21128 15960
rect 20441 15923 20499 15929
rect 21100 15904 21128 15932
rect 21284 15932 21496 15960
rect 21928 15960 21956 15991
rect 22112 15960 22140 16068
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 22738 16056 22744 16108
rect 22796 16096 22802 16108
rect 23477 16099 23535 16105
rect 23477 16096 23489 16099
rect 22796 16068 23489 16096
rect 22796 16056 22802 16068
rect 23477 16065 23489 16068
rect 23523 16065 23535 16099
rect 23477 16059 23535 16065
rect 22186 15988 22192 16040
rect 22244 15988 22250 16040
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 15997 22339 16031
rect 22281 15991 22339 15997
rect 21928 15932 22140 15960
rect 22296 15960 22324 15991
rect 22462 15988 22468 16040
rect 22520 16028 22526 16040
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 22520 16000 22569 16028
rect 22520 15988 22526 16000
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 22830 15988 22836 16040
rect 22888 16028 22894 16040
rect 23017 16031 23075 16037
rect 22888 16000 22968 16028
rect 22888 15988 22894 16000
rect 22940 15960 22968 16000
rect 23017 15997 23029 16031
rect 23063 15997 23075 16031
rect 23017 15991 23075 15997
rect 22296 15932 22968 15960
rect 23032 15960 23060 15991
rect 23290 15988 23296 16040
rect 23348 15988 23354 16040
rect 23566 15988 23572 16040
rect 23624 15988 23630 16040
rect 23860 16037 23888 16136
rect 24302 16124 24308 16136
rect 24360 16124 24366 16176
rect 24026 16056 24032 16108
rect 24084 16096 24090 16108
rect 25222 16096 25228 16108
rect 24084 16068 24164 16096
rect 24084 16056 24090 16068
rect 24136 16037 24164 16068
rect 24228 16068 25228 16096
rect 23845 16031 23903 16037
rect 23845 15997 23857 16031
rect 23891 15997 23903 16031
rect 23845 15991 23903 15997
rect 24121 16031 24179 16037
rect 24121 15997 24133 16031
rect 24167 15997 24179 16031
rect 24121 15991 24179 15997
rect 23937 15963 23995 15969
rect 23032 15932 23888 15960
rect 21284 15904 21312 15932
rect 20165 15895 20223 15901
rect 20165 15892 20177 15895
rect 19536 15864 20177 15892
rect 20165 15861 20177 15864
rect 20211 15861 20223 15895
rect 20165 15855 20223 15861
rect 20254 15852 20260 15904
rect 20312 15892 20318 15904
rect 20717 15895 20775 15901
rect 20717 15892 20729 15895
rect 20312 15864 20729 15892
rect 20312 15852 20318 15864
rect 20717 15861 20729 15864
rect 20763 15861 20775 15895
rect 20717 15855 20775 15861
rect 21082 15852 21088 15904
rect 21140 15852 21146 15904
rect 21266 15852 21272 15904
rect 21324 15852 21330 15904
rect 21542 15852 21548 15904
rect 21600 15852 21606 15904
rect 21818 15852 21824 15904
rect 21876 15852 21882 15904
rect 21910 15852 21916 15904
rect 21968 15892 21974 15904
rect 22296 15892 22324 15932
rect 21968 15864 22324 15892
rect 22373 15895 22431 15901
rect 21968 15852 21974 15864
rect 22373 15861 22385 15895
rect 22419 15892 22431 15895
rect 22554 15892 22560 15904
rect 22419 15864 22560 15892
rect 22419 15861 22431 15864
rect 22373 15855 22431 15861
rect 22554 15852 22560 15864
rect 22612 15852 22618 15904
rect 22649 15895 22707 15901
rect 22649 15861 22661 15895
rect 22695 15892 22707 15895
rect 22830 15892 22836 15904
rect 22695 15864 22836 15892
rect 22695 15861 22707 15864
rect 22649 15855 22707 15861
rect 22830 15852 22836 15864
rect 22888 15852 22894 15904
rect 22940 15901 22968 15932
rect 22925 15895 22983 15901
rect 22925 15861 22937 15895
rect 22971 15861 22983 15895
rect 23860 15892 23888 15932
rect 23937 15929 23949 15963
rect 23983 15960 23995 15963
rect 24228 15960 24256 16068
rect 25222 16056 25228 16068
rect 25280 16056 25286 16108
rect 24302 15988 24308 16040
rect 24360 16028 24366 16040
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 24360 16000 24593 16028
rect 24360 15988 24366 16000
rect 24581 15997 24593 16000
rect 24627 16028 24639 16031
rect 26418 16028 26424 16040
rect 24627 16000 26424 16028
rect 24627 15997 24639 16000
rect 24581 15991 24639 15997
rect 26418 15988 26424 16000
rect 26476 15988 26482 16040
rect 23983 15932 24256 15960
rect 23983 15929 23995 15932
rect 23937 15923 23995 15929
rect 24118 15892 24124 15904
rect 23860 15864 24124 15892
rect 22925 15855 22983 15861
rect 24118 15852 24124 15864
rect 24176 15852 24182 15904
rect 24213 15895 24271 15901
rect 24213 15861 24225 15895
rect 24259 15892 24271 15895
rect 26602 15892 26608 15904
rect 24259 15864 26608 15892
rect 24259 15861 24271 15864
rect 24213 15855 24271 15861
rect 26602 15852 26608 15864
rect 26660 15852 26666 15904
rect 552 15802 31531 15824
rect 552 15750 8102 15802
rect 8154 15750 8166 15802
rect 8218 15750 8230 15802
rect 8282 15750 8294 15802
rect 8346 15750 8358 15802
rect 8410 15750 15807 15802
rect 15859 15750 15871 15802
rect 15923 15750 15935 15802
rect 15987 15750 15999 15802
rect 16051 15750 16063 15802
rect 16115 15750 23512 15802
rect 23564 15750 23576 15802
rect 23628 15750 23640 15802
rect 23692 15750 23704 15802
rect 23756 15750 23768 15802
rect 23820 15750 31217 15802
rect 31269 15750 31281 15802
rect 31333 15750 31345 15802
rect 31397 15750 31409 15802
rect 31461 15750 31473 15802
rect 31525 15750 31531 15802
rect 552 15728 31531 15750
rect 8757 15691 8815 15697
rect 8757 15657 8769 15691
rect 8803 15688 8815 15691
rect 9766 15688 9772 15700
rect 8803 15660 9772 15688
rect 8803 15657 8815 15660
rect 8757 15651 8815 15657
rect 9766 15648 9772 15660
rect 9824 15648 9830 15700
rect 9861 15691 9919 15697
rect 9861 15657 9873 15691
rect 9907 15688 9919 15691
rect 9950 15688 9956 15700
rect 9907 15660 9956 15688
rect 9907 15657 9919 15660
rect 9861 15651 9919 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10318 15688 10324 15700
rect 10152 15660 10324 15688
rect 9585 15623 9643 15629
rect 9585 15589 9597 15623
rect 9631 15620 9643 15623
rect 10152 15620 10180 15660
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 10594 15688 10600 15700
rect 10520 15660 10600 15688
rect 10520 15620 10548 15660
rect 10594 15648 10600 15660
rect 10652 15648 10658 15700
rect 10870 15648 10876 15700
rect 10928 15648 10934 15700
rect 11422 15688 11428 15700
rect 11256 15660 11428 15688
rect 10888 15620 10916 15648
rect 9631 15592 10180 15620
rect 10253 15592 10548 15620
rect 10612 15592 10916 15620
rect 9631 15589 9643 15592
rect 9585 15583 9643 15589
rect 8665 15555 8723 15561
rect 8665 15521 8677 15555
rect 8711 15521 8723 15555
rect 8665 15515 8723 15521
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 8680 15484 8708 15515
rect 8938 15512 8944 15564
rect 8996 15512 9002 15564
rect 9401 15555 9459 15561
rect 9401 15521 9413 15555
rect 9447 15552 9459 15555
rect 9490 15552 9496 15564
rect 9447 15524 9496 15552
rect 9447 15521 9459 15524
rect 9401 15515 9459 15521
rect 9490 15512 9496 15524
rect 9548 15512 9554 15564
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 9769 15555 9827 15561
rect 9769 15552 9781 15555
rect 9732 15524 9781 15552
rect 9732 15512 9738 15524
rect 9769 15521 9781 15524
rect 9815 15521 9827 15555
rect 9769 15515 9827 15521
rect 10042 15512 10048 15564
rect 10100 15512 10106 15564
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 10253 15552 10281 15592
rect 10183 15524 10281 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 10318 15512 10324 15564
rect 10376 15512 10382 15564
rect 10505 15555 10563 15561
rect 10505 15521 10517 15555
rect 10551 15552 10563 15555
rect 10612 15552 10640 15592
rect 11054 15580 11060 15632
rect 11112 15580 11118 15632
rect 10551 15524 10640 15552
rect 10551 15521 10563 15524
rect 10505 15515 10563 15521
rect 10686 15512 10692 15564
rect 10744 15512 10750 15564
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15552 10839 15555
rect 11072 15552 11100 15580
rect 11256 15561 11284 15660
rect 11422 15648 11428 15660
rect 11480 15648 11486 15700
rect 11701 15691 11759 15697
rect 11701 15657 11713 15691
rect 11747 15688 11759 15691
rect 12618 15688 12624 15700
rect 11747 15660 12624 15688
rect 11747 15657 11759 15660
rect 11701 15651 11759 15657
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 13541 15691 13599 15697
rect 13541 15657 13553 15691
rect 13587 15688 13599 15691
rect 13725 15691 13783 15697
rect 13725 15688 13737 15691
rect 13587 15660 13737 15688
rect 13587 15657 13599 15660
rect 13541 15651 13599 15657
rect 13725 15657 13737 15660
rect 13771 15657 13783 15691
rect 13725 15651 13783 15657
rect 14093 15691 14151 15697
rect 14093 15657 14105 15691
rect 14139 15688 14151 15691
rect 14826 15688 14832 15700
rect 14139 15660 14832 15688
rect 14139 15657 14151 15660
rect 14093 15651 14151 15657
rect 14826 15648 14832 15660
rect 14884 15648 14890 15700
rect 15105 15691 15163 15697
rect 15105 15657 15117 15691
rect 15151 15688 15163 15691
rect 15289 15691 15347 15697
rect 15289 15688 15301 15691
rect 15151 15660 15301 15688
rect 15151 15657 15163 15660
rect 15105 15651 15163 15657
rect 15289 15657 15301 15660
rect 15335 15657 15347 15691
rect 15289 15651 15347 15657
rect 15470 15648 15476 15700
rect 15528 15648 15534 15700
rect 15654 15648 15660 15700
rect 15712 15688 15718 15700
rect 16761 15691 16819 15697
rect 16761 15688 16773 15691
rect 15712 15660 16773 15688
rect 15712 15648 15718 15660
rect 16761 15657 16773 15660
rect 16807 15657 16819 15691
rect 18322 15688 18328 15700
rect 16761 15651 16819 15657
rect 18248 15660 18328 15688
rect 11882 15620 11888 15632
rect 11348 15592 11888 15620
rect 11348 15561 11376 15592
rect 11882 15580 11888 15592
rect 11940 15580 11946 15632
rect 12805 15623 12863 15629
rect 12805 15620 12817 15623
rect 12084 15592 12817 15620
rect 10827 15524 11100 15552
rect 11241 15555 11299 15561
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 11241 15521 11253 15555
rect 11287 15521 11299 15555
rect 11241 15515 11299 15521
rect 11333 15555 11391 15561
rect 11333 15521 11345 15555
rect 11379 15521 11391 15555
rect 11333 15515 11391 15521
rect 11422 15512 11428 15564
rect 11480 15512 11486 15564
rect 11698 15552 11704 15564
rect 11532 15524 11704 15552
rect 9692 15484 9720 15512
rect 10413 15487 10471 15493
rect 10413 15484 10425 15487
rect 8536 15456 9720 15484
rect 9784 15456 10425 15484
rect 8536 15444 8542 15456
rect 8570 15376 8576 15428
rect 8628 15416 8634 15428
rect 9309 15419 9367 15425
rect 9309 15416 9321 15419
rect 8628 15388 9321 15416
rect 8628 15376 8634 15388
rect 9309 15385 9321 15388
rect 9355 15385 9367 15419
rect 9309 15379 9367 15385
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 9784 15416 9812 15456
rect 10413 15453 10425 15456
rect 10459 15453 10471 15487
rect 10704 15484 10732 15512
rect 11054 15484 11060 15496
rect 10704 15456 11060 15484
rect 10413 15447 10471 15453
rect 11054 15444 11060 15456
rect 11112 15444 11118 15496
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15484 11207 15487
rect 11532 15484 11560 15524
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 11790 15512 11796 15564
rect 11848 15512 11854 15564
rect 12084 15561 12112 15592
rect 12805 15589 12817 15592
rect 12851 15589 12863 15623
rect 14734 15620 14740 15632
rect 12805 15583 12863 15589
rect 14476 15592 14740 15620
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15521 12127 15555
rect 12069 15515 12127 15521
rect 11195 15456 11560 15484
rect 11195 15453 11207 15456
rect 11149 15447 11207 15453
rect 11974 15444 11980 15496
rect 12032 15444 12038 15496
rect 10689 15419 10747 15425
rect 10689 15416 10701 15419
rect 9640 15388 9812 15416
rect 9876 15388 10701 15416
rect 9640 15376 9646 15388
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 9033 15351 9091 15357
rect 9033 15348 9045 15351
rect 8352 15320 9045 15348
rect 8352 15308 8358 15320
rect 9033 15317 9045 15320
rect 9079 15317 9091 15351
rect 9033 15311 9091 15317
rect 9122 15308 9128 15360
rect 9180 15348 9186 15360
rect 9876 15348 9904 15388
rect 10689 15385 10701 15388
rect 10735 15385 10747 15419
rect 10689 15379 10747 15385
rect 10778 15376 10784 15428
rect 10836 15416 10842 15428
rect 12084 15416 12112 15515
rect 12158 15512 12164 15564
rect 12216 15512 12222 15564
rect 12434 15512 12440 15564
rect 12492 15512 12498 15564
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 12894 15552 12900 15564
rect 12759 15524 12900 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 12986 15512 12992 15564
rect 13044 15552 13050 15564
rect 13173 15555 13231 15561
rect 13173 15552 13185 15555
rect 13044 15524 13185 15552
rect 13044 15512 13050 15524
rect 13173 15521 13185 15524
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 13262 15512 13268 15564
rect 13320 15552 13326 15564
rect 13449 15555 13507 15561
rect 13449 15552 13461 15555
rect 13320 15524 13461 15552
rect 13320 15512 13326 15524
rect 13449 15521 13461 15524
rect 13495 15521 13507 15555
rect 13449 15515 13507 15521
rect 13722 15512 13728 15564
rect 13780 15512 13786 15564
rect 13906 15512 13912 15564
rect 13964 15512 13970 15564
rect 14476 15561 14504 15592
rect 14734 15580 14740 15592
rect 14792 15620 14798 15632
rect 15488 15620 15516 15648
rect 14792 15592 15056 15620
rect 14792 15580 14798 15592
rect 15028 15561 15056 15592
rect 15304 15592 15516 15620
rect 15856 15592 16436 15620
rect 15304 15561 15332 15592
rect 14185 15555 14243 15561
rect 14185 15521 14197 15555
rect 14231 15552 14243 15555
rect 14369 15555 14427 15561
rect 14369 15552 14381 15555
rect 14231 15524 14381 15552
rect 14231 15521 14243 15524
rect 14185 15515 14243 15521
rect 14369 15521 14381 15524
rect 14415 15521 14427 15555
rect 14369 15515 14427 15521
rect 14461 15555 14519 15561
rect 14461 15521 14473 15555
rect 14507 15521 14519 15555
rect 14461 15515 14519 15521
rect 14553 15555 14611 15561
rect 14553 15521 14565 15555
rect 14599 15521 14611 15555
rect 14553 15515 14611 15521
rect 15013 15555 15071 15561
rect 15013 15521 15025 15555
rect 15059 15521 15071 15555
rect 15013 15515 15071 15521
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15521 15347 15555
rect 15289 15515 15347 15521
rect 15473 15555 15531 15561
rect 15473 15521 15485 15555
rect 15519 15521 15531 15555
rect 15473 15515 15531 15521
rect 15565 15555 15623 15561
rect 15565 15521 15577 15555
rect 15611 15552 15623 15555
rect 15611 15524 15792 15552
rect 15611 15521 15623 15524
rect 15565 15515 15623 15521
rect 14568 15484 14596 15515
rect 14292 15456 14596 15484
rect 14292 15428 14320 15456
rect 10836 15388 12112 15416
rect 10836 15376 10842 15388
rect 14274 15376 14280 15428
rect 14332 15376 14338 15428
rect 9180 15320 9904 15348
rect 9180 15308 9186 15320
rect 11422 15308 11428 15360
rect 11480 15348 11486 15360
rect 12253 15351 12311 15357
rect 12253 15348 12265 15351
rect 11480 15320 12265 15348
rect 11480 15308 11486 15320
rect 12253 15317 12265 15320
rect 12299 15317 12311 15351
rect 12253 15311 12311 15317
rect 12526 15308 12532 15360
rect 12584 15308 12590 15360
rect 13262 15308 13268 15360
rect 13320 15308 13326 15360
rect 14182 15308 14188 15360
rect 14240 15348 14246 15360
rect 14645 15351 14703 15357
rect 14645 15348 14657 15351
rect 14240 15320 14657 15348
rect 14240 15308 14246 15320
rect 14645 15317 14657 15320
rect 14691 15317 14703 15351
rect 15028 15348 15056 15515
rect 15488 15484 15516 15515
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 15488 15456 15669 15484
rect 15657 15453 15669 15456
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 15470 15376 15476 15428
rect 15528 15416 15534 15428
rect 15764 15416 15792 15524
rect 15528 15388 15792 15416
rect 15528 15376 15534 15388
rect 15856 15348 15884 15592
rect 16408 15561 16436 15592
rect 16301 15555 16359 15561
rect 16301 15521 16313 15555
rect 16347 15521 16359 15555
rect 16301 15515 16359 15521
rect 16393 15555 16451 15561
rect 16393 15521 16405 15555
rect 16439 15521 16451 15555
rect 16393 15515 16451 15521
rect 16316 15484 16344 15515
rect 16666 15512 16672 15564
rect 16724 15550 16730 15564
rect 16724 15522 16767 15550
rect 16724 15512 16730 15522
rect 16850 15512 16856 15564
rect 16908 15552 16914 15564
rect 16945 15555 17003 15561
rect 16945 15552 16957 15555
rect 16908 15524 16957 15552
rect 16908 15512 16914 15524
rect 16945 15521 16957 15524
rect 16991 15521 17003 15555
rect 16945 15515 17003 15521
rect 17405 15555 17463 15561
rect 17405 15521 17417 15555
rect 17451 15552 17463 15555
rect 17589 15555 17647 15561
rect 17589 15552 17601 15555
rect 17451 15524 17601 15552
rect 17451 15521 17463 15524
rect 17405 15515 17463 15521
rect 17589 15521 17601 15524
rect 17635 15521 17647 15555
rect 17589 15515 17647 15521
rect 17681 15555 17739 15561
rect 17681 15521 17693 15555
rect 17727 15552 17739 15555
rect 17773 15555 17831 15561
rect 17773 15552 17785 15555
rect 17727 15524 17785 15552
rect 17727 15521 17739 15524
rect 17681 15515 17739 15521
rect 17773 15521 17785 15524
rect 17819 15552 17831 15555
rect 17954 15552 17960 15564
rect 17819 15524 17960 15552
rect 17819 15521 17831 15524
rect 17773 15515 17831 15521
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 18248 15561 18276 15660
rect 18322 15648 18328 15660
rect 18380 15688 18386 15700
rect 18966 15688 18972 15700
rect 18380 15660 18972 15688
rect 18380 15648 18386 15660
rect 18966 15648 18972 15660
rect 19024 15648 19030 15700
rect 19058 15648 19064 15700
rect 19116 15688 19122 15700
rect 19153 15691 19211 15697
rect 19153 15688 19165 15691
rect 19116 15660 19165 15688
rect 19116 15648 19122 15660
rect 19153 15657 19165 15660
rect 19199 15657 19211 15691
rect 19153 15651 19211 15657
rect 19518 15648 19524 15700
rect 19576 15688 19582 15700
rect 20349 15691 20407 15697
rect 20349 15688 20361 15691
rect 19576 15660 20361 15688
rect 19576 15648 19582 15660
rect 20349 15657 20361 15660
rect 20395 15657 20407 15691
rect 20530 15688 20536 15700
rect 20349 15651 20407 15657
rect 20456 15660 20536 15688
rect 18414 15580 18420 15632
rect 18472 15620 18478 15632
rect 18472 15592 19748 15620
rect 18472 15580 18478 15592
rect 18233 15555 18291 15561
rect 18233 15521 18245 15555
rect 18279 15521 18291 15555
rect 18233 15515 18291 15521
rect 18322 15512 18328 15564
rect 18380 15512 18386 15564
rect 18785 15555 18843 15561
rect 18785 15521 18797 15555
rect 18831 15552 18843 15555
rect 18969 15555 19027 15561
rect 18969 15552 18981 15555
rect 18831 15524 18981 15552
rect 18831 15521 18843 15524
rect 18785 15515 18843 15521
rect 18969 15521 18981 15524
rect 19015 15521 19027 15555
rect 18969 15515 19027 15521
rect 19058 15512 19064 15564
rect 19116 15512 19122 15564
rect 19153 15555 19211 15561
rect 19153 15521 19165 15555
rect 19199 15521 19211 15555
rect 19153 15515 19211 15521
rect 19337 15555 19395 15561
rect 19337 15521 19349 15555
rect 19383 15552 19395 15555
rect 19426 15552 19432 15564
rect 19383 15524 19432 15552
rect 19383 15521 19395 15524
rect 19337 15515 19395 15521
rect 17037 15487 17095 15493
rect 17037 15484 17049 15487
rect 16316 15456 17049 15484
rect 17037 15453 17049 15456
rect 17083 15453 17095 15487
rect 17037 15447 17095 15453
rect 17865 15487 17923 15493
rect 17865 15453 17877 15487
rect 17911 15484 17923 15487
rect 18874 15484 18880 15496
rect 17911 15456 18880 15484
rect 17911 15453 17923 15456
rect 17865 15447 17923 15453
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 19168 15484 19196 15515
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 19720 15561 19748 15592
rect 19794 15580 19800 15632
rect 19852 15580 19858 15632
rect 20070 15620 20076 15632
rect 19904 15592 20076 15620
rect 19613 15555 19671 15561
rect 19613 15521 19625 15555
rect 19659 15521 19671 15555
rect 19613 15515 19671 15521
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15521 19763 15555
rect 19705 15515 19763 15521
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 19168 15456 19533 15484
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 16209 15419 16267 15425
rect 16209 15385 16221 15419
rect 16255 15416 16267 15419
rect 17494 15416 17500 15428
rect 16255 15388 17500 15416
rect 16255 15385 16267 15388
rect 16209 15379 16267 15385
rect 17494 15376 17500 15388
rect 17552 15376 17558 15428
rect 18417 15419 18475 15425
rect 18417 15385 18429 15419
rect 18463 15416 18475 15419
rect 18463 15388 19288 15416
rect 18463 15385 18475 15388
rect 18417 15379 18475 15385
rect 15028 15320 15884 15348
rect 16485 15351 16543 15357
rect 14645 15311 14703 15317
rect 16485 15317 16497 15351
rect 16531 15348 16543 15351
rect 16666 15348 16672 15360
rect 16531 15320 16672 15348
rect 16531 15317 16543 15320
rect 16485 15311 16543 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 17310 15308 17316 15360
rect 17368 15308 17374 15360
rect 18138 15308 18144 15360
rect 18196 15308 18202 15360
rect 18693 15351 18751 15357
rect 18693 15317 18705 15351
rect 18739 15348 18751 15351
rect 19058 15348 19064 15360
rect 18739 15320 19064 15348
rect 18739 15317 18751 15320
rect 18693 15311 18751 15317
rect 19058 15308 19064 15320
rect 19116 15308 19122 15360
rect 19260 15348 19288 15388
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 19628 15416 19656 15515
rect 19904 15484 19932 15592
rect 20070 15580 20076 15592
rect 20128 15580 20134 15632
rect 20456 15561 20484 15660
rect 20530 15648 20536 15660
rect 20588 15688 20594 15700
rect 22094 15688 22100 15700
rect 20588 15660 22100 15688
rect 20588 15648 20594 15660
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 22278 15648 22284 15700
rect 22336 15688 22342 15700
rect 22336 15660 22692 15688
rect 22336 15648 22342 15660
rect 22462 15620 22468 15632
rect 20732 15592 22468 15620
rect 20732 15564 20760 15592
rect 19981 15555 20039 15561
rect 19981 15521 19993 15555
rect 20027 15552 20039 15555
rect 20441 15555 20499 15561
rect 20441 15552 20453 15555
rect 20027 15524 20453 15552
rect 20027 15521 20039 15524
rect 19981 15515 20039 15521
rect 20441 15521 20453 15524
rect 20487 15521 20499 15555
rect 20441 15515 20499 15521
rect 20533 15555 20591 15561
rect 20533 15521 20545 15555
rect 20579 15521 20591 15555
rect 20533 15515 20591 15521
rect 20548 15484 20576 15515
rect 20714 15512 20720 15564
rect 20772 15512 20778 15564
rect 20809 15555 20867 15561
rect 20809 15521 20821 15555
rect 20855 15552 20867 15555
rect 21266 15552 21272 15564
rect 20855 15524 21272 15552
rect 20855 15521 20867 15524
rect 20809 15515 20867 15521
rect 21266 15512 21272 15524
rect 21324 15512 21330 15564
rect 21560 15561 21588 15592
rect 22462 15580 22468 15592
rect 22520 15580 22526 15632
rect 21545 15555 21603 15561
rect 21545 15521 21557 15555
rect 21591 15521 21603 15555
rect 21545 15515 21603 15521
rect 21910 15512 21916 15564
rect 21968 15512 21974 15564
rect 22002 15512 22008 15564
rect 22060 15512 22066 15564
rect 22278 15512 22284 15564
rect 22336 15512 22342 15564
rect 22370 15512 22376 15564
rect 22428 15512 22434 15564
rect 22664 15561 22692 15660
rect 22922 15648 22928 15700
rect 22980 15688 22986 15700
rect 23017 15691 23075 15697
rect 23017 15688 23029 15691
rect 22980 15660 23029 15688
rect 22980 15648 22986 15660
rect 23017 15657 23029 15660
rect 23063 15657 23075 15691
rect 23017 15651 23075 15657
rect 23290 15648 23296 15700
rect 23348 15688 23354 15700
rect 24397 15691 24455 15697
rect 24397 15688 24409 15691
rect 23348 15660 24409 15688
rect 23348 15648 23354 15660
rect 24397 15657 24409 15660
rect 24443 15657 24455 15691
rect 24397 15651 24455 15657
rect 24946 15648 24952 15700
rect 25004 15648 25010 15700
rect 24026 15620 24032 15632
rect 23124 15592 24032 15620
rect 23124 15561 23152 15592
rect 24026 15580 24032 15592
rect 24084 15580 24090 15632
rect 24118 15580 24124 15632
rect 24176 15580 24182 15632
rect 25682 15620 25688 15632
rect 24504 15592 25688 15620
rect 22557 15555 22615 15561
rect 22557 15521 22569 15555
rect 22603 15521 22615 15555
rect 22557 15515 22615 15521
rect 22649 15555 22707 15561
rect 22649 15521 22661 15555
rect 22695 15521 22707 15555
rect 22649 15515 22707 15521
rect 23109 15555 23167 15561
rect 23109 15521 23121 15555
rect 23155 15521 23167 15555
rect 23109 15515 23167 15521
rect 23385 15555 23443 15561
rect 23385 15521 23397 15555
rect 23431 15552 23443 15555
rect 23569 15555 23627 15561
rect 23569 15552 23581 15555
rect 23431 15524 23581 15552
rect 23431 15521 23443 15524
rect 23385 15515 23443 15521
rect 23569 15521 23581 15524
rect 23615 15521 23627 15555
rect 23569 15515 23627 15521
rect 23661 15555 23719 15561
rect 23661 15521 23673 15555
rect 23707 15552 23719 15555
rect 23937 15555 23995 15561
rect 23707 15524 23888 15552
rect 23707 15521 23719 15524
rect 23661 15515 23719 15521
rect 19904 15456 20576 15484
rect 22572 15484 22600 15515
rect 23860 15496 23888 15524
rect 23937 15521 23949 15555
rect 23983 15521 23995 15555
rect 23937 15515 23995 15521
rect 23290 15484 23296 15496
rect 22572 15456 23296 15484
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 23842 15444 23848 15496
rect 23900 15444 23906 15496
rect 23952 15484 23980 15515
rect 24210 15512 24216 15564
rect 24268 15552 24274 15564
rect 24305 15555 24363 15561
rect 24305 15552 24317 15555
rect 24268 15524 24317 15552
rect 24268 15512 24274 15524
rect 24305 15521 24317 15524
rect 24351 15521 24363 15555
rect 24305 15515 24363 15521
rect 24504 15484 24532 15592
rect 25682 15580 25688 15592
rect 25740 15580 25746 15632
rect 24578 15512 24584 15564
rect 24636 15512 24642 15564
rect 24854 15512 24860 15564
rect 24912 15512 24918 15564
rect 23952 15456 24532 15484
rect 24673 15487 24731 15493
rect 24673 15453 24685 15487
rect 24719 15484 24731 15487
rect 26326 15484 26332 15496
rect 24719 15456 26332 15484
rect 24719 15453 24731 15456
rect 24673 15447 24731 15453
rect 26326 15444 26332 15456
rect 26384 15444 26390 15496
rect 19392 15388 19656 15416
rect 20073 15419 20131 15425
rect 19392 15376 19398 15388
rect 19536 15360 19564 15388
rect 20073 15385 20085 15419
rect 20119 15416 20131 15419
rect 20990 15416 20996 15428
rect 20119 15388 20996 15416
rect 20119 15385 20131 15388
rect 20073 15379 20131 15385
rect 20990 15376 20996 15388
rect 21048 15376 21054 15428
rect 22186 15376 22192 15428
rect 22244 15376 22250 15428
rect 22465 15419 22523 15425
rect 22465 15385 22477 15419
rect 22511 15416 22523 15419
rect 25314 15416 25320 15428
rect 22511 15388 25320 15416
rect 22511 15385 22523 15388
rect 22465 15379 22523 15385
rect 25314 15376 25320 15388
rect 25372 15376 25378 15428
rect 19426 15348 19432 15360
rect 19260 15320 19432 15348
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 19518 15308 19524 15360
rect 19576 15308 19582 15360
rect 20346 15308 20352 15360
rect 20404 15348 20410 15360
rect 20625 15351 20683 15357
rect 20625 15348 20637 15351
rect 20404 15320 20637 15348
rect 20404 15308 20410 15320
rect 20625 15317 20637 15320
rect 20671 15317 20683 15351
rect 20625 15311 20683 15317
rect 20901 15351 20959 15357
rect 20901 15317 20913 15351
rect 20947 15348 20959 15351
rect 21174 15348 21180 15360
rect 20947 15320 21180 15348
rect 20947 15317 20959 15320
rect 20901 15311 20959 15317
rect 21174 15308 21180 15320
rect 21232 15308 21238 15360
rect 21358 15308 21364 15360
rect 21416 15308 21422 15360
rect 21634 15308 21640 15360
rect 21692 15308 21698 15360
rect 22094 15308 22100 15360
rect 22152 15348 22158 15360
rect 22741 15351 22799 15357
rect 22741 15348 22753 15351
rect 22152 15320 22753 15348
rect 22152 15308 22158 15320
rect 22741 15317 22753 15320
rect 22787 15317 22799 15351
rect 22741 15311 22799 15317
rect 23293 15351 23351 15357
rect 23293 15317 23305 15351
rect 23339 15348 23351 15351
rect 23474 15348 23480 15360
rect 23339 15320 23480 15348
rect 23339 15317 23351 15320
rect 23293 15311 23351 15317
rect 23474 15308 23480 15320
rect 23532 15308 23538 15360
rect 23845 15351 23903 15357
rect 23845 15317 23857 15351
rect 23891 15348 23903 15351
rect 24210 15348 24216 15360
rect 23891 15320 24216 15348
rect 23891 15317 23903 15320
rect 23845 15311 23903 15317
rect 24210 15308 24216 15320
rect 24268 15308 24274 15360
rect 552 15258 31372 15280
rect 552 15206 4250 15258
rect 4302 15206 4314 15258
rect 4366 15206 4378 15258
rect 4430 15206 4442 15258
rect 4494 15206 4506 15258
rect 4558 15206 11955 15258
rect 12007 15206 12019 15258
rect 12071 15206 12083 15258
rect 12135 15206 12147 15258
rect 12199 15206 12211 15258
rect 12263 15206 19660 15258
rect 19712 15206 19724 15258
rect 19776 15206 19788 15258
rect 19840 15206 19852 15258
rect 19904 15206 19916 15258
rect 19968 15206 27365 15258
rect 27417 15206 27429 15258
rect 27481 15206 27493 15258
rect 27545 15206 27557 15258
rect 27609 15206 27621 15258
rect 27673 15206 31372 15258
rect 552 15184 31372 15206
rect 8662 15104 8668 15156
rect 8720 15104 8726 15156
rect 9033 15147 9091 15153
rect 9033 15113 9045 15147
rect 9079 15144 9091 15147
rect 9766 15144 9772 15156
rect 9079 15116 9772 15144
rect 9079 15113 9091 15116
rect 9033 15107 9091 15113
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 10137 15147 10195 15153
rect 10137 15113 10149 15147
rect 10183 15144 10195 15147
rect 10226 15144 10232 15156
rect 10183 15116 10232 15144
rect 10183 15113 10195 15116
rect 10137 15107 10195 15113
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 10502 15104 10508 15156
rect 10560 15104 10566 15156
rect 10689 15147 10747 15153
rect 10689 15113 10701 15147
rect 10735 15144 10747 15147
rect 12710 15144 12716 15156
rect 10735 15116 12716 15144
rect 10735 15113 10747 15116
rect 10689 15107 10747 15113
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 13630 15104 13636 15156
rect 13688 15104 13694 15156
rect 13722 15104 13728 15156
rect 13780 15104 13786 15156
rect 13906 15104 13912 15156
rect 13964 15104 13970 15156
rect 16577 15147 16635 15153
rect 16577 15113 16589 15147
rect 16623 15144 16635 15147
rect 17402 15144 17408 15156
rect 16623 15116 17408 15144
rect 16623 15113 16635 15116
rect 16577 15107 16635 15113
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 18322 15104 18328 15156
rect 18380 15144 18386 15156
rect 18417 15147 18475 15153
rect 18417 15144 18429 15147
rect 18380 15116 18429 15144
rect 18380 15104 18386 15116
rect 18417 15113 18429 15116
rect 18463 15113 18475 15147
rect 18417 15107 18475 15113
rect 19334 15104 19340 15156
rect 19392 15144 19398 15156
rect 20073 15147 20131 15153
rect 19392 15116 19656 15144
rect 19392 15104 19398 15116
rect 8680 15008 8708 15104
rect 10520 15076 10548 15104
rect 9140 15048 10548 15076
rect 12621 15079 12679 15085
rect 7944 14980 8432 15008
rect 8680 14980 8892 15008
rect 7944 14949 7972 14980
rect 8404 14949 8432 14980
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14909 7987 14943
rect 7929 14903 7987 14909
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14909 8079 14943
rect 8021 14903 8079 14909
rect 8389 14943 8447 14949
rect 8389 14909 8401 14943
rect 8435 14940 8447 14943
rect 8478 14940 8484 14952
rect 8435 14912 8484 14940
rect 8435 14909 8447 14912
rect 8389 14903 8447 14909
rect 7837 14875 7895 14881
rect 7837 14841 7849 14875
rect 7883 14872 7895 14875
rect 8036 14872 8064 14903
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 8665 14943 8723 14949
rect 8665 14909 8677 14943
rect 8711 14940 8723 14943
rect 8754 14940 8760 14952
rect 8711 14912 8760 14940
rect 8711 14909 8723 14912
rect 8665 14903 8723 14909
rect 8754 14900 8760 14912
rect 8812 14900 8818 14952
rect 8864 14949 8892 14980
rect 9140 14949 9168 15048
rect 12621 15045 12633 15079
rect 12667 15076 12679 15079
rect 13740 15076 13768 15104
rect 12667 15048 13768 15076
rect 12667 15045 12679 15048
rect 12621 15039 12679 15045
rect 9582 14968 9588 15020
rect 9640 14968 9646 15020
rect 10873 15011 10931 15017
rect 10873 15008 10885 15011
rect 9784 14980 10088 15008
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14909 8907 14943
rect 8849 14903 8907 14909
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14909 9183 14943
rect 9125 14903 9183 14909
rect 9306 14900 9312 14952
rect 9364 14940 9370 14952
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 9364 14912 9413 14940
rect 9364 14900 9370 14912
rect 9401 14909 9413 14912
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 9674 14900 9680 14952
rect 9732 14900 9738 14952
rect 7883 14844 8064 14872
rect 8113 14875 8171 14881
rect 7883 14841 7895 14844
rect 7837 14835 7895 14841
rect 8113 14841 8125 14875
rect 8159 14872 8171 14875
rect 8159 14844 9444 14872
rect 8159 14841 8171 14844
rect 8113 14835 8171 14841
rect 7190 14764 7196 14816
rect 7248 14804 7254 14816
rect 8294 14804 8300 14816
rect 7248 14776 8300 14804
rect 7248 14764 7254 14776
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 8481 14807 8539 14813
rect 8481 14773 8493 14807
rect 8527 14804 8539 14807
rect 8665 14807 8723 14813
rect 8665 14804 8677 14807
rect 8527 14776 8677 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 8665 14773 8677 14776
rect 8711 14773 8723 14807
rect 8665 14767 8723 14773
rect 9306 14764 9312 14816
rect 9364 14764 9370 14816
rect 9416 14804 9444 14844
rect 9490 14832 9496 14884
rect 9548 14872 9554 14884
rect 9784 14872 9812 14980
rect 9950 14900 9956 14952
rect 10008 14900 10014 14952
rect 10060 14949 10088 14980
rect 10152 14980 10885 15008
rect 10152 14952 10180 14980
rect 10873 14977 10885 14980
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 12897 15011 12955 15017
rect 12897 14977 12909 15011
rect 12943 15008 12955 15011
rect 13924 15008 13952 15104
rect 18141 15079 18199 15085
rect 18141 15045 18153 15079
rect 18187 15076 18199 15079
rect 18598 15076 18604 15088
rect 18187 15048 18604 15076
rect 18187 15045 18199 15048
rect 18141 15039 18199 15045
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 19628 15076 19656 15116
rect 20073 15113 20085 15147
rect 20119 15144 20131 15147
rect 20806 15144 20812 15156
rect 20119 15116 20812 15144
rect 20119 15113 20131 15116
rect 20073 15107 20131 15113
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 22186 15144 22192 15156
rect 21836 15116 22192 15144
rect 20346 15076 20352 15088
rect 19628 15048 20352 15076
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 21836 15017 21864 15116
rect 22186 15104 22192 15116
rect 22244 15104 22250 15156
rect 22554 15104 22560 15156
rect 22612 15144 22618 15156
rect 23477 15147 23535 15153
rect 23477 15144 23489 15147
rect 22612 15116 23489 15144
rect 22612 15104 22618 15116
rect 23477 15113 23489 15116
rect 23523 15113 23535 15147
rect 23477 15107 23535 15113
rect 23934 15104 23940 15156
rect 23992 15104 23998 15156
rect 24210 15104 24216 15156
rect 24268 15144 24274 15156
rect 28258 15144 28264 15156
rect 24268 15116 28264 15144
rect 24268 15104 24274 15116
rect 28258 15104 28264 15116
rect 28316 15104 28322 15156
rect 23198 15036 23204 15088
rect 23256 15036 23262 15088
rect 24765 15079 24823 15085
rect 24765 15076 24777 15079
rect 23308 15048 24777 15076
rect 18693 15011 18751 15017
rect 18693 15008 18705 15011
rect 12943 14980 13952 15008
rect 17880 14980 18705 15008
rect 12943 14977 12955 14980
rect 12897 14971 12955 14977
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14909 10103 14943
rect 10045 14903 10103 14909
rect 10134 14900 10140 14952
rect 10192 14900 10198 14952
rect 10318 14900 10324 14952
rect 10376 14900 10382 14952
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14909 10563 14943
rect 10505 14903 10563 14909
rect 9548 14844 9812 14872
rect 9861 14875 9919 14881
rect 9548 14832 9554 14844
rect 9861 14841 9873 14875
rect 9907 14841 9919 14875
rect 10336 14872 10364 14900
rect 9861 14835 9919 14841
rect 10152 14844 10364 14872
rect 10520 14872 10548 14903
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 10781 14943 10839 14949
rect 10781 14940 10793 14943
rect 10744 14912 10793 14940
rect 10744 14900 10750 14912
rect 10781 14909 10793 14912
rect 10827 14909 10839 14943
rect 11514 14940 11520 14952
rect 10781 14903 10839 14909
rect 10888 14912 11520 14940
rect 10888 14872 10916 14912
rect 11514 14900 11520 14912
rect 11572 14900 11578 14952
rect 11606 14900 11612 14952
rect 11664 14900 11670 14952
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 10520 14844 10916 14872
rect 9766 14804 9772 14816
rect 9416 14776 9772 14804
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 9876 14804 9904 14835
rect 10152 14804 10180 14844
rect 10962 14832 10968 14884
rect 11020 14872 11026 14884
rect 11118 14875 11176 14881
rect 11118 14872 11130 14875
rect 11020 14844 11130 14872
rect 11020 14832 11026 14844
rect 11118 14841 11130 14844
rect 11164 14841 11176 14875
rect 11118 14835 11176 14841
rect 9876 14776 10180 14804
rect 10410 14764 10416 14816
rect 10468 14764 10474 14816
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 11330 14804 11336 14816
rect 10652 14776 11336 14804
rect 10652 14764 10658 14776
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 11624 14804 11652 14900
rect 11790 14832 11796 14884
rect 11848 14872 11854 14884
rect 12544 14872 12572 14903
rect 11848 14844 12572 14872
rect 13004 14872 13032 14903
rect 13078 14900 13084 14952
rect 13136 14900 13142 14952
rect 13814 14900 13820 14952
rect 13872 14900 13878 14952
rect 15013 14943 15071 14949
rect 15013 14940 15025 14943
rect 14016 14912 15025 14940
rect 13832 14872 13860 14900
rect 14016 14884 14044 14912
rect 15013 14909 15025 14912
rect 15059 14940 15071 14943
rect 15197 14943 15255 14949
rect 15197 14940 15209 14943
rect 15059 14912 15209 14940
rect 15059 14909 15071 14912
rect 15013 14903 15071 14909
rect 15197 14909 15209 14912
rect 15243 14909 15255 14943
rect 15197 14903 15255 14909
rect 16761 14943 16819 14949
rect 16761 14909 16773 14943
rect 16807 14940 16819 14943
rect 17770 14940 17776 14952
rect 16807 14912 17776 14940
rect 16807 14909 16819 14912
rect 16761 14903 16819 14909
rect 17770 14900 17776 14912
rect 17828 14940 17834 14952
rect 17880 14940 17908 14980
rect 18693 14977 18705 14980
rect 18739 14977 18751 15011
rect 18693 14971 18751 14977
rect 21729 15011 21787 15017
rect 21729 14977 21741 15011
rect 21775 15008 21787 15011
rect 21821 15011 21879 15017
rect 21821 15008 21833 15011
rect 21775 14980 21833 15008
rect 21775 14977 21787 14980
rect 21729 14971 21787 14977
rect 21821 14977 21833 14980
rect 21867 14977 21879 15011
rect 21821 14971 21879 14977
rect 17828 14912 17908 14940
rect 17828 14900 17834 14912
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 18325 14943 18383 14949
rect 18325 14940 18337 14943
rect 18196 14912 18337 14940
rect 18196 14900 18202 14912
rect 18325 14909 18337 14912
rect 18371 14909 18383 14943
rect 18325 14903 18383 14909
rect 18960 14943 19018 14949
rect 18960 14909 18972 14943
rect 19006 14940 19018 14943
rect 20254 14940 20260 14952
rect 19006 14912 20260 14940
rect 19006 14909 19018 14912
rect 18960 14903 19018 14909
rect 20254 14900 20260 14912
rect 20312 14900 20318 14952
rect 21473 14943 21531 14949
rect 21473 14909 21485 14943
rect 21519 14940 21531 14943
rect 23308 14940 23336 15048
rect 24765 15045 24777 15048
rect 24811 15045 24823 15079
rect 24765 15039 24823 15045
rect 25038 15036 25044 15088
rect 25096 15036 25102 15088
rect 25130 15036 25136 15088
rect 25188 15076 25194 15088
rect 25317 15079 25375 15085
rect 25317 15076 25329 15079
rect 25188 15048 25329 15076
rect 25188 15036 25194 15048
rect 25317 15045 25329 15048
rect 25363 15045 25375 15079
rect 25317 15039 25375 15045
rect 23474 14968 23480 15020
rect 23532 15008 23538 15020
rect 23532 14980 23612 15008
rect 23532 14968 23538 14980
rect 21519 14912 23336 14940
rect 21519 14909 21531 14912
rect 21473 14903 21531 14909
rect 23382 14900 23388 14952
rect 23440 14900 23446 14952
rect 23584 14949 23612 14980
rect 24044 14980 28304 15008
rect 23569 14943 23627 14949
rect 23569 14909 23581 14943
rect 23615 14909 23627 14943
rect 23569 14903 23627 14909
rect 23750 14900 23756 14952
rect 23808 14940 23814 14952
rect 23845 14943 23903 14949
rect 23845 14940 23857 14943
rect 23808 14912 23857 14940
rect 23808 14900 23814 14912
rect 23845 14909 23857 14912
rect 23891 14909 23903 14943
rect 23845 14903 23903 14909
rect 13004 14844 13860 14872
rect 11848 14832 11854 14844
rect 12253 14807 12311 14813
rect 12253 14804 12265 14807
rect 11624 14776 12265 14804
rect 12253 14773 12265 14776
rect 12299 14773 12311 14807
rect 12544 14804 12572 14844
rect 13998 14832 14004 14884
rect 14056 14832 14062 14884
rect 14768 14875 14826 14881
rect 14768 14841 14780 14875
rect 14814 14872 14826 14875
rect 15464 14875 15522 14881
rect 14814 14844 15240 14872
rect 14814 14841 14826 14844
rect 14768 14835 14826 14841
rect 15212 14816 15240 14844
rect 15464 14841 15476 14875
rect 15510 14872 15522 14875
rect 15562 14872 15568 14884
rect 15510 14844 15568 14872
rect 15510 14841 15522 14844
rect 15464 14835 15522 14841
rect 15562 14832 15568 14844
rect 15620 14832 15626 14884
rect 17028 14875 17086 14881
rect 17028 14841 17040 14875
rect 17074 14872 17086 14875
rect 17126 14872 17132 14884
rect 17074 14844 17132 14872
rect 17074 14841 17086 14844
rect 17028 14835 17086 14841
rect 17126 14832 17132 14844
rect 17184 14832 17190 14884
rect 21726 14872 21732 14884
rect 20364 14844 21732 14872
rect 12986 14804 12992 14816
rect 12544 14776 12992 14804
rect 12253 14767 12311 14773
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 13170 14764 13176 14816
rect 13228 14764 13234 14816
rect 13538 14764 13544 14816
rect 13596 14804 13602 14816
rect 14274 14804 14280 14816
rect 13596 14776 14280 14804
rect 13596 14764 13602 14776
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 15194 14764 15200 14816
rect 15252 14764 15258 14816
rect 20364 14813 20392 14844
rect 21726 14832 21732 14844
rect 21784 14832 21790 14884
rect 22088 14875 22146 14881
rect 22088 14841 22100 14875
rect 22134 14872 22146 14875
rect 23014 14872 23020 14884
rect 22134 14844 23020 14872
rect 22134 14841 22146 14844
rect 22088 14835 22146 14841
rect 23014 14832 23020 14844
rect 23072 14832 23078 14884
rect 20349 14807 20407 14813
rect 20349 14773 20361 14807
rect 20395 14773 20407 14807
rect 20349 14767 20407 14773
rect 21174 14764 21180 14816
rect 21232 14804 21238 14816
rect 22646 14804 22652 14816
rect 21232 14776 22652 14804
rect 21232 14764 21238 14776
rect 22646 14764 22652 14776
rect 22704 14764 22710 14816
rect 23382 14764 23388 14816
rect 23440 14804 23446 14816
rect 24044 14804 24072 14980
rect 24118 14900 24124 14952
rect 24176 14940 24182 14952
rect 24305 14943 24363 14949
rect 24305 14940 24317 14943
rect 24176 14912 24317 14940
rect 24176 14900 24182 14912
rect 24305 14909 24317 14912
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 24486 14900 24492 14952
rect 24544 14900 24550 14952
rect 24578 14900 24584 14952
rect 24636 14900 24642 14952
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 24762 14900 24768 14952
rect 24820 14940 24826 14952
rect 24949 14943 25007 14949
rect 24949 14940 24961 14943
rect 24820 14912 24961 14940
rect 24820 14900 24826 14912
rect 24949 14909 24961 14912
rect 24995 14909 25007 14943
rect 24949 14903 25007 14909
rect 25222 14900 25228 14952
rect 25280 14900 25286 14952
rect 25501 14943 25559 14949
rect 25501 14909 25513 14943
rect 25547 14909 25559 14943
rect 25501 14903 25559 14909
rect 24504 14872 24532 14900
rect 25516 14872 25544 14903
rect 25866 14872 25872 14884
rect 24504 14844 25872 14872
rect 25866 14832 25872 14844
rect 25924 14832 25930 14884
rect 28276 14816 28304 14980
rect 23440 14776 24072 14804
rect 24213 14807 24271 14813
rect 23440 14764 23446 14776
rect 24213 14773 24225 14807
rect 24259 14804 24271 14807
rect 24394 14804 24400 14816
rect 24259 14776 24400 14804
rect 24259 14773 24271 14776
rect 24213 14767 24271 14773
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 24946 14764 24952 14816
rect 25004 14804 25010 14816
rect 25498 14804 25504 14816
rect 25004 14776 25504 14804
rect 25004 14764 25010 14776
rect 25498 14764 25504 14776
rect 25556 14764 25562 14816
rect 25593 14807 25651 14813
rect 25593 14773 25605 14807
rect 25639 14804 25651 14807
rect 25774 14804 25780 14816
rect 25639 14776 25780 14804
rect 25639 14773 25651 14776
rect 25593 14767 25651 14773
rect 25774 14764 25780 14776
rect 25832 14764 25838 14816
rect 28258 14764 28264 14816
rect 28316 14764 28322 14816
rect 29638 14764 29644 14816
rect 29696 14804 29702 14816
rect 31662 14804 31668 14816
rect 29696 14776 31668 14804
rect 29696 14764 29702 14776
rect 31662 14764 31668 14776
rect 31720 14764 31726 14816
rect 552 14714 31531 14736
rect 552 14662 8102 14714
rect 8154 14662 8166 14714
rect 8218 14662 8230 14714
rect 8282 14662 8294 14714
rect 8346 14662 8358 14714
rect 8410 14662 15807 14714
rect 15859 14662 15871 14714
rect 15923 14662 15935 14714
rect 15987 14662 15999 14714
rect 16051 14662 16063 14714
rect 16115 14662 23512 14714
rect 23564 14662 23576 14714
rect 23628 14662 23640 14714
rect 23692 14662 23704 14714
rect 23756 14662 23768 14714
rect 23820 14662 31217 14714
rect 31269 14662 31281 14714
rect 31333 14662 31345 14714
rect 31397 14662 31409 14714
rect 31461 14662 31473 14714
rect 31525 14662 31531 14714
rect 552 14640 31531 14662
rect 7834 14600 7840 14612
rect 7484 14572 7840 14600
rect 7484 14473 7512 14572
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 7926 14560 7932 14612
rect 7984 14560 7990 14612
rect 8938 14600 8944 14612
rect 8312 14572 8944 14600
rect 7558 14492 7564 14544
rect 7616 14492 7622 14544
rect 7653 14535 7711 14541
rect 7653 14501 7665 14535
rect 7699 14532 7711 14535
rect 8312 14532 8340 14572
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 9033 14603 9091 14609
rect 9033 14569 9045 14603
rect 9079 14600 9091 14603
rect 10226 14600 10232 14612
rect 9079 14572 10232 14600
rect 9079 14569 9091 14572
rect 9033 14563 9091 14569
rect 10226 14560 10232 14572
rect 10284 14560 10290 14612
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 10686 14600 10692 14612
rect 10643 14572 10692 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 13078 14600 13084 14612
rect 11388 14572 13084 14600
rect 11388 14560 11394 14572
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 13357 14603 13415 14609
rect 13357 14569 13369 14603
rect 13403 14600 13415 14603
rect 15470 14600 15476 14612
rect 13403 14572 15476 14600
rect 13403 14569 13415 14572
rect 13357 14563 13415 14569
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 16206 14600 16212 14612
rect 15795 14572 16212 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 16666 14560 16672 14612
rect 16724 14560 16730 14612
rect 16761 14603 16819 14609
rect 16761 14569 16773 14603
rect 16807 14600 16819 14603
rect 16850 14600 16856 14612
rect 16807 14572 16856 14600
rect 16807 14569 16819 14572
rect 16761 14563 16819 14569
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 17310 14560 17316 14612
rect 17368 14560 17374 14612
rect 17681 14603 17739 14609
rect 17681 14569 17693 14603
rect 17727 14600 17739 14603
rect 18969 14603 19027 14609
rect 18969 14600 18981 14603
rect 17727 14572 18981 14600
rect 17727 14569 17739 14572
rect 17681 14563 17739 14569
rect 18969 14569 18981 14572
rect 19015 14569 19027 14603
rect 18969 14563 19027 14569
rect 19058 14560 19064 14612
rect 19116 14560 19122 14612
rect 19150 14560 19156 14612
rect 19208 14600 19214 14612
rect 19208 14572 20024 14600
rect 19208 14560 19214 14572
rect 11054 14532 11060 14544
rect 7699 14504 8340 14532
rect 8588 14504 11060 14532
rect 7699 14501 7711 14504
rect 7653 14495 7711 14501
rect 7469 14467 7527 14473
rect 7469 14433 7481 14467
rect 7515 14433 7527 14467
rect 7576 14464 7604 14492
rect 7745 14467 7803 14473
rect 7745 14464 7757 14467
rect 7576 14436 7757 14464
rect 7469 14427 7527 14433
rect 7745 14433 7757 14436
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 7834 14424 7840 14476
rect 7892 14424 7898 14476
rect 8018 14424 8024 14476
rect 8076 14424 8082 14476
rect 8110 14424 8116 14476
rect 8168 14424 8174 14476
rect 8588 14473 8616 14504
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8266 14436 8585 14464
rect 8266 14396 8294 14436
rect 8573 14433 8585 14436
rect 8619 14433 8631 14467
rect 8573 14427 8631 14433
rect 8662 14424 8668 14476
rect 8720 14424 8726 14476
rect 7116 14368 8294 14396
rect 7116 14272 7144 14368
rect 7377 14331 7435 14337
rect 7377 14297 7389 14331
rect 7423 14328 7435 14331
rect 8294 14328 8300 14340
rect 7423 14300 8300 14328
rect 7423 14297 7435 14300
rect 7377 14291 7435 14297
rect 8294 14288 8300 14300
rect 8352 14288 8358 14340
rect 8680 14328 8708 14424
rect 8864 14408 8892 14504
rect 11054 14492 11060 14504
rect 11112 14532 11118 14544
rect 11241 14535 11299 14541
rect 11241 14532 11253 14535
rect 11112 14504 11253 14532
rect 11112 14492 11118 14504
rect 9122 14424 9128 14476
rect 9180 14424 9186 14476
rect 9473 14467 9531 14473
rect 9473 14433 9485 14467
rect 9519 14464 9531 14467
rect 9766 14464 9772 14476
rect 9519 14436 9772 14464
rect 9519 14433 9531 14436
rect 9473 14427 9531 14433
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 11164 14473 11192 14504
rect 11241 14501 11253 14504
rect 11287 14501 11299 14535
rect 11241 14495 11299 14501
rect 12989 14535 13047 14541
rect 12989 14501 13001 14535
rect 13035 14532 13047 14535
rect 15194 14532 15200 14544
rect 13035 14504 15200 14532
rect 13035 14501 13047 14504
rect 12989 14495 13047 14501
rect 15194 14492 15200 14504
rect 15252 14492 15258 14544
rect 16684 14532 16712 14560
rect 16684 14504 17264 14532
rect 11149 14467 11207 14473
rect 11149 14433 11161 14467
rect 11195 14433 11207 14467
rect 13262 14464 13268 14476
rect 11149 14427 11207 14433
rect 12406 14436 13268 14464
rect 8846 14356 8852 14408
rect 8904 14356 8910 14408
rect 8938 14356 8944 14408
rect 8996 14356 9002 14408
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 8404 14300 8708 14328
rect 8956 14328 8984 14356
rect 9232 14328 9260 14359
rect 10870 14356 10876 14408
rect 10928 14396 10934 14408
rect 12406 14396 12434 14436
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 13446 14424 13452 14476
rect 13504 14424 13510 14476
rect 13725 14467 13783 14473
rect 13725 14433 13737 14467
rect 13771 14433 13783 14467
rect 13725 14427 13783 14433
rect 10928 14368 12434 14396
rect 10928 14356 10934 14368
rect 12802 14356 12808 14408
rect 12860 14396 12866 14408
rect 13633 14399 13691 14405
rect 13633 14396 13645 14399
rect 12860 14368 13645 14396
rect 12860 14356 12866 14368
rect 13633 14365 13645 14368
rect 13679 14365 13691 14399
rect 13740 14396 13768 14427
rect 13814 14424 13820 14476
rect 13872 14424 13878 14476
rect 14182 14464 14188 14476
rect 13924 14436 14188 14464
rect 13924 14396 13952 14436
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 14274 14424 14280 14476
rect 14332 14424 14338 14476
rect 14642 14473 14648 14476
rect 14636 14464 14648 14473
rect 14603 14436 14648 14464
rect 14636 14427 14648 14436
rect 14642 14424 14648 14427
rect 14700 14424 14706 14476
rect 16301 14467 16359 14473
rect 16301 14433 16313 14467
rect 16347 14433 16359 14467
rect 16301 14427 16359 14433
rect 13740 14368 13952 14396
rect 13633 14359 13691 14365
rect 13998 14356 14004 14408
rect 14056 14396 14062 14408
rect 14369 14399 14427 14405
rect 14369 14396 14381 14399
rect 14056 14368 14381 14396
rect 14056 14356 14062 14368
rect 14369 14365 14381 14368
rect 14415 14365 14427 14399
rect 16316 14396 16344 14427
rect 16390 14424 16396 14476
rect 16448 14424 16454 14476
rect 16853 14467 16911 14473
rect 16853 14433 16865 14467
rect 16899 14433 16911 14467
rect 16853 14427 16911 14433
rect 16485 14399 16543 14405
rect 16485 14396 16497 14399
rect 16316 14368 16497 14396
rect 14369 14359 14427 14365
rect 16485 14365 16497 14368
rect 16531 14365 16543 14399
rect 16868 14396 16896 14427
rect 16942 14424 16948 14476
rect 17000 14424 17006 14476
rect 17236 14473 17264 14504
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14433 17279 14467
rect 17328 14464 17356 14560
rect 18414 14532 18420 14544
rect 17696 14504 18420 14532
rect 17696 14473 17724 14504
rect 18414 14492 18420 14504
rect 18472 14492 18478 14544
rect 18524 14504 18920 14532
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 17328 14436 17509 14464
rect 17221 14427 17279 14433
rect 17497 14433 17509 14436
rect 17543 14433 17555 14467
rect 17497 14427 17555 14433
rect 17681 14467 17739 14473
rect 17681 14433 17693 14467
rect 17727 14433 17739 14467
rect 17681 14427 17739 14433
rect 17954 14424 17960 14476
rect 18012 14424 18018 14476
rect 18046 14424 18052 14476
rect 18104 14424 18110 14476
rect 18322 14424 18328 14476
rect 18380 14464 18386 14476
rect 18524 14473 18552 14504
rect 18892 14473 18920 14504
rect 18509 14467 18567 14473
rect 18509 14464 18521 14467
rect 18380 14436 18521 14464
rect 18380 14424 18386 14436
rect 18509 14433 18521 14436
rect 18555 14433 18567 14467
rect 18509 14427 18567 14433
rect 18785 14467 18843 14473
rect 18785 14433 18797 14467
rect 18831 14433 18843 14467
rect 18785 14427 18843 14433
rect 18877 14467 18935 14473
rect 18877 14433 18889 14467
rect 18923 14433 18935 14467
rect 19076 14464 19104 14560
rect 19797 14535 19855 14541
rect 19797 14532 19809 14535
rect 19352 14504 19809 14532
rect 19352 14473 19380 14504
rect 19797 14501 19809 14504
rect 19843 14501 19855 14535
rect 19797 14495 19855 14501
rect 19153 14467 19211 14473
rect 19153 14464 19165 14467
rect 19076 14436 19165 14464
rect 18877 14427 18935 14433
rect 19153 14433 19165 14436
rect 19199 14433 19211 14467
rect 19153 14427 19211 14433
rect 19337 14467 19395 14473
rect 19337 14433 19349 14467
rect 19383 14433 19395 14467
rect 19337 14427 19395 14433
rect 17865 14399 17923 14405
rect 17865 14396 17877 14399
rect 16868 14368 17877 14396
rect 16485 14359 16543 14365
rect 17865 14365 17877 14368
rect 17911 14365 17923 14399
rect 17972 14396 18000 14424
rect 17972 14368 18460 14396
rect 17865 14359 17923 14365
rect 8956 14300 9260 14328
rect 7098 14220 7104 14272
rect 7156 14220 7162 14272
rect 8018 14220 8024 14272
rect 8076 14260 8082 14272
rect 8205 14263 8263 14269
rect 8205 14260 8217 14263
rect 8076 14232 8217 14260
rect 8076 14220 8082 14232
rect 8205 14229 8217 14232
rect 8251 14260 8263 14263
rect 8404 14260 8432 14300
rect 11606 14288 11612 14340
rect 11664 14328 11670 14340
rect 13538 14328 13544 14340
rect 11664 14300 13544 14328
rect 11664 14288 11670 14300
rect 13538 14288 13544 14300
rect 13596 14288 13602 14340
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 14185 14331 14243 14337
rect 14185 14328 14197 14331
rect 13872 14300 14197 14328
rect 13872 14288 13878 14300
rect 14185 14297 14197 14300
rect 14231 14297 14243 14331
rect 14185 14291 14243 14297
rect 17037 14331 17095 14337
rect 17037 14297 17049 14331
rect 17083 14328 17095 14331
rect 18322 14328 18328 14340
rect 17083 14300 18328 14328
rect 17083 14297 17095 14300
rect 17037 14291 17095 14297
rect 18322 14288 18328 14300
rect 18380 14288 18386 14340
rect 18432 14328 18460 14368
rect 18598 14356 18604 14408
rect 18656 14396 18662 14408
rect 18800 14396 18828 14427
rect 19426 14424 19432 14476
rect 19484 14424 19490 14476
rect 19518 14424 19524 14476
rect 19576 14464 19582 14476
rect 19996 14473 20024 14572
rect 21082 14560 21088 14612
rect 21140 14600 21146 14612
rect 21726 14600 21732 14612
rect 21140 14572 21732 14600
rect 21140 14560 21146 14572
rect 21726 14560 21732 14572
rect 21784 14560 21790 14612
rect 22094 14560 22100 14612
rect 22152 14600 22158 14612
rect 22152 14572 22324 14600
rect 22152 14560 22158 14572
rect 20714 14492 20720 14544
rect 20772 14492 20778 14544
rect 21913 14535 21971 14541
rect 21913 14532 21925 14535
rect 21008 14504 21925 14532
rect 19889 14467 19947 14473
rect 19889 14464 19901 14467
rect 19576 14436 19901 14464
rect 19576 14424 19582 14436
rect 19889 14433 19901 14436
rect 19935 14433 19947 14467
rect 19889 14427 19947 14433
rect 19981 14467 20039 14473
rect 19981 14433 19993 14467
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 20441 14467 20499 14473
rect 20441 14433 20453 14467
rect 20487 14433 20499 14467
rect 20732 14463 20760 14492
rect 21008 14473 21036 14504
rect 21913 14501 21925 14504
rect 21959 14501 21971 14535
rect 21913 14495 21971 14501
rect 22189 14535 22247 14541
rect 22189 14501 22201 14535
rect 22235 14501 22247 14535
rect 22189 14495 22247 14501
rect 20993 14467 21051 14473
rect 20441 14427 20499 14433
rect 20717 14457 20775 14463
rect 19536 14396 19564 14424
rect 18656 14368 19564 14396
rect 18656 14356 18662 14368
rect 18782 14328 18788 14340
rect 18432 14300 18788 14328
rect 18782 14288 18788 14300
rect 18840 14288 18846 14340
rect 20456 14328 20484 14427
rect 20717 14423 20729 14457
rect 20763 14423 20775 14457
rect 20993 14433 21005 14467
rect 21039 14433 21051 14467
rect 20993 14427 21051 14433
rect 21453 14467 21511 14473
rect 21453 14433 21465 14467
rect 21499 14433 21511 14467
rect 21453 14427 21511 14433
rect 20717 14417 20775 14423
rect 21468 14396 21496 14427
rect 21542 14424 21548 14476
rect 21600 14424 21606 14476
rect 21818 14424 21824 14476
rect 21876 14464 21882 14476
rect 22005 14467 22063 14473
rect 22005 14464 22017 14467
rect 21876 14436 22017 14464
rect 21876 14424 21882 14436
rect 22005 14433 22017 14436
rect 22051 14433 22063 14467
rect 22005 14427 22063 14433
rect 22094 14396 22100 14408
rect 21468 14368 22100 14396
rect 22094 14356 22100 14368
rect 22152 14356 22158 14408
rect 20714 14328 20720 14340
rect 20456 14300 20720 14328
rect 20714 14288 20720 14300
rect 20772 14288 20778 14340
rect 21726 14288 21732 14340
rect 21784 14328 21790 14340
rect 22204 14328 22232 14495
rect 22296 14473 22324 14572
rect 22554 14560 22560 14612
rect 22612 14560 22618 14612
rect 22830 14560 22836 14612
rect 22888 14600 22894 14612
rect 22888 14572 23980 14600
rect 22888 14560 22894 14572
rect 22572 14532 22600 14560
rect 22388 14504 22600 14532
rect 22640 14535 22698 14541
rect 22388 14473 22416 14504
rect 22640 14501 22652 14535
rect 22686 14532 22698 14535
rect 23106 14532 23112 14544
rect 22686 14504 23112 14532
rect 22686 14501 22698 14504
rect 22640 14495 22698 14501
rect 23106 14492 23112 14504
rect 23164 14492 23170 14544
rect 23952 14532 23980 14572
rect 24026 14560 24032 14612
rect 24084 14560 24090 14612
rect 24118 14560 24124 14612
rect 24176 14600 24182 14612
rect 24302 14600 24308 14612
rect 24176 14572 24308 14600
rect 24176 14560 24182 14572
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 24578 14560 24584 14612
rect 24636 14600 24642 14612
rect 25409 14603 25467 14609
rect 25409 14600 25421 14603
rect 24636 14572 25421 14600
rect 24636 14560 24642 14572
rect 25409 14569 25421 14572
rect 25455 14569 25467 14603
rect 25409 14563 25467 14569
rect 25682 14560 25688 14612
rect 25740 14560 25746 14612
rect 25774 14560 25780 14612
rect 25832 14560 25838 14612
rect 25792 14532 25820 14560
rect 23952 14504 24072 14532
rect 22281 14467 22339 14473
rect 22281 14433 22293 14467
rect 22327 14433 22339 14467
rect 22281 14427 22339 14433
rect 22373 14467 22431 14473
rect 22373 14433 22385 14467
rect 22419 14433 22431 14467
rect 23934 14464 23940 14476
rect 22373 14427 22431 14433
rect 22480 14436 23940 14464
rect 22480 14396 22508 14436
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 21784 14300 22232 14328
rect 22296 14368 22508 14396
rect 24044 14396 24072 14504
rect 24412 14504 25084 14532
rect 24412 14476 24440 14504
rect 24118 14424 24124 14476
rect 24176 14424 24182 14476
rect 24213 14467 24271 14473
rect 24213 14433 24225 14467
rect 24259 14433 24271 14467
rect 24213 14427 24271 14433
rect 24228 14396 24256 14427
rect 24394 14424 24400 14476
rect 24452 14424 24458 14476
rect 24673 14467 24731 14473
rect 24673 14433 24685 14467
rect 24719 14433 24731 14467
rect 24673 14427 24731 14433
rect 24044 14368 24256 14396
rect 24688 14396 24716 14427
rect 24946 14424 24952 14476
rect 25004 14424 25010 14476
rect 25056 14473 25084 14504
rect 25424 14504 25636 14532
rect 25792 14504 25912 14532
rect 25049 14467 25107 14473
rect 25049 14433 25061 14467
rect 25095 14464 25107 14467
rect 25424 14464 25452 14504
rect 25095 14462 25176 14464
rect 25240 14462 25452 14464
rect 25095 14436 25452 14462
rect 25095 14433 25107 14436
rect 25148 14434 25268 14436
rect 25049 14427 25107 14433
rect 25498 14424 25504 14476
rect 25556 14424 25562 14476
rect 25608 14464 25636 14504
rect 25774 14464 25780 14476
rect 25608 14436 25780 14464
rect 25774 14424 25780 14436
rect 25832 14424 25838 14476
rect 25884 14473 25912 14504
rect 25869 14467 25927 14473
rect 25869 14433 25881 14467
rect 25915 14433 25927 14467
rect 25869 14427 25927 14433
rect 24808 14396 24814 14408
rect 24688 14368 24814 14396
rect 21784 14288 21790 14300
rect 8251 14232 8432 14260
rect 8251 14229 8263 14232
rect 8205 14223 8263 14229
rect 8478 14220 8484 14272
rect 8536 14220 8542 14272
rect 8757 14263 8815 14269
rect 8757 14229 8769 14263
rect 8803 14260 8815 14263
rect 9490 14260 9496 14272
rect 8803 14232 9496 14260
rect 8803 14229 8815 14232
rect 8757 14223 8815 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 11054 14220 11060 14272
rect 11112 14220 11118 14272
rect 13722 14220 13728 14272
rect 13780 14260 13786 14272
rect 13909 14263 13967 14269
rect 13909 14260 13921 14263
rect 13780 14232 13921 14260
rect 13780 14220 13786 14232
rect 13909 14229 13921 14232
rect 13955 14229 13967 14263
rect 13909 14223 13967 14229
rect 16206 14220 16212 14272
rect 16264 14220 16270 14272
rect 17310 14220 17316 14272
rect 17368 14220 17374 14272
rect 17494 14220 17500 14272
rect 17552 14260 17558 14272
rect 18141 14263 18199 14269
rect 18141 14260 18153 14263
rect 17552 14232 18153 14260
rect 17552 14220 17558 14232
rect 18141 14229 18153 14232
rect 18187 14229 18199 14263
rect 18141 14223 18199 14229
rect 18414 14220 18420 14272
rect 18472 14220 18478 14272
rect 18506 14220 18512 14272
rect 18564 14260 18570 14272
rect 18693 14263 18751 14269
rect 18693 14260 18705 14263
rect 18564 14232 18705 14260
rect 18564 14220 18570 14232
rect 18693 14229 18705 14232
rect 18739 14229 18751 14263
rect 18693 14223 18751 14229
rect 19242 14220 19248 14272
rect 19300 14220 19306 14272
rect 19521 14263 19579 14269
rect 19521 14229 19533 14263
rect 19567 14260 19579 14263
rect 20073 14263 20131 14269
rect 20073 14260 20085 14263
rect 19567 14232 20085 14260
rect 19567 14229 19579 14232
rect 19521 14223 19579 14229
rect 20073 14229 20085 14232
rect 20119 14229 20131 14263
rect 20073 14223 20131 14229
rect 20346 14220 20352 14272
rect 20404 14220 20410 14272
rect 20438 14220 20444 14272
rect 20496 14260 20502 14272
rect 20625 14263 20683 14269
rect 20625 14260 20637 14263
rect 20496 14232 20637 14260
rect 20496 14220 20502 14232
rect 20625 14229 20637 14232
rect 20671 14229 20683 14263
rect 20625 14223 20683 14229
rect 20901 14263 20959 14269
rect 20901 14229 20913 14263
rect 20947 14260 20959 14263
rect 21174 14260 21180 14272
rect 20947 14232 21180 14260
rect 20947 14229 20959 14232
rect 20901 14223 20959 14229
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 21361 14263 21419 14269
rect 21361 14229 21373 14263
rect 21407 14260 21419 14263
rect 21450 14260 21456 14272
rect 21407 14232 21456 14260
rect 21407 14229 21419 14232
rect 21361 14223 21419 14229
rect 21450 14220 21456 14232
rect 21508 14220 21514 14272
rect 21637 14263 21695 14269
rect 21637 14229 21649 14263
rect 21683 14260 21695 14263
rect 22296 14260 22324 14368
rect 24808 14356 24814 14368
rect 24866 14356 24872 14408
rect 25682 14356 25688 14408
rect 25740 14396 25746 14408
rect 25961 14399 26019 14405
rect 25961 14396 25973 14399
rect 25740 14368 25973 14396
rect 25740 14356 25746 14368
rect 25961 14365 25973 14368
rect 26007 14365 26019 14399
rect 25961 14359 26019 14365
rect 24305 14331 24363 14337
rect 24305 14328 24317 14331
rect 23391 14300 24317 14328
rect 21683 14232 22324 14260
rect 21683 14229 21695 14232
rect 21637 14223 21695 14229
rect 22370 14220 22376 14272
rect 22428 14260 22434 14272
rect 23391 14260 23419 14300
rect 24305 14297 24317 14300
rect 24351 14297 24363 14331
rect 24946 14328 24952 14340
rect 24305 14291 24363 14297
rect 24872 14300 24952 14328
rect 22428 14232 23419 14260
rect 23753 14263 23811 14269
rect 22428 14220 22434 14232
rect 23753 14229 23765 14263
rect 23799 14260 23811 14263
rect 24210 14260 24216 14272
rect 23799 14232 24216 14260
rect 23799 14229 23811 14232
rect 23753 14223 23811 14229
rect 24210 14220 24216 14232
rect 24268 14220 24274 14272
rect 24578 14220 24584 14272
rect 24636 14220 24642 14272
rect 24872 14269 24900 14300
rect 24946 14288 24952 14300
rect 25004 14288 25010 14340
rect 24857 14263 24915 14269
rect 24857 14229 24869 14263
rect 24903 14229 24915 14263
rect 24857 14223 24915 14229
rect 25130 14220 25136 14272
rect 25188 14220 25194 14272
rect 552 14170 31372 14192
rect 552 14118 4250 14170
rect 4302 14118 4314 14170
rect 4366 14118 4378 14170
rect 4430 14118 4442 14170
rect 4494 14118 4506 14170
rect 4558 14118 11955 14170
rect 12007 14118 12019 14170
rect 12071 14118 12083 14170
rect 12135 14118 12147 14170
rect 12199 14118 12211 14170
rect 12263 14118 19660 14170
rect 19712 14118 19724 14170
rect 19776 14118 19788 14170
rect 19840 14118 19852 14170
rect 19904 14118 19916 14170
rect 19968 14118 27365 14170
rect 27417 14118 27429 14170
rect 27481 14118 27493 14170
rect 27545 14118 27557 14170
rect 27609 14118 27621 14170
rect 27673 14118 31372 14170
rect 552 14096 31372 14118
rect 7009 14059 7067 14065
rect 7009 14025 7021 14059
rect 7055 14056 7067 14059
rect 7834 14056 7840 14068
rect 7055 14028 7840 14056
rect 7055 14025 7067 14028
rect 7009 14019 7067 14025
rect 7834 14016 7840 14028
rect 7892 14016 7898 14068
rect 7926 14016 7932 14068
rect 7984 14056 7990 14068
rect 8113 14059 8171 14065
rect 8113 14056 8125 14059
rect 7984 14028 8125 14056
rect 7984 14016 7990 14028
rect 8113 14025 8125 14028
rect 8159 14025 8171 14059
rect 8113 14019 8171 14025
rect 8570 14016 8576 14068
rect 8628 14016 8634 14068
rect 8938 14056 8944 14068
rect 8680 14028 8944 14056
rect 7190 13948 7196 14000
rect 7248 13948 7254 14000
rect 7285 13991 7343 13997
rect 7285 13957 7297 13991
rect 7331 13988 7343 13991
rect 8588 13988 8616 14016
rect 7331 13960 8616 13988
rect 7331 13957 7343 13960
rect 7285 13951 7343 13957
rect 7098 13812 7104 13864
rect 7156 13812 7162 13864
rect 7208 13861 7236 13948
rect 7466 13880 7472 13932
rect 7524 13880 7530 13932
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 8110 13920 8116 13932
rect 7607 13892 8116 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 8294 13880 8300 13932
rect 8352 13880 8358 13932
rect 8680 13929 8708 14028
rect 8938 14016 8944 14028
rect 8996 14056 9002 14068
rect 9766 14056 9772 14068
rect 8996 14028 9772 14056
rect 8996 14016 9002 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 9858 14016 9864 14068
rect 9916 14056 9922 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 9916 14028 10057 14056
rect 9916 14016 9922 14028
rect 10045 14025 10057 14028
rect 10091 14025 10103 14059
rect 10045 14019 10103 14025
rect 10226 14016 10232 14068
rect 10284 14056 10290 14068
rect 10284 14028 11652 14056
rect 10284 14016 10290 14028
rect 9784 13988 9812 14016
rect 10134 13988 10140 14000
rect 9784 13960 10140 13988
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 10502 13948 10508 14000
rect 10560 13948 10566 14000
rect 10778 13948 10784 14000
rect 10836 13988 10842 14000
rect 11624 13997 11652 14028
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11756 14028 12173 14056
rect 11756 14016 11762 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 12483 14028 14136 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 11333 13991 11391 13997
rect 11333 13988 11345 13991
rect 10836 13960 11345 13988
rect 10836 13948 10842 13960
rect 11333 13957 11345 13960
rect 11379 13957 11391 13991
rect 11333 13951 11391 13957
rect 11609 13991 11667 13997
rect 11609 13957 11621 13991
rect 11655 13957 11667 13991
rect 11609 13951 11667 13957
rect 11790 13948 11796 14000
rect 11848 13988 11854 14000
rect 12989 13991 13047 13997
rect 12989 13988 13001 13991
rect 11848 13960 13001 13988
rect 11848 13948 11854 13960
rect 12989 13957 13001 13960
rect 13035 13957 13047 13991
rect 12989 13951 13047 13957
rect 13265 13991 13323 13997
rect 13265 13957 13277 13991
rect 13311 13988 13323 13991
rect 13446 13988 13452 14000
rect 13311 13960 13452 13988
rect 13311 13957 13323 13960
rect 13265 13951 13323 13957
rect 13446 13948 13452 13960
rect 13504 13948 13510 14000
rect 13817 13991 13875 13997
rect 13817 13957 13829 13991
rect 13863 13988 13875 13991
rect 13906 13988 13912 14000
rect 13863 13960 13912 13988
rect 13863 13957 13875 13960
rect 13817 13951 13875 13957
rect 13906 13948 13912 13960
rect 13964 13948 13970 14000
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13889 8723 13923
rect 11882 13920 11888 13932
rect 8665 13883 8723 13889
rect 10612 13892 11100 13920
rect 7193 13855 7251 13861
rect 7193 13821 7205 13855
rect 7239 13821 7251 13855
rect 7193 13815 7251 13821
rect 7374 13812 7380 13864
rect 7432 13855 7438 13864
rect 7432 13812 7443 13855
rect 7385 13809 7443 13812
rect 7484 13716 7512 13880
rect 7650 13812 7656 13864
rect 7708 13812 7714 13864
rect 7926 13812 7932 13864
rect 7984 13812 7990 13864
rect 8021 13855 8079 13861
rect 8021 13821 8033 13855
rect 8067 13852 8079 13855
rect 8202 13852 8208 13864
rect 8067 13824 8208 13852
rect 8067 13821 8079 13824
rect 8021 13815 8079 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 7558 13744 7564 13796
rect 7616 13784 7622 13796
rect 8312 13784 8340 13880
rect 8389 13855 8447 13861
rect 8389 13821 8401 13855
rect 8435 13852 8447 13855
rect 8570 13852 8576 13864
rect 8435 13824 8576 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 8570 13812 8576 13824
rect 8628 13812 8634 13864
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 9306 13852 9312 13864
rect 8812 13824 9312 13852
rect 8812 13812 8818 13824
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 10612 13861 10640 13892
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13821 10655 13855
rect 10597 13815 10655 13821
rect 10686 13812 10692 13864
rect 10744 13812 10750 13864
rect 10781 13855 10839 13861
rect 10781 13821 10793 13855
rect 10827 13852 10839 13855
rect 10870 13852 10876 13864
rect 10827 13824 10876 13852
rect 10827 13821 10839 13824
rect 10781 13815 10839 13821
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 10965 13855 11023 13861
rect 10965 13821 10977 13855
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 8910 13787 8968 13793
rect 8910 13784 8922 13787
rect 7616 13756 8248 13784
rect 8312 13756 8922 13784
rect 7616 13744 7622 13756
rect 7837 13719 7895 13725
rect 7837 13716 7849 13719
rect 7484 13688 7849 13716
rect 7837 13685 7849 13688
rect 7883 13685 7895 13719
rect 8220 13716 8248 13756
rect 8910 13753 8922 13756
rect 8956 13753 8968 13787
rect 8910 13747 8968 13753
rect 10134 13744 10140 13796
rect 10192 13784 10198 13796
rect 10980 13784 11008 13815
rect 11072 13793 11100 13892
rect 11440 13892 11888 13920
rect 11440 13861 11468 13892
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 12342 13880 12348 13932
rect 12400 13920 12406 13932
rect 12713 13923 12771 13929
rect 12713 13920 12725 13923
rect 12400 13892 12725 13920
rect 12400 13880 12406 13892
rect 12713 13889 12725 13892
rect 12759 13889 12771 13923
rect 13538 13920 13544 13932
rect 12713 13883 12771 13889
rect 12820 13892 13544 13920
rect 11425 13855 11483 13861
rect 11425 13821 11437 13855
rect 11471 13821 11483 13855
rect 11425 13815 11483 13821
rect 11606 13812 11612 13864
rect 11664 13852 11670 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11664 13824 11713 13852
rect 11664 13812 11670 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 11977 13855 12035 13861
rect 11977 13821 11989 13855
rect 12023 13821 12035 13855
rect 11977 13815 12035 13821
rect 10192 13756 11008 13784
rect 11057 13787 11115 13793
rect 10192 13744 10198 13756
rect 11057 13753 11069 13787
rect 11103 13784 11115 13787
rect 11624 13784 11652 13812
rect 11103 13756 11652 13784
rect 11992 13784 12020 13815
rect 12066 13812 12072 13864
rect 12124 13812 12130 13864
rect 12820 13861 12848 13892
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14108 13920 14136 14028
rect 14182 14016 14188 14068
rect 14240 14056 14246 14068
rect 14240 14028 15424 14056
rect 14240 14016 14246 14028
rect 15396 13997 15424 14028
rect 17310 14016 17316 14068
rect 17368 14016 17374 14068
rect 17865 14059 17923 14065
rect 17865 14025 17877 14059
rect 17911 14056 17923 14059
rect 17954 14056 17960 14068
rect 17911 14028 17960 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 18046 14016 18052 14068
rect 18104 14056 18110 14068
rect 18141 14059 18199 14065
rect 18141 14056 18153 14059
rect 18104 14028 18153 14056
rect 18104 14016 18110 14028
rect 18141 14025 18153 14028
rect 18187 14025 18199 14059
rect 18141 14019 18199 14025
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 20625 14059 20683 14065
rect 20625 14056 20637 14059
rect 19300 14028 20637 14056
rect 19300 14016 19306 14028
rect 20625 14025 20637 14028
rect 20671 14025 20683 14059
rect 20625 14019 20683 14025
rect 20714 14016 20720 14068
rect 20772 14056 20778 14068
rect 20901 14059 20959 14065
rect 20901 14056 20913 14059
rect 20772 14028 20913 14056
rect 20772 14016 20778 14028
rect 20901 14025 20913 14028
rect 20947 14025 20959 14059
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 20901 14019 20959 14025
rect 21008 14028 21465 14056
rect 15381 13991 15439 13997
rect 15381 13957 15393 13991
rect 15427 13957 15439 13991
rect 16390 13988 16396 14000
rect 15381 13951 15439 13957
rect 15856 13960 16396 13988
rect 14108 13892 14228 13920
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13852 12587 13855
rect 12805 13855 12863 13861
rect 12575 13824 12756 13852
rect 12575 13821 12587 13824
rect 12529 13815 12587 13821
rect 12158 13784 12164 13796
rect 11992 13756 12164 13784
rect 11103 13753 11115 13756
rect 11057 13747 11115 13753
rect 12158 13744 12164 13756
rect 12216 13744 12222 13796
rect 12728 13784 12756 13824
rect 12805 13821 12817 13855
rect 12851 13852 12863 13855
rect 12986 13852 12992 13864
rect 12851 13824 12992 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 12986 13812 12992 13824
rect 13044 13812 13050 13864
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 13357 13855 13415 13861
rect 13357 13821 13369 13855
rect 13403 13852 13415 13855
rect 13722 13852 13728 13864
rect 13403 13824 13728 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 13096 13784 13124 13815
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 14200 13852 14228 13892
rect 14200 13824 14596 13852
rect 13630 13784 13636 13796
rect 12728 13756 12848 13784
rect 13096 13756 13636 13784
rect 8481 13719 8539 13725
rect 8481 13716 8493 13719
rect 8220 13688 8493 13716
rect 7837 13679 7895 13685
rect 8481 13685 8493 13688
rect 8527 13685 8539 13719
rect 8481 13679 8539 13685
rect 9214 13676 9220 13728
rect 9272 13716 9278 13728
rect 10042 13716 10048 13728
rect 9272 13688 10048 13716
rect 9272 13676 9278 13688
rect 10042 13676 10048 13688
rect 10100 13716 10106 13728
rect 11514 13716 11520 13728
rect 10100 13688 11520 13716
rect 10100 13676 10106 13688
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 11885 13719 11943 13725
rect 11885 13685 11897 13719
rect 11931 13716 11943 13719
rect 12618 13716 12624 13728
rect 11931 13688 12624 13716
rect 11931 13685 11943 13688
rect 11885 13679 11943 13685
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 12820 13716 12848 13756
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 14458 13784 14464 13796
rect 13740 13756 14464 13784
rect 13740 13716 13768 13756
rect 14458 13744 14464 13756
rect 14516 13744 14522 13796
rect 14568 13784 14596 13824
rect 14642 13812 14648 13864
rect 14700 13852 14706 13864
rect 15197 13855 15255 13861
rect 14700 13824 15056 13852
rect 14700 13812 14706 13824
rect 14930 13787 14988 13793
rect 14930 13784 14942 13787
rect 14568 13756 14942 13784
rect 14930 13753 14942 13756
rect 14976 13753 14988 13787
rect 15028 13784 15056 13824
rect 15197 13821 15209 13855
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 15212 13784 15240 13815
rect 15286 13812 15292 13864
rect 15344 13852 15350 13864
rect 15856 13861 15884 13960
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 17328 13988 17356 14016
rect 17328 13960 18460 13988
rect 18432 13929 18460 13960
rect 19518 13948 19524 14000
rect 19576 13988 19582 14000
rect 19981 13991 20039 13997
rect 19981 13988 19993 13991
rect 19576 13960 19993 13988
rect 19576 13948 19582 13960
rect 19981 13957 19993 13960
rect 20027 13957 20039 13991
rect 19981 13951 20039 13957
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16577 13923 16635 13929
rect 16577 13920 16589 13923
rect 16071 13892 16589 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 16577 13889 16589 13892
rect 16623 13889 16635 13923
rect 17589 13923 17647 13929
rect 17589 13920 17601 13923
rect 16577 13883 16635 13889
rect 17144 13892 17601 13920
rect 15473 13855 15531 13861
rect 15473 13852 15485 13855
rect 15344 13824 15485 13852
rect 15344 13812 15350 13824
rect 15473 13821 15485 13824
rect 15519 13821 15531 13855
rect 15473 13815 15531 13821
rect 15841 13855 15899 13861
rect 15841 13821 15853 13855
rect 15887 13821 15899 13855
rect 15841 13815 15899 13821
rect 15856 13784 15884 13815
rect 15930 13812 15936 13864
rect 15988 13812 15994 13864
rect 17144 13861 17172 13892
rect 17589 13889 17601 13892
rect 17635 13889 17647 13923
rect 17589 13883 17647 13889
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 18782 13880 18788 13932
rect 18840 13920 18846 13932
rect 21008 13920 21036 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 23750 14056 23756 14068
rect 21453 14019 21511 14025
rect 22066 14028 23756 14056
rect 21177 13991 21235 13997
rect 21177 13957 21189 13991
rect 21223 13988 21235 13991
rect 22066 13988 22094 14028
rect 23750 14016 23756 14028
rect 23808 14016 23814 14068
rect 23842 14016 23848 14068
rect 23900 14056 23906 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 23900 14028 25053 14056
rect 23900 14016 23906 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25041 14019 25099 14025
rect 25130 14016 25136 14068
rect 25188 14016 25194 14068
rect 25314 14016 25320 14068
rect 25372 14016 25378 14068
rect 25590 14016 25596 14068
rect 25648 14016 25654 14068
rect 26142 14016 26148 14068
rect 26200 14016 26206 14068
rect 26418 14016 26424 14068
rect 26476 14016 26482 14068
rect 21223 13960 22094 13988
rect 21223 13957 21235 13960
rect 21177 13951 21235 13957
rect 23474 13948 23480 14000
rect 23532 13988 23538 14000
rect 23569 13991 23627 13997
rect 23569 13988 23581 13991
rect 23532 13960 23581 13988
rect 23532 13948 23538 13960
rect 23569 13957 23581 13960
rect 23615 13957 23627 13991
rect 23569 13951 23627 13957
rect 24213 13991 24271 13997
rect 24213 13957 24225 13991
rect 24259 13988 24271 13991
rect 24762 13988 24768 14000
rect 24259 13960 24768 13988
rect 24259 13957 24271 13960
rect 24213 13951 24271 13957
rect 24762 13948 24768 13960
rect 24820 13948 24826 14000
rect 21450 13920 21456 13932
rect 18840 13892 21036 13920
rect 21284 13892 21456 13920
rect 18840 13880 18846 13892
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 16301 13855 16359 13861
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 16485 13855 16543 13861
rect 16485 13852 16497 13855
rect 16347 13824 16497 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 16485 13821 16497 13824
rect 16531 13821 16543 13855
rect 16485 13815 16543 13821
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13821 17187 13855
rect 17129 13815 17187 13821
rect 15028 13756 15240 13784
rect 15304 13756 15884 13784
rect 16224 13784 16252 13815
rect 17218 13812 17224 13864
rect 17276 13812 17282 13864
rect 17678 13812 17684 13864
rect 17736 13812 17742 13864
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13852 18015 13855
rect 18046 13852 18052 13864
rect 18003 13824 18052 13852
rect 18003 13821 18015 13824
rect 17957 13815 18015 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18230 13812 18236 13864
rect 18288 13812 18294 13864
rect 18322 13812 18328 13864
rect 18380 13812 18386 13864
rect 20732 13861 20760 13892
rect 18693 13855 18751 13861
rect 18693 13821 18705 13855
rect 18739 13821 18751 13855
rect 18693 13815 18751 13821
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 20809 13855 20867 13861
rect 20809 13821 20821 13855
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 16390 13784 16396 13796
rect 16224 13756 16396 13784
rect 14930 13747 14988 13753
rect 12820 13688 13768 13716
rect 13906 13676 13912 13728
rect 13964 13716 13970 13728
rect 14734 13716 14740 13728
rect 13964 13688 14740 13716
rect 13964 13676 13970 13688
rect 14734 13676 14740 13688
rect 14792 13716 14798 13728
rect 15304 13716 15332 13756
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 16942 13744 16948 13796
rect 17000 13784 17006 13796
rect 18708 13784 18736 13815
rect 17000 13756 18736 13784
rect 17000 13744 17006 13756
rect 20254 13744 20260 13796
rect 20312 13784 20318 13796
rect 20824 13784 20852 13815
rect 20990 13812 20996 13864
rect 21048 13852 21054 13864
rect 21284 13861 21312 13892
rect 21450 13880 21456 13892
rect 21508 13880 21514 13932
rect 25148 13920 25176 14016
rect 25222 13948 25228 14000
rect 25280 13988 25286 14000
rect 25869 13991 25927 13997
rect 25869 13988 25881 13991
rect 25280 13960 25881 13988
rect 25280 13948 25286 13960
rect 25869 13957 25881 13960
rect 25915 13957 25927 13991
rect 25869 13951 25927 13957
rect 25148 13892 26096 13920
rect 21269 13855 21327 13861
rect 21048 13824 21220 13852
rect 21048 13812 21054 13824
rect 20312 13756 20852 13784
rect 21192 13784 21220 13824
rect 21269 13821 21281 13855
rect 21315 13821 21327 13855
rect 21269 13815 21327 13821
rect 21361 13855 21419 13861
rect 21361 13821 21373 13855
rect 21407 13821 21419 13855
rect 21361 13815 21419 13821
rect 21376 13784 21404 13815
rect 21726 13812 21732 13864
rect 21784 13852 21790 13864
rect 21821 13855 21879 13861
rect 21821 13852 21833 13855
rect 21784 13824 21833 13852
rect 21784 13812 21790 13824
rect 21821 13821 21833 13824
rect 21867 13821 21879 13855
rect 21821 13815 21879 13821
rect 21913 13855 21971 13861
rect 21913 13821 21925 13855
rect 21959 13821 21971 13855
rect 21913 13815 21971 13821
rect 21192 13756 21404 13784
rect 20312 13744 20318 13756
rect 21450 13744 21456 13796
rect 21508 13784 21514 13796
rect 21928 13784 21956 13815
rect 22186 13812 22192 13864
rect 22244 13812 22250 13864
rect 22278 13812 22284 13864
rect 22336 13852 22342 13864
rect 22456 13855 22514 13861
rect 22336 13824 22416 13852
rect 22336 13812 22342 13824
rect 21508 13756 21956 13784
rect 22388 13784 22416 13824
rect 22456 13821 22468 13855
rect 22502 13852 22514 13855
rect 23290 13852 23296 13864
rect 22502 13824 23296 13852
rect 22502 13821 22514 13824
rect 22456 13815 22514 13821
rect 23290 13812 23296 13824
rect 23348 13812 23354 13864
rect 24029 13855 24087 13861
rect 24029 13821 24041 13855
rect 24075 13821 24087 13855
rect 24029 13815 24087 13821
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13852 24179 13855
rect 24394 13852 24400 13864
rect 24167 13824 24400 13852
rect 24167 13821 24179 13824
rect 24121 13815 24179 13821
rect 23937 13787 23995 13793
rect 23937 13784 23949 13787
rect 22388 13756 23949 13784
rect 21508 13744 21514 13756
rect 23937 13753 23949 13756
rect 23983 13753 23995 13787
rect 24044 13784 24072 13815
rect 24210 13784 24216 13796
rect 24044 13756 24216 13784
rect 23937 13747 23995 13753
rect 24210 13744 24216 13756
rect 24268 13744 24274 13796
rect 14792 13688 15332 13716
rect 14792 13676 14798 13688
rect 15470 13676 15476 13728
rect 15528 13716 15534 13728
rect 15749 13719 15807 13725
rect 15749 13716 15761 13719
rect 15528 13688 15761 13716
rect 15528 13676 15534 13688
rect 15749 13685 15761 13688
rect 15795 13685 15807 13719
rect 15749 13679 15807 13685
rect 17037 13719 17095 13725
rect 17037 13685 17049 13719
rect 17083 13716 17095 13719
rect 17126 13716 17132 13728
rect 17083 13688 17132 13716
rect 17083 13685 17095 13688
rect 17037 13679 17095 13685
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 17313 13719 17371 13725
rect 17313 13685 17325 13719
rect 17359 13716 17371 13719
rect 19334 13716 19340 13728
rect 17359 13688 19340 13716
rect 17359 13685 17371 13688
rect 17313 13679 17371 13685
rect 19334 13676 19340 13688
rect 19392 13676 19398 13728
rect 21726 13676 21732 13728
rect 21784 13676 21790 13728
rect 22002 13676 22008 13728
rect 22060 13676 22066 13728
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 24320 13716 24348 13824
rect 24394 13812 24400 13824
rect 24452 13812 24458 13864
rect 24486 13812 24492 13864
rect 24544 13812 24550 13864
rect 24581 13855 24639 13861
rect 24581 13821 24593 13855
rect 24627 13852 24639 13855
rect 24627 13824 24808 13852
rect 24627 13821 24639 13824
rect 24581 13815 24639 13821
rect 24504 13784 24532 13812
rect 24780 13784 24808 13824
rect 24854 13812 24860 13864
rect 24912 13812 24918 13864
rect 25133 13855 25191 13861
rect 25133 13821 25145 13855
rect 25179 13821 25191 13855
rect 25133 13815 25191 13821
rect 25409 13855 25467 13861
rect 25409 13821 25421 13855
rect 25455 13852 25467 13855
rect 25590 13852 25596 13864
rect 25455 13824 25596 13852
rect 25455 13821 25467 13824
rect 25409 13815 25467 13821
rect 25148 13784 25176 13815
rect 25590 13812 25596 13824
rect 25648 13812 25654 13864
rect 25685 13855 25743 13861
rect 25685 13821 25697 13855
rect 25731 13852 25743 13855
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 25731 13824 25789 13852
rect 25731 13821 25743 13824
rect 25685 13815 25743 13821
rect 25777 13821 25789 13824
rect 25823 13852 25835 13855
rect 25866 13852 25872 13864
rect 25823 13824 25872 13852
rect 25823 13821 25835 13824
rect 25777 13815 25835 13821
rect 25866 13812 25872 13824
rect 25924 13812 25930 13864
rect 26068 13861 26096 13892
rect 26053 13855 26111 13861
rect 26053 13821 26065 13855
rect 26099 13821 26111 13855
rect 26053 13815 26111 13821
rect 26326 13812 26332 13864
rect 26384 13812 26390 13864
rect 26602 13812 26608 13864
rect 26660 13812 26666 13864
rect 24504 13756 24624 13784
rect 24780 13756 25084 13784
rect 25148 13756 25728 13784
rect 24489 13719 24547 13725
rect 24489 13716 24501 13719
rect 22152 13688 24501 13716
rect 22152 13676 22158 13688
rect 24489 13685 24501 13688
rect 24535 13685 24547 13719
rect 24596 13716 24624 13756
rect 24765 13719 24823 13725
rect 24765 13716 24777 13719
rect 24596 13688 24777 13716
rect 24489 13679 24547 13685
rect 24765 13685 24777 13688
rect 24811 13685 24823 13719
rect 25056 13716 25084 13756
rect 25700 13728 25728 13756
rect 25406 13716 25412 13728
rect 25056 13688 25412 13716
rect 24765 13679 24823 13685
rect 25406 13676 25412 13688
rect 25464 13676 25470 13728
rect 25682 13676 25688 13728
rect 25740 13676 25746 13728
rect 26694 13676 26700 13728
rect 26752 13676 26758 13728
rect 552 13626 31531 13648
rect 552 13574 8102 13626
rect 8154 13574 8166 13626
rect 8218 13574 8230 13626
rect 8282 13574 8294 13626
rect 8346 13574 8358 13626
rect 8410 13574 15807 13626
rect 15859 13574 15871 13626
rect 15923 13574 15935 13626
rect 15987 13574 15999 13626
rect 16051 13574 16063 13626
rect 16115 13574 23512 13626
rect 23564 13574 23576 13626
rect 23628 13574 23640 13626
rect 23692 13574 23704 13626
rect 23756 13574 23768 13626
rect 23820 13574 31217 13626
rect 31269 13574 31281 13626
rect 31333 13574 31345 13626
rect 31397 13574 31409 13626
rect 31461 13574 31473 13626
rect 31525 13574 31531 13626
rect 552 13552 31531 13574
rect 7926 13472 7932 13524
rect 7984 13512 7990 13524
rect 8386 13512 8392 13524
rect 7984 13484 8392 13512
rect 7984 13472 7990 13484
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8478 13472 8484 13524
rect 8536 13472 8542 13524
rect 8662 13472 8668 13524
rect 8720 13472 8726 13524
rect 8772 13484 9536 13512
rect 7650 13404 7656 13456
rect 7708 13404 7714 13456
rect 8496 13444 8524 13472
rect 7760 13416 8524 13444
rect 7469 13379 7527 13385
rect 7469 13345 7481 13379
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13376 7619 13379
rect 7668 13376 7696 13404
rect 7760 13385 7788 13416
rect 7607 13348 7696 13376
rect 7745 13379 7803 13385
rect 7607 13345 7619 13348
rect 7561 13339 7619 13345
rect 7745 13345 7757 13379
rect 7791 13345 7803 13379
rect 7745 13339 7803 13345
rect 7484 13240 7512 13339
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 8021 13379 8079 13385
rect 8021 13376 8033 13379
rect 7984 13348 8033 13376
rect 7984 13336 7990 13348
rect 8021 13345 8033 13348
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 8110 13336 8116 13388
rect 8168 13336 8174 13388
rect 8205 13379 8263 13385
rect 8205 13345 8217 13379
rect 8251 13376 8263 13379
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 8251 13348 8401 13376
rect 8251 13345 8263 13348
rect 8205 13339 8263 13345
rect 8389 13345 8401 13348
rect 8435 13345 8447 13379
rect 8389 13339 8447 13345
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13308 7711 13311
rect 8680 13308 8708 13472
rect 7699 13280 8708 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 8018 13240 8024 13252
rect 7484 13212 8024 13240
rect 8018 13200 8024 13212
rect 8076 13240 8082 13252
rect 8772 13240 8800 13484
rect 9122 13404 9128 13456
rect 9180 13404 9186 13456
rect 8849 13379 8907 13385
rect 8849 13345 8861 13379
rect 8895 13345 8907 13379
rect 9140 13375 9168 13404
rect 8849 13339 8907 13345
rect 9125 13369 9183 13375
rect 8076 13212 8800 13240
rect 8864 13240 8892 13339
rect 9125 13335 9137 13369
rect 9171 13335 9183 13369
rect 9214 13336 9220 13388
rect 9272 13336 9278 13388
rect 9508 13385 9536 13484
rect 9582 13472 9588 13524
rect 9640 13472 9646 13524
rect 10134 13472 10140 13524
rect 10192 13472 10198 13524
rect 10413 13515 10471 13521
rect 10413 13481 10425 13515
rect 10459 13512 10471 13515
rect 10686 13512 10692 13524
rect 10459 13484 10692 13512
rect 10459 13481 10471 13484
rect 10413 13475 10471 13481
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 11054 13512 11060 13524
rect 10796 13484 11060 13512
rect 10796 13444 10824 13484
rect 11054 13472 11060 13484
rect 11112 13472 11118 13524
rect 12526 13512 12532 13524
rect 11155 13484 12532 13512
rect 11155 13444 11183 13484
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 13354 13472 13360 13524
rect 13412 13472 13418 13524
rect 13725 13515 13783 13521
rect 13725 13481 13737 13515
rect 13771 13512 13783 13515
rect 13906 13512 13912 13524
rect 13771 13484 13912 13512
rect 13771 13481 13783 13484
rect 13725 13475 13783 13481
rect 13906 13472 13912 13484
rect 13964 13472 13970 13524
rect 14001 13515 14059 13521
rect 14001 13481 14013 13515
rect 14047 13512 14059 13515
rect 15654 13512 15660 13524
rect 14047 13484 15660 13512
rect 14047 13481 14059 13484
rect 14001 13475 14059 13481
rect 15654 13472 15660 13484
rect 15712 13472 15718 13524
rect 16758 13472 16764 13524
rect 16816 13512 16822 13524
rect 17497 13515 17555 13521
rect 17497 13512 17509 13515
rect 16816 13484 17509 13512
rect 16816 13472 16822 13484
rect 17497 13481 17509 13484
rect 17543 13481 17555 13515
rect 17497 13475 17555 13481
rect 18046 13472 18052 13524
rect 18104 13512 18110 13524
rect 18414 13512 18420 13524
rect 18104 13484 18420 13512
rect 18104 13472 18110 13484
rect 18414 13472 18420 13484
rect 18472 13472 18478 13524
rect 19058 13472 19064 13524
rect 19116 13472 19122 13524
rect 20530 13472 20536 13524
rect 20588 13512 20594 13524
rect 20625 13515 20683 13521
rect 20625 13512 20637 13515
rect 20588 13484 20637 13512
rect 20588 13472 20594 13484
rect 20625 13481 20637 13484
rect 20671 13481 20683 13515
rect 20625 13475 20683 13481
rect 21542 13472 21548 13524
rect 21600 13512 21606 13524
rect 21729 13515 21787 13521
rect 21729 13512 21741 13515
rect 21600 13484 21741 13512
rect 21600 13472 21606 13484
rect 21729 13481 21741 13484
rect 21775 13481 21787 13515
rect 21729 13475 21787 13481
rect 22002 13472 22008 13524
rect 22060 13512 22066 13524
rect 22060 13484 22140 13512
rect 22060 13472 22066 13484
rect 12250 13453 12256 13456
rect 9784 13416 10824 13444
rect 11072 13416 11183 13444
rect 11241 13447 11299 13453
rect 9784 13385 9812 13416
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13345 9551 13379
rect 9493 13339 9551 13345
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 9953 13379 10011 13385
rect 9953 13345 9965 13379
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 9125 13329 9183 13335
rect 9306 13268 9312 13320
rect 9364 13268 9370 13320
rect 9968 13308 9996 13339
rect 10042 13336 10048 13388
rect 10100 13336 10106 13388
rect 10321 13379 10379 13385
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 10502 13376 10508 13388
rect 10367 13348 10508 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 10502 13336 10508 13348
rect 10560 13382 10566 13388
rect 10597 13382 10655 13385
rect 10560 13379 10655 13382
rect 10560 13354 10609 13379
rect 10560 13336 10566 13354
rect 10597 13345 10609 13354
rect 10643 13345 10655 13379
rect 11072 13376 11100 13416
rect 11241 13413 11253 13447
rect 11287 13444 11299 13447
rect 12244 13444 12256 13453
rect 11287 13416 11744 13444
rect 12211 13416 12256 13444
rect 11287 13413 11299 13416
rect 11241 13407 11299 13413
rect 10597 13339 10655 13345
rect 10704 13348 11100 13376
rect 11149 13379 11207 13385
rect 10704 13308 10732 13348
rect 11149 13345 11161 13379
rect 11195 13376 11207 13379
rect 11606 13376 11612 13388
rect 11195 13348 11612 13376
rect 11195 13345 11207 13348
rect 11149 13339 11207 13345
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 11716 13385 11744 13416
rect 12244 13407 12256 13416
rect 12250 13404 12256 13407
rect 12308 13404 12314 13456
rect 15933 13447 15991 13453
rect 15933 13444 15945 13447
rect 12728 13416 15945 13444
rect 12728 13388 12756 13416
rect 15933 13413 15945 13416
rect 15979 13444 15991 13447
rect 17586 13444 17592 13456
rect 15979 13416 17592 13444
rect 15979 13413 15991 13416
rect 15933 13407 15991 13413
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 19512 13447 19570 13453
rect 17788 13416 19288 13444
rect 17788 13388 17816 13416
rect 11701 13379 11759 13385
rect 11701 13345 11713 13379
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 12710 13336 12716 13388
rect 12768 13336 12774 13388
rect 13814 13336 13820 13388
rect 13872 13336 13878 13388
rect 13909 13379 13967 13385
rect 13909 13345 13921 13379
rect 13955 13345 13967 13379
rect 13909 13339 13967 13345
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 9968 13280 10732 13308
rect 11624 13280 11989 13308
rect 10689 13243 10747 13249
rect 8864 13212 9996 13240
rect 8076 13200 8082 13212
rect 7374 13132 7380 13184
rect 7432 13132 7438 13184
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 7929 13175 7987 13181
rect 7929 13172 7941 13175
rect 7800 13144 7941 13172
rect 7800 13132 7806 13144
rect 7929 13141 7941 13144
rect 7975 13141 7987 13175
rect 7929 13135 7987 13141
rect 8110 13132 8116 13184
rect 8168 13172 8174 13184
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 8168 13144 8493 13172
rect 8168 13132 8174 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8481 13135 8539 13141
rect 8757 13175 8815 13181
rect 8757 13141 8769 13175
rect 8803 13172 8815 13175
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8803 13144 9045 13172
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 9033 13141 9045 13144
rect 9079 13141 9091 13175
rect 9033 13135 9091 13141
rect 9858 13132 9864 13184
rect 9916 13132 9922 13184
rect 9968 13172 9996 13212
rect 10689 13209 10701 13243
rect 10735 13240 10747 13243
rect 11238 13240 11244 13252
rect 10735 13212 11244 13240
rect 10735 13209 10747 13212
rect 10689 13203 10747 13209
rect 11238 13200 11244 13212
rect 11296 13200 11302 13252
rect 11624 13184 11652 13280
rect 11977 13277 11989 13280
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 13924 13252 13952 13339
rect 16206 13336 16212 13388
rect 16264 13376 16270 13388
rect 16373 13379 16431 13385
rect 16373 13376 16385 13379
rect 16264 13348 16385 13376
rect 16264 13336 16270 13348
rect 16373 13345 16385 13348
rect 16419 13345 16431 13379
rect 16373 13339 16431 13345
rect 17681 13379 17739 13385
rect 17681 13345 17693 13379
rect 17727 13376 17739 13379
rect 17770 13376 17776 13388
rect 17727 13348 17776 13376
rect 17727 13345 17739 13348
rect 17681 13339 17739 13345
rect 17770 13336 17776 13348
rect 17828 13336 17834 13388
rect 17954 13385 17960 13388
rect 17948 13376 17960 13385
rect 17915 13348 17960 13376
rect 17948 13339 17960 13348
rect 17954 13336 17960 13339
rect 18012 13336 18018 13388
rect 19260 13385 19288 13416
rect 19512 13413 19524 13447
rect 19558 13444 19570 13447
rect 20346 13444 20352 13456
rect 19558 13416 20352 13444
rect 19558 13413 19570 13416
rect 19512 13407 19570 13413
rect 20346 13404 20352 13416
rect 20404 13404 20410 13456
rect 19245 13379 19303 13385
rect 19245 13345 19257 13379
rect 19291 13345 19303 13379
rect 19245 13339 19303 13345
rect 20993 13379 21051 13385
rect 20993 13345 21005 13379
rect 21039 13345 21051 13379
rect 20993 13339 21051 13345
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 14185 13311 14243 13317
rect 14185 13308 14197 13311
rect 14056 13280 14197 13308
rect 14056 13268 14062 13280
rect 14185 13277 14197 13280
rect 14231 13308 14243 13311
rect 14642 13308 14648 13320
rect 14231 13280 14648 13308
rect 14231 13277 14243 13280
rect 14185 13271 14243 13277
rect 14642 13268 14648 13280
rect 14700 13308 14706 13320
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 14700 13280 16129 13308
rect 14700 13268 14706 13280
rect 16117 13277 16129 13280
rect 16163 13277 16175 13311
rect 21008 13308 21036 13339
rect 21450 13336 21456 13388
rect 21508 13376 21514 13388
rect 21545 13379 21603 13385
rect 21545 13376 21557 13379
rect 21508 13348 21557 13376
rect 21508 13336 21514 13348
rect 21545 13345 21557 13348
rect 21591 13345 21603 13379
rect 21545 13339 21603 13345
rect 21637 13379 21695 13385
rect 21637 13345 21649 13379
rect 21683 13376 21695 13379
rect 21726 13376 21732 13388
rect 21683 13348 21732 13376
rect 21683 13345 21695 13348
rect 21637 13339 21695 13345
rect 21082 13308 21088 13320
rect 21008 13280 21088 13308
rect 16117 13271 16175 13277
rect 21082 13268 21088 13280
rect 21140 13308 21146 13320
rect 21266 13308 21272 13320
rect 21140 13280 21272 13308
rect 21140 13268 21146 13280
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 21560 13308 21588 13339
rect 21726 13336 21732 13348
rect 21784 13336 21790 13388
rect 22112 13385 22140 13484
rect 23198 13472 23204 13524
rect 23256 13512 23262 13524
rect 23256 13484 24808 13512
rect 23256 13472 23262 13484
rect 22554 13444 22560 13456
rect 22204 13416 22560 13444
rect 22097 13379 22155 13385
rect 22097 13345 22109 13379
rect 22143 13345 22155 13379
rect 22097 13339 22155 13345
rect 22204 13320 22232 13416
rect 22554 13404 22560 13416
rect 22612 13444 22618 13456
rect 24210 13444 24216 13456
rect 22612 13416 23796 13444
rect 22612 13404 22618 13416
rect 22456 13379 22514 13385
rect 22456 13345 22468 13379
rect 22502 13376 22514 13379
rect 23658 13376 23664 13388
rect 22502 13348 23664 13376
rect 22502 13345 22514 13348
rect 22456 13339 22514 13345
rect 23658 13336 23664 13348
rect 23716 13336 23722 13388
rect 23768 13385 23796 13416
rect 23860 13416 24216 13444
rect 23753 13379 23811 13385
rect 23753 13345 23765 13379
rect 23799 13345 23811 13379
rect 23753 13339 23811 13345
rect 21818 13308 21824 13320
rect 21560 13280 21824 13308
rect 21818 13268 21824 13280
rect 21876 13268 21882 13320
rect 22186 13268 22192 13320
rect 22244 13268 22250 13320
rect 23860 13308 23888 13416
rect 24210 13404 24216 13416
rect 24268 13444 24274 13456
rect 24578 13444 24584 13456
rect 24268 13416 24584 13444
rect 24268 13404 24274 13416
rect 24578 13404 24584 13416
rect 24636 13444 24642 13456
rect 24780 13444 24808 13484
rect 25314 13472 25320 13524
rect 25372 13472 25378 13524
rect 25406 13472 25412 13524
rect 25464 13512 25470 13524
rect 25685 13515 25743 13521
rect 25685 13512 25697 13515
rect 25464 13484 25697 13512
rect 25464 13472 25470 13484
rect 25685 13481 25697 13484
rect 25731 13481 25743 13515
rect 25685 13475 25743 13481
rect 25958 13472 25964 13524
rect 26016 13472 26022 13524
rect 26418 13472 26424 13524
rect 26476 13512 26482 13524
rect 31662 13512 31668 13524
rect 26476 13484 31668 13512
rect 26476 13472 26482 13484
rect 31662 13472 31668 13484
rect 31720 13472 31726 13524
rect 24636 13416 24716 13444
rect 24780 13416 25360 13444
rect 24636 13404 24642 13416
rect 24020 13379 24078 13385
rect 24020 13345 24032 13379
rect 24066 13376 24078 13379
rect 24486 13376 24492 13388
rect 24066 13348 24492 13376
rect 24066 13345 24078 13348
rect 24020 13339 24078 13345
rect 24486 13336 24492 13348
rect 24544 13336 24550 13388
rect 24688 13376 24716 13416
rect 24854 13376 24860 13388
rect 24688 13348 24860 13376
rect 24826 13336 24860 13348
rect 24912 13336 24918 13388
rect 25332 13385 25360 13416
rect 25774 13404 25780 13456
rect 25832 13444 25838 13456
rect 25832 13416 26464 13444
rect 25832 13404 25838 13416
rect 25317 13379 25375 13385
rect 25317 13345 25329 13379
rect 25363 13345 25375 13379
rect 25317 13339 25375 13345
rect 25498 13336 25504 13388
rect 25556 13336 25562 13388
rect 25593 13379 25651 13385
rect 25593 13345 25605 13379
rect 25639 13345 25651 13379
rect 25593 13339 25651 13345
rect 23492 13280 23888 13308
rect 24826 13308 24854 13336
rect 25608 13308 25636 13339
rect 25682 13336 25688 13388
rect 25740 13376 25746 13388
rect 26436 13385 26464 13416
rect 25869 13379 25927 13385
rect 25869 13376 25881 13379
rect 25740 13348 25881 13376
rect 25740 13336 25746 13348
rect 25869 13345 25881 13348
rect 25915 13345 25927 13379
rect 25869 13339 25927 13345
rect 26421 13379 26479 13385
rect 26421 13345 26433 13379
rect 26467 13345 26479 13379
rect 26421 13339 26479 13345
rect 24826 13280 25636 13308
rect 25884 13308 25912 13339
rect 25958 13308 25964 13320
rect 25884 13280 25964 13308
rect 13906 13200 13912 13252
rect 13964 13240 13970 13252
rect 21910 13240 21916 13252
rect 13964 13212 15792 13240
rect 13964 13200 13970 13212
rect 11330 13172 11336 13184
rect 9968 13144 11336 13172
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 11514 13132 11520 13184
rect 11572 13132 11578 13184
rect 11606 13132 11612 13184
rect 11664 13132 11670 13184
rect 11793 13175 11851 13181
rect 11793 13141 11805 13175
rect 11839 13172 11851 13175
rect 12986 13172 12992 13184
rect 11839 13144 12992 13172
rect 11839 13141 11851 13144
rect 11793 13135 11851 13141
rect 12986 13132 12992 13144
rect 13044 13132 13050 13184
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 15470 13172 15476 13184
rect 14332 13144 15476 13172
rect 14332 13132 14338 13144
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 15764 13172 15792 13212
rect 20732 13212 21916 13240
rect 20732 13184 20760 13212
rect 21910 13200 21916 13212
rect 21968 13240 21974 13252
rect 22005 13243 22063 13249
rect 22005 13240 22017 13243
rect 21968 13212 22017 13240
rect 21968 13200 21974 13212
rect 22005 13209 22017 13212
rect 22051 13209 22063 13243
rect 22005 13203 22063 13209
rect 16850 13172 16856 13184
rect 15764 13144 16856 13172
rect 16850 13132 16856 13144
rect 16908 13132 16914 13184
rect 20714 13132 20720 13184
rect 20772 13132 20778 13184
rect 20898 13132 20904 13184
rect 20956 13132 20962 13184
rect 21450 13132 21456 13184
rect 21508 13132 21514 13184
rect 22020 13172 22048 13203
rect 23492 13172 23520 13280
rect 25958 13268 25964 13280
rect 26016 13268 26022 13320
rect 24826 13212 28304 13240
rect 22020 13144 23520 13172
rect 23569 13175 23627 13181
rect 23569 13141 23581 13175
rect 23615 13172 23627 13175
rect 24826 13172 24854 13212
rect 28276 13184 28304 13212
rect 23615 13144 24854 13172
rect 25133 13175 25191 13181
rect 23615 13141 23627 13144
rect 23569 13135 23627 13141
rect 25133 13141 25145 13175
rect 25179 13172 25191 13175
rect 26418 13172 26424 13184
rect 25179 13144 26424 13172
rect 25179 13141 25191 13144
rect 25133 13135 25191 13141
rect 26418 13132 26424 13144
rect 26476 13132 26482 13184
rect 26510 13132 26516 13184
rect 26568 13132 26574 13184
rect 28258 13132 28264 13184
rect 28316 13132 28322 13184
rect 552 13082 31372 13104
rect 552 13030 4250 13082
rect 4302 13030 4314 13082
rect 4366 13030 4378 13082
rect 4430 13030 4442 13082
rect 4494 13030 4506 13082
rect 4558 13030 11955 13082
rect 12007 13030 12019 13082
rect 12071 13030 12083 13082
rect 12135 13030 12147 13082
rect 12199 13030 12211 13082
rect 12263 13030 19660 13082
rect 19712 13030 19724 13082
rect 19776 13030 19788 13082
rect 19840 13030 19852 13082
rect 19904 13030 19916 13082
rect 19968 13030 27365 13082
rect 27417 13030 27429 13082
rect 27481 13030 27493 13082
rect 27545 13030 27557 13082
rect 27609 13030 27621 13082
rect 27673 13030 31372 13082
rect 552 13008 31372 13030
rect 7558 12928 7564 12980
rect 7616 12928 7622 12980
rect 7742 12928 7748 12980
rect 7800 12928 7806 12980
rect 8938 12928 8944 12980
rect 8996 12928 9002 12980
rect 9398 12928 9404 12980
rect 9456 12928 9462 12980
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 10962 12968 10968 12980
rect 10827 12940 10968 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 12989 12971 13047 12977
rect 12989 12937 13001 12971
rect 13035 12968 13047 12971
rect 13446 12968 13452 12980
rect 13035 12940 13452 12968
rect 13035 12937 13047 12940
rect 12989 12931 13047 12937
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 15013 12971 15071 12977
rect 15013 12937 15025 12971
rect 15059 12968 15071 12971
rect 15378 12968 15384 12980
rect 15059 12940 15384 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 16850 12928 16856 12980
rect 16908 12968 16914 12980
rect 17678 12968 17684 12980
rect 16908 12940 17684 12968
rect 16908 12928 16914 12940
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 18138 12928 18144 12980
rect 18196 12968 18202 12980
rect 18417 12971 18475 12977
rect 18417 12968 18429 12971
rect 18196 12940 18429 12968
rect 18196 12928 18202 12940
rect 18417 12937 18429 12940
rect 18463 12937 18475 12971
rect 18417 12931 18475 12937
rect 20073 12971 20131 12977
rect 20073 12937 20085 12971
rect 20119 12968 20131 12971
rect 20162 12968 20168 12980
rect 20119 12940 20168 12968
rect 20119 12937 20131 12940
rect 20073 12931 20131 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 24486 12928 24492 12980
rect 24544 12928 24550 12980
rect 24670 12928 24676 12980
rect 24728 12968 24734 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 24728 12940 24777 12968
rect 24728 12928 24734 12940
rect 24765 12937 24777 12940
rect 24811 12937 24823 12971
rect 24765 12931 24823 12937
rect 25866 12928 25872 12980
rect 25924 12928 25930 12980
rect 7760 12832 7788 12928
rect 7883 12903 7941 12909
rect 7883 12869 7895 12903
rect 7929 12900 7941 12903
rect 9030 12900 9036 12912
rect 7929 12872 9036 12900
rect 7929 12869 7941 12872
rect 7883 12863 7941 12869
rect 9030 12860 9036 12872
rect 9088 12860 9094 12912
rect 9416 12900 9444 12928
rect 9140 12872 9444 12900
rect 10505 12903 10563 12909
rect 8846 12832 8852 12844
rect 7668 12804 7788 12832
rect 7852 12804 8852 12832
rect 7668 12773 7696 12804
rect 7653 12767 7711 12773
rect 7852 12767 7880 12804
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 7653 12733 7665 12767
rect 7699 12733 7711 12767
rect 7653 12727 7711 12733
rect 7812 12761 7880 12767
rect 7812 12727 7824 12761
rect 7858 12730 7880 12761
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 8110 12764 8116 12776
rect 8067 12736 8116 12764
rect 8067 12733 8079 12736
rect 7858 12727 7870 12730
rect 8021 12727 8079 12733
rect 7812 12721 7870 12727
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8205 12767 8263 12773
rect 8205 12733 8217 12767
rect 8251 12733 8263 12767
rect 8205 12727 8263 12733
rect 8220 12696 8248 12727
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 8444 12736 8585 12764
rect 8444 12724 8450 12736
rect 8573 12733 8585 12736
rect 8619 12764 8631 12767
rect 9140 12764 9168 12872
rect 10505 12869 10517 12903
rect 10551 12900 10563 12903
rect 11054 12900 11060 12912
rect 10551 12872 11060 12900
rect 10551 12869 10563 12872
rect 10505 12863 10563 12869
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 13630 12900 13636 12912
rect 12676 12872 13636 12900
rect 12676 12860 12682 12872
rect 13630 12860 13636 12872
rect 13688 12860 13694 12912
rect 15286 12860 15292 12912
rect 15344 12900 15350 12912
rect 16485 12903 16543 12909
rect 16485 12900 16497 12903
rect 15344 12872 16497 12900
rect 15344 12860 15350 12872
rect 16485 12869 16497 12872
rect 16531 12869 16543 12903
rect 16485 12863 16543 12869
rect 21358 12860 21364 12912
rect 21416 12900 21422 12912
rect 21416 12872 24808 12900
rect 21416 12860 21422 12872
rect 10594 12832 10600 12844
rect 10428 12804 10600 12832
rect 10428 12776 10456 12804
rect 10594 12792 10600 12804
rect 10652 12792 10658 12844
rect 21082 12792 21088 12844
rect 21140 12832 21146 12844
rect 21140 12804 21956 12832
rect 21140 12792 21146 12804
rect 21376 12776 21404 12804
rect 8619 12736 9168 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 9766 12724 9772 12776
rect 9824 12764 9830 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 9824 12736 10333 12764
rect 9824 12724 9830 12736
rect 8754 12696 8760 12708
rect 8220 12668 8760 12696
rect 8754 12656 8760 12668
rect 8812 12656 8818 12708
rect 9122 12656 9128 12708
rect 9180 12696 9186 12708
rect 10054 12699 10112 12705
rect 10054 12696 10066 12699
rect 9180 12668 10066 12696
rect 9180 12656 9186 12668
rect 10054 12665 10066 12668
rect 10100 12665 10112 12699
rect 10054 12659 10112 12665
rect 10152 12696 10180 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 10410 12724 10416 12776
rect 10468 12724 10474 12776
rect 10873 12767 10931 12773
rect 10873 12733 10885 12767
rect 10919 12764 10931 12767
rect 11238 12764 11244 12776
rect 10919 12736 11244 12764
rect 10919 12733 10931 12736
rect 10873 12727 10931 12733
rect 11238 12724 11244 12736
rect 11296 12764 11302 12776
rect 11296 12736 12434 12764
rect 11296 12724 11302 12736
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 10152 12668 10977 12696
rect 10152 12640 10180 12668
rect 10965 12665 10977 12668
rect 11011 12696 11023 12699
rect 11146 12696 11152 12708
rect 11011 12668 11152 12696
rect 11011 12665 11023 12668
rect 10965 12659 11023 12665
rect 11146 12656 11152 12668
rect 11204 12696 11210 12708
rect 11606 12696 11612 12708
rect 11204 12668 11612 12696
rect 11204 12656 11210 12668
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 8205 12631 8263 12637
rect 8205 12597 8217 12631
rect 8251 12628 8263 12631
rect 8478 12628 8484 12640
rect 8251 12600 8484 12628
rect 8251 12597 8263 12600
rect 8205 12591 8263 12597
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 8665 12631 8723 12637
rect 8665 12597 8677 12631
rect 8711 12628 8723 12631
rect 9398 12628 9404 12640
rect 8711 12600 9404 12628
rect 8711 12597 8723 12600
rect 8665 12591 8723 12597
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 10134 12588 10140 12640
rect 10192 12588 10198 12640
rect 12406 12628 12434 12736
rect 12710 12724 12716 12776
rect 12768 12724 12774 12776
rect 12894 12724 12900 12776
rect 12952 12724 12958 12776
rect 13170 12724 13176 12776
rect 13228 12724 13234 12776
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 13679 12736 14044 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 14016 12708 14044 12736
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 16942 12764 16948 12776
rect 15252 12736 16948 12764
rect 15252 12724 15258 12736
rect 16942 12724 16948 12736
rect 17000 12724 17006 12776
rect 17034 12724 17040 12776
rect 17092 12764 17098 12776
rect 17770 12764 17776 12776
rect 17092 12736 17776 12764
rect 17092 12724 17098 12736
rect 17770 12724 17776 12736
rect 17828 12764 17834 12776
rect 18693 12767 18751 12773
rect 18693 12764 18705 12767
rect 17828 12736 18705 12764
rect 17828 12724 17834 12736
rect 18693 12733 18705 12736
rect 18739 12733 18751 12767
rect 18693 12727 18751 12733
rect 20441 12767 20499 12773
rect 20441 12733 20453 12767
rect 20487 12764 20499 12767
rect 20625 12767 20683 12773
rect 20625 12764 20637 12767
rect 20487 12736 20637 12764
rect 20487 12733 20499 12736
rect 20441 12727 20499 12733
rect 20625 12733 20637 12736
rect 20671 12733 20683 12767
rect 20625 12727 20683 12733
rect 20714 12724 20720 12776
rect 20772 12724 20778 12776
rect 20990 12724 20996 12776
rect 21048 12724 21054 12776
rect 21269 12767 21327 12773
rect 21269 12733 21281 12767
rect 21315 12733 21327 12767
rect 21269 12727 21327 12733
rect 12986 12656 12992 12708
rect 13044 12696 13050 12708
rect 13878 12699 13936 12705
rect 13878 12696 13890 12699
rect 13044 12668 13890 12696
rect 13044 12656 13050 12668
rect 13878 12665 13890 12668
rect 13924 12665 13936 12699
rect 13878 12659 13936 12665
rect 13998 12656 14004 12708
rect 14056 12656 14062 12708
rect 17126 12656 17132 12708
rect 17184 12696 17190 12708
rect 17282 12699 17340 12705
rect 17282 12696 17294 12699
rect 17184 12668 17294 12696
rect 17184 12656 17190 12668
rect 17282 12665 17294 12668
rect 17328 12665 17340 12699
rect 17282 12659 17340 12665
rect 18960 12699 19018 12705
rect 18960 12665 18972 12699
rect 19006 12696 19018 12699
rect 20349 12699 20407 12705
rect 20349 12696 20361 12699
rect 19006 12668 20361 12696
rect 19006 12665 19018 12668
rect 18960 12659 19018 12665
rect 20349 12665 20361 12668
rect 20395 12665 20407 12699
rect 20349 12659 20407 12665
rect 20806 12656 20812 12708
rect 20864 12696 20870 12708
rect 21284 12696 21312 12727
rect 21358 12724 21364 12776
rect 21416 12724 21422 12776
rect 21542 12724 21548 12776
rect 21600 12724 21606 12776
rect 21818 12724 21824 12776
rect 21876 12724 21882 12776
rect 21928 12764 21956 12804
rect 22646 12792 22652 12844
rect 22704 12832 22710 12844
rect 24213 12835 24271 12841
rect 22704 12804 24164 12832
rect 22704 12792 22710 12804
rect 21928 12736 23704 12764
rect 23676 12705 23704 12736
rect 23842 12724 23848 12776
rect 23900 12724 23906 12776
rect 23934 12724 23940 12776
rect 23992 12724 23998 12776
rect 24026 12724 24032 12776
rect 24084 12724 24090 12776
rect 24136 12773 24164 12804
rect 24213 12801 24225 12835
rect 24259 12832 24271 12835
rect 24259 12804 24624 12832
rect 24259 12801 24271 12804
rect 24213 12795 24271 12801
rect 24121 12767 24179 12773
rect 24121 12733 24133 12767
rect 24167 12733 24179 12767
rect 24121 12727 24179 12733
rect 24302 12724 24308 12776
rect 24360 12724 24366 12776
rect 24397 12767 24455 12773
rect 24397 12733 24409 12767
rect 24443 12733 24455 12767
rect 24397 12727 24455 12733
rect 21729 12699 21787 12705
rect 21729 12696 21741 12699
rect 20864 12668 21220 12696
rect 21284 12668 21741 12696
rect 20864 12656 20870 12668
rect 12618 12628 12624 12640
rect 12406 12600 12624 12628
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 13262 12588 13268 12640
rect 13320 12588 13326 12640
rect 20901 12631 20959 12637
rect 20901 12597 20913 12631
rect 20947 12628 20959 12631
rect 21082 12628 21088 12640
rect 20947 12600 21088 12628
rect 20947 12597 20959 12600
rect 20901 12591 20959 12597
rect 21082 12588 21088 12600
rect 21140 12588 21146 12640
rect 21192 12637 21220 12668
rect 21729 12665 21741 12668
rect 21775 12665 21787 12699
rect 21729 12659 21787 12665
rect 21913 12699 21971 12705
rect 21913 12665 21925 12699
rect 21959 12665 21971 12699
rect 21913 12659 21971 12665
rect 23661 12699 23719 12705
rect 23661 12665 23673 12699
rect 23707 12665 23719 12699
rect 24044 12696 24072 12724
rect 24412 12696 24440 12727
rect 24044 12668 24440 12696
rect 24596 12696 24624 12804
rect 24673 12767 24731 12773
rect 24673 12733 24685 12767
rect 24719 12764 24731 12767
rect 24780 12764 24808 12872
rect 24854 12860 24860 12912
rect 24912 12860 24918 12912
rect 25884 12900 25912 12928
rect 25424 12872 25912 12900
rect 26160 12872 26648 12900
rect 24872 12773 24900 12860
rect 24719 12736 24808 12764
rect 24857 12767 24915 12773
rect 24719 12733 24731 12736
rect 24673 12727 24731 12733
rect 24857 12733 24869 12767
rect 24903 12733 24915 12767
rect 24857 12727 24915 12733
rect 24946 12724 24952 12776
rect 25004 12724 25010 12776
rect 25424 12773 25452 12872
rect 25590 12792 25596 12844
rect 25648 12792 25654 12844
rect 25774 12792 25780 12844
rect 25832 12832 25838 12844
rect 26160 12841 26188 12872
rect 26145 12835 26203 12841
rect 26145 12832 26157 12835
rect 25832 12804 26157 12832
rect 25832 12792 25838 12804
rect 25976 12773 26004 12804
rect 26145 12801 26157 12804
rect 26191 12801 26203 12835
rect 26421 12835 26479 12841
rect 26421 12832 26433 12835
rect 26145 12795 26203 12801
rect 26252 12804 26433 12832
rect 26252 12773 26280 12804
rect 26421 12801 26433 12804
rect 26467 12801 26479 12835
rect 26421 12795 26479 12801
rect 25409 12767 25467 12773
rect 25409 12733 25421 12767
rect 25455 12733 25467 12767
rect 25409 12727 25467 12733
rect 25685 12767 25743 12773
rect 25685 12733 25697 12767
rect 25731 12764 25743 12767
rect 25869 12767 25927 12773
rect 25869 12764 25881 12767
rect 25731 12736 25881 12764
rect 25731 12733 25743 12736
rect 25685 12727 25743 12733
rect 25869 12733 25881 12736
rect 25915 12733 25927 12767
rect 25869 12727 25927 12733
rect 25961 12767 26019 12773
rect 25961 12733 25973 12767
rect 26007 12733 26019 12767
rect 25961 12727 26019 12733
rect 26237 12767 26295 12773
rect 26237 12733 26249 12767
rect 26283 12733 26295 12767
rect 26237 12727 26295 12733
rect 26326 12724 26332 12776
rect 26384 12724 26390 12776
rect 26620 12773 26648 12872
rect 26605 12767 26663 12773
rect 26605 12733 26617 12767
rect 26651 12733 26663 12767
rect 26605 12727 26663 12733
rect 25317 12699 25375 12705
rect 25317 12696 25329 12699
rect 24596 12668 25329 12696
rect 23661 12659 23719 12665
rect 25317 12665 25329 12668
rect 25363 12665 25375 12699
rect 25317 12659 25375 12665
rect 21177 12631 21235 12637
rect 21177 12597 21189 12631
rect 21223 12597 21235 12631
rect 21177 12591 21235 12597
rect 21453 12631 21511 12637
rect 21453 12597 21465 12631
rect 21499 12628 21511 12631
rect 21634 12628 21640 12640
rect 21499 12600 21640 12628
rect 21499 12597 21511 12600
rect 21453 12591 21511 12597
rect 21634 12588 21640 12600
rect 21692 12588 21698 12640
rect 21928 12628 21956 12659
rect 22370 12628 22376 12640
rect 21928 12600 22376 12628
rect 22370 12588 22376 12600
rect 22428 12588 22434 12640
rect 23676 12628 23704 12659
rect 26050 12656 26056 12708
rect 26108 12696 26114 12708
rect 26697 12699 26755 12705
rect 26697 12696 26709 12699
rect 26108 12668 26709 12696
rect 26108 12656 26114 12668
rect 26697 12665 26709 12668
rect 26743 12665 26755 12699
rect 26697 12659 26755 12665
rect 24302 12628 24308 12640
rect 23676 12600 24308 12628
rect 24302 12588 24308 12600
rect 24360 12588 24366 12640
rect 24394 12588 24400 12640
rect 24452 12628 24458 12640
rect 25041 12631 25099 12637
rect 25041 12628 25053 12631
rect 24452 12600 25053 12628
rect 24452 12588 24458 12600
rect 25041 12597 25053 12600
rect 25087 12597 25099 12631
rect 25041 12591 25099 12597
rect 552 12538 31531 12560
rect 552 12486 8102 12538
rect 8154 12486 8166 12538
rect 8218 12486 8230 12538
rect 8282 12486 8294 12538
rect 8346 12486 8358 12538
rect 8410 12486 15807 12538
rect 15859 12486 15871 12538
rect 15923 12486 15935 12538
rect 15987 12486 15999 12538
rect 16051 12486 16063 12538
rect 16115 12486 23512 12538
rect 23564 12486 23576 12538
rect 23628 12486 23640 12538
rect 23692 12486 23704 12538
rect 23756 12486 23768 12538
rect 23820 12486 31217 12538
rect 31269 12486 31281 12538
rect 31333 12486 31345 12538
rect 31397 12486 31409 12538
rect 31461 12486 31473 12538
rect 31525 12486 31531 12538
rect 552 12464 31531 12486
rect 8478 12384 8484 12436
rect 8536 12384 8542 12436
rect 8570 12384 8576 12436
rect 8628 12384 8634 12436
rect 8754 12384 8760 12436
rect 8812 12384 8818 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9263 12427 9321 12433
rect 9263 12424 9275 12427
rect 8904 12396 9275 12424
rect 8904 12384 8910 12396
rect 9263 12393 9275 12396
rect 9309 12393 9321 12427
rect 9263 12387 9321 12393
rect 9398 12384 9404 12436
rect 9456 12384 9462 12436
rect 9585 12427 9643 12433
rect 9585 12393 9597 12427
rect 9631 12424 9643 12427
rect 9858 12424 9864 12436
rect 9631 12396 9864 12424
rect 9631 12393 9643 12396
rect 9585 12387 9643 12393
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10042 12384 10048 12436
rect 10100 12384 10106 12436
rect 10226 12384 10232 12436
rect 10284 12384 10290 12436
rect 11149 12427 11207 12433
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 11238 12424 11244 12436
rect 11195 12396 11244 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 11422 12384 11428 12436
rect 11480 12384 11486 12436
rect 11974 12384 11980 12436
rect 12032 12384 12038 12436
rect 12529 12427 12587 12433
rect 12529 12393 12541 12427
rect 12575 12424 12587 12427
rect 12710 12424 12716 12436
rect 12575 12396 12716 12424
rect 12575 12393 12587 12396
rect 12529 12387 12587 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12424 12863 12427
rect 12851 12396 12940 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 8205 12359 8263 12365
rect 8205 12325 8217 12359
rect 8251 12356 8263 12359
rect 8588 12356 8616 12384
rect 9416 12356 9444 12384
rect 10060 12356 10088 12384
rect 10778 12356 10784 12368
rect 8251 12328 8616 12356
rect 8772 12328 9168 12356
rect 9416 12328 9812 12356
rect 8251 12325 8263 12328
rect 8205 12319 8263 12325
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 7837 12291 7895 12297
rect 7837 12288 7849 12291
rect 7432 12260 7849 12288
rect 7432 12248 7438 12260
rect 7837 12257 7849 12260
rect 7883 12257 7895 12291
rect 7837 12251 7895 12257
rect 8110 12248 8116 12300
rect 8168 12248 8174 12300
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12288 8631 12291
rect 8772 12288 8800 12328
rect 9140 12297 9168 12328
rect 8619 12260 8800 12288
rect 8849 12291 8907 12297
rect 8619 12257 8631 12260
rect 8573 12251 8631 12257
rect 8849 12257 8861 12291
rect 8895 12257 8907 12291
rect 8849 12251 8907 12257
rect 9125 12291 9183 12297
rect 9125 12257 9137 12291
rect 9171 12288 9183 12291
rect 9214 12288 9220 12300
rect 9171 12260 9220 12288
rect 9171 12257 9183 12260
rect 9125 12251 9183 12257
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 8864 12220 8892 12251
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 9398 12297 9404 12300
rect 9366 12291 9404 12297
rect 9366 12257 9378 12291
rect 9366 12251 9404 12257
rect 9398 12248 9404 12251
rect 9456 12248 9462 12300
rect 9784 12297 9812 12328
rect 9876 12328 10088 12356
rect 10244 12328 10784 12356
rect 9876 12297 9904 12328
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12257 9827 12291
rect 9769 12251 9827 12257
rect 9861 12291 9919 12297
rect 9861 12257 9873 12291
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 8720 12192 8892 12220
rect 9692 12220 9720 12251
rect 10042 12248 10048 12300
rect 10100 12248 10106 12300
rect 10244 12297 10272 12328
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 12912 12356 12940 12396
rect 12986 12384 12992 12436
rect 13044 12424 13050 12436
rect 13170 12424 13176 12436
rect 13044 12396 13176 12424
rect 13044 12384 13050 12396
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 13354 12384 13360 12436
rect 13412 12424 13418 12436
rect 15013 12427 15071 12433
rect 13412 12396 14412 12424
rect 13412 12384 13418 12396
rect 14182 12356 14188 12368
rect 12360 12328 12848 12356
rect 12912 12328 13400 12356
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12257 10287 12291
rect 10229 12251 10287 12257
rect 10318 12248 10324 12300
rect 10376 12248 10382 12300
rect 10413 12291 10471 12297
rect 10413 12257 10425 12291
rect 10459 12288 10471 12291
rect 10597 12291 10655 12297
rect 10597 12288 10609 12291
rect 10459 12260 10609 12288
rect 10459 12257 10471 12260
rect 10413 12251 10471 12257
rect 10597 12257 10609 12260
rect 10643 12257 10655 12291
rect 10597 12251 10655 12257
rect 11054 12248 11060 12300
rect 11112 12248 11118 12300
rect 11514 12248 11520 12300
rect 11572 12248 11578 12300
rect 11606 12248 11612 12300
rect 11664 12248 11670 12300
rect 11885 12291 11943 12297
rect 11885 12257 11897 12291
rect 11931 12257 11943 12291
rect 11885 12251 11943 12257
rect 10336 12220 10364 12248
rect 9692 12192 10364 12220
rect 11900 12220 11928 12251
rect 12066 12248 12072 12300
rect 12124 12248 12130 12300
rect 12360 12297 12388 12328
rect 12345 12291 12403 12297
rect 12345 12257 12357 12291
rect 12391 12257 12403 12291
rect 12345 12251 12403 12257
rect 12434 12248 12440 12300
rect 12492 12288 12498 12300
rect 12705 12289 12763 12295
rect 12492 12286 12664 12288
rect 12705 12286 12717 12289
rect 12492 12260 12717 12286
rect 12492 12248 12498 12260
rect 12636 12258 12717 12260
rect 12705 12255 12717 12258
rect 12751 12255 12763 12289
rect 12820 12288 12848 12328
rect 12989 12291 13047 12297
rect 12989 12288 13001 12291
rect 12820 12260 13001 12288
rect 12705 12249 12763 12255
rect 12989 12257 13001 12260
rect 13035 12288 13047 12291
rect 13170 12288 13176 12300
rect 13035 12260 13176 12288
rect 13035 12257 13047 12260
rect 12989 12251 13047 12257
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 13262 12248 13268 12300
rect 13320 12248 13326 12300
rect 12802 12220 12808 12232
rect 11900 12192 12808 12220
rect 8720 12180 8726 12192
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 13372 12220 13400 12328
rect 13464 12328 14188 12356
rect 13464 12297 13492 12328
rect 14182 12316 14188 12328
rect 14240 12316 14246 12368
rect 14274 12316 14280 12368
rect 14332 12316 14338 12368
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 13541 12291 13599 12297
rect 13541 12257 13553 12291
rect 13587 12257 13599 12291
rect 13541 12251 13599 12257
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 13906 12288 13912 12300
rect 13679 12260 13912 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 13556 12220 13584 12251
rect 13906 12248 13912 12260
rect 13964 12288 13970 12300
rect 14001 12291 14059 12297
rect 14001 12288 14013 12291
rect 13964 12260 14013 12288
rect 13964 12248 13970 12260
rect 14001 12257 14013 12260
rect 14047 12288 14059 12291
rect 14090 12288 14096 12300
rect 14047 12260 14096 12288
rect 14047 12257 14059 12260
rect 14001 12251 14059 12257
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 14292 12287 14320 12316
rect 14384 12297 14412 12396
rect 15013 12393 15025 12427
rect 15059 12424 15071 12427
rect 15197 12427 15255 12433
rect 15197 12424 15209 12427
rect 15059 12396 15209 12424
rect 15059 12393 15071 12396
rect 15013 12387 15071 12393
rect 15197 12393 15209 12396
rect 15243 12393 15255 12427
rect 15197 12387 15255 12393
rect 15565 12427 15623 12433
rect 15565 12393 15577 12427
rect 15611 12424 15623 12427
rect 16761 12427 16819 12433
rect 16761 12424 16773 12427
rect 15611 12396 16773 12424
rect 15611 12393 15623 12396
rect 15565 12387 15623 12393
rect 16761 12393 16773 12396
rect 16807 12393 16819 12427
rect 16761 12387 16819 12393
rect 17770 12384 17776 12436
rect 17828 12424 17834 12436
rect 18877 12427 18935 12433
rect 18877 12424 18889 12427
rect 17828 12396 18889 12424
rect 17828 12384 17834 12396
rect 18877 12393 18889 12396
rect 18923 12393 18935 12427
rect 18877 12387 18935 12393
rect 20901 12427 20959 12433
rect 20901 12393 20913 12427
rect 20947 12424 20959 12427
rect 21634 12424 21640 12436
rect 20947 12396 21640 12424
rect 20947 12393 20959 12396
rect 20901 12387 20959 12393
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 21726 12384 21732 12436
rect 21784 12424 21790 12436
rect 24394 12424 24400 12436
rect 21784 12396 24400 12424
rect 21784 12384 21790 12396
rect 24394 12384 24400 12396
rect 24452 12384 24458 12436
rect 24489 12427 24547 12433
rect 24489 12393 24501 12427
rect 24535 12424 24547 12427
rect 28258 12424 28264 12436
rect 24535 12396 28264 12424
rect 24535 12393 24547 12396
rect 24489 12387 24547 12393
rect 28258 12384 28264 12396
rect 28316 12384 28322 12436
rect 15470 12316 15476 12368
rect 15528 12356 15534 12368
rect 18598 12356 18604 12368
rect 15528 12328 16252 12356
rect 15528 12316 15534 12328
rect 14369 12291 14427 12297
rect 14277 12281 14335 12287
rect 14277 12247 14289 12281
rect 14323 12247 14335 12281
rect 14369 12257 14381 12291
rect 14415 12257 14427 12291
rect 14369 12251 14427 12257
rect 14461 12291 14519 12297
rect 14461 12257 14473 12291
rect 14507 12288 14519 12291
rect 14645 12291 14703 12297
rect 14645 12288 14657 12291
rect 14507 12260 14657 12288
rect 14507 12257 14519 12260
rect 14461 12251 14519 12257
rect 14645 12257 14657 12260
rect 14691 12257 14703 12291
rect 14645 12251 14703 12257
rect 14277 12241 14335 12247
rect 13372 12192 13584 12220
rect 14384 12220 14412 12251
rect 14734 12248 14740 12300
rect 14792 12248 14798 12300
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 14752 12220 14780 12248
rect 14384 12192 14780 12220
rect 12253 12155 12311 12161
rect 12253 12121 12265 12155
rect 12299 12152 12311 12155
rect 12894 12152 12900 12164
rect 12299 12124 12900 12152
rect 12299 12121 12311 12124
rect 12253 12115 12311 12121
rect 12894 12112 12900 12124
rect 12952 12112 12958 12164
rect 13004 12124 13492 12152
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 8938 12084 8944 12096
rect 7975 12056 8944 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 8938 12044 8944 12056
rect 8996 12044 9002 12096
rect 9033 12087 9091 12093
rect 9033 12053 9045 12087
rect 9079 12084 9091 12087
rect 9214 12084 9220 12096
rect 9079 12056 9220 12084
rect 9079 12053 9091 12056
rect 9033 12047 9091 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 10686 12044 10692 12096
rect 10744 12044 10750 12096
rect 11701 12087 11759 12093
rect 11701 12053 11713 12087
rect 11747 12084 11759 12087
rect 13004 12084 13032 12124
rect 13464 12096 13492 12124
rect 13814 12112 13820 12164
rect 13872 12152 13878 12164
rect 14185 12155 14243 12161
rect 14185 12152 14197 12155
rect 13872 12124 14197 12152
rect 13872 12112 13878 12124
rect 14185 12121 14197 12124
rect 14231 12121 14243 12155
rect 14185 12115 14243 12121
rect 11747 12056 13032 12084
rect 13081 12087 13139 12093
rect 11747 12053 11759 12056
rect 11701 12047 11759 12053
rect 13081 12053 13093 12087
rect 13127 12084 13139 12087
rect 13357 12087 13415 12093
rect 13357 12084 13369 12087
rect 13127 12056 13369 12084
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 13357 12053 13369 12056
rect 13403 12053 13415 12087
rect 13357 12047 13415 12053
rect 13446 12044 13452 12096
rect 13504 12044 13510 12096
rect 13906 12044 13912 12096
rect 13964 12044 13970 12096
rect 14737 12087 14795 12093
rect 14737 12053 14749 12087
rect 14783 12084 14795 12087
rect 14936 12084 14964 12251
rect 15194 12248 15200 12300
rect 15252 12248 15258 12300
rect 15381 12291 15439 12297
rect 15381 12257 15393 12291
rect 15427 12257 15439 12291
rect 15381 12251 15439 12257
rect 15010 12180 15016 12232
rect 15068 12220 15074 12232
rect 15396 12220 15424 12251
rect 15654 12248 15660 12300
rect 15712 12248 15718 12300
rect 15746 12248 15752 12300
rect 15804 12248 15810 12300
rect 15838 12248 15844 12300
rect 15896 12248 15902 12300
rect 16117 12291 16175 12297
rect 16117 12257 16129 12291
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 15068 12192 15424 12220
rect 15068 12180 15074 12192
rect 15102 12112 15108 12164
rect 15160 12152 15166 12164
rect 16132 12152 16160 12251
rect 16224 12220 16252 12328
rect 16592 12328 18604 12356
rect 16592 12297 16620 12328
rect 17236 12297 17264 12328
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 21269 12359 21327 12365
rect 21269 12356 21281 12359
rect 18708 12328 21281 12356
rect 16577 12291 16635 12297
rect 16577 12257 16589 12291
rect 16623 12257 16635 12291
rect 16577 12251 16635 12257
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 17221 12291 17279 12297
rect 17221 12257 17233 12291
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 16684 12220 16712 12251
rect 16224 12192 16712 12220
rect 17144 12164 17172 12251
rect 17586 12248 17592 12300
rect 17644 12288 17650 12300
rect 18708 12288 18736 12328
rect 21269 12325 21281 12328
rect 21315 12325 21327 12359
rect 21269 12319 21327 12325
rect 23376 12359 23434 12365
rect 23376 12325 23388 12359
rect 23422 12356 23434 12359
rect 25869 12359 25927 12365
rect 25869 12356 25881 12359
rect 23422 12328 25881 12356
rect 23422 12325 23434 12328
rect 23376 12319 23434 12325
rect 25869 12325 25881 12328
rect 25915 12325 25927 12359
rect 25869 12319 25927 12325
rect 26050 12316 26056 12368
rect 26108 12316 26114 12368
rect 26142 12316 26148 12368
rect 26200 12316 26206 12368
rect 26510 12356 26516 12368
rect 26252 12328 26516 12356
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 17644 12260 18736 12288
rect 18800 12260 19441 12288
rect 17644 12248 17650 12260
rect 15160 12124 16160 12152
rect 15160 12112 15166 12124
rect 16298 12112 16304 12164
rect 16356 12152 16362 12164
rect 17037 12155 17095 12161
rect 17037 12152 17049 12155
rect 16356 12124 17049 12152
rect 16356 12112 16362 12124
rect 17037 12121 17049 12124
rect 17083 12121 17095 12155
rect 17037 12115 17095 12121
rect 17126 12112 17132 12164
rect 17184 12112 17190 12164
rect 18800 12152 18828 12260
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 19518 12248 19524 12300
rect 19576 12288 19582 12300
rect 19705 12291 19763 12297
rect 19705 12288 19717 12291
rect 19576 12260 19717 12288
rect 19576 12248 19582 12260
rect 19705 12257 19717 12260
rect 19751 12257 19763 12291
rect 19705 12251 19763 12257
rect 20165 12291 20223 12297
rect 20165 12257 20177 12291
rect 20211 12257 20223 12291
rect 20165 12251 20223 12257
rect 20180 12220 20208 12251
rect 20622 12248 20628 12300
rect 20680 12248 20686 12300
rect 20714 12248 20720 12300
rect 20772 12248 20778 12300
rect 20898 12248 20904 12300
rect 20956 12248 20962 12300
rect 21542 12248 21548 12300
rect 21600 12288 21606 12300
rect 24486 12288 24492 12300
rect 21600 12260 24492 12288
rect 21600 12248 21606 12260
rect 24486 12248 24492 12260
rect 24544 12248 24550 12300
rect 24578 12248 24584 12300
rect 24636 12288 24642 12300
rect 24673 12291 24731 12297
rect 24673 12288 24685 12291
rect 24636 12260 24685 12288
rect 24636 12248 24642 12260
rect 24673 12257 24685 12260
rect 24719 12257 24731 12291
rect 24673 12251 24731 12257
rect 24762 12248 24768 12300
rect 24820 12248 24826 12300
rect 25133 12291 25191 12297
rect 25133 12257 25145 12291
rect 25179 12288 25191 12291
rect 25317 12291 25375 12297
rect 25317 12288 25329 12291
rect 25179 12260 25329 12288
rect 25179 12257 25191 12260
rect 25133 12251 25191 12257
rect 25317 12257 25329 12260
rect 25363 12257 25375 12291
rect 25317 12251 25375 12257
rect 25409 12291 25467 12297
rect 25409 12257 25421 12291
rect 25455 12288 25467 12291
rect 25501 12291 25559 12297
rect 25501 12288 25513 12291
rect 25455 12260 25513 12288
rect 25455 12257 25467 12260
rect 25409 12251 25467 12257
rect 25501 12257 25513 12260
rect 25547 12257 25559 12291
rect 25501 12251 25559 12257
rect 25961 12291 26019 12297
rect 25961 12257 25973 12291
rect 26007 12288 26019 12291
rect 26068 12288 26096 12316
rect 26252 12297 26280 12328
rect 26510 12316 26516 12328
rect 26568 12316 26574 12368
rect 26007 12260 26096 12288
rect 26237 12291 26295 12297
rect 26007 12257 26019 12260
rect 25961 12251 26019 12257
rect 26237 12257 26249 12291
rect 26283 12257 26295 12291
rect 26237 12251 26295 12257
rect 23109 12223 23167 12229
rect 23109 12220 23121 12223
rect 20180 12192 20944 12220
rect 20916 12164 20944 12192
rect 22572 12192 23121 12220
rect 17236 12124 18828 12152
rect 15010 12084 15016 12096
rect 14783 12056 15016 12084
rect 14783 12053 14795 12056
rect 14737 12047 14795 12053
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 15562 12044 15568 12096
rect 15620 12084 15626 12096
rect 16209 12087 16267 12093
rect 16209 12084 16221 12087
rect 15620 12056 16221 12084
rect 15620 12044 15626 12056
rect 16209 12053 16221 12056
rect 16255 12053 16267 12087
rect 16209 12047 16267 12053
rect 16482 12044 16488 12096
rect 16540 12044 16546 12096
rect 16850 12044 16856 12096
rect 16908 12084 16914 12096
rect 17236 12084 17264 12124
rect 18874 12112 18880 12164
rect 18932 12152 18938 12164
rect 19797 12155 19855 12161
rect 19797 12152 19809 12155
rect 18932 12124 19809 12152
rect 18932 12112 18938 12124
rect 19797 12121 19809 12124
rect 19843 12121 19855 12155
rect 19797 12115 19855 12121
rect 20898 12112 20904 12164
rect 20956 12112 20962 12164
rect 16908 12056 17264 12084
rect 17313 12087 17371 12093
rect 16908 12044 16914 12056
rect 17313 12053 17325 12087
rect 17359 12084 17371 12087
rect 18046 12084 18052 12096
rect 17359 12056 18052 12084
rect 17359 12053 17371 12056
rect 17313 12047 17371 12053
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 19518 12044 19524 12096
rect 19576 12044 19582 12096
rect 20070 12044 20076 12096
rect 20128 12044 20134 12096
rect 20530 12044 20536 12096
rect 20588 12044 20594 12096
rect 22186 12044 22192 12096
rect 22244 12084 22250 12096
rect 22572 12093 22600 12192
rect 23109 12189 23121 12192
rect 23155 12189 23167 12223
rect 23109 12183 23167 12189
rect 25516 12220 25544 12251
rect 26326 12248 26332 12300
rect 26384 12248 26390 12300
rect 26344 12220 26372 12248
rect 25516 12192 26372 12220
rect 24670 12112 24676 12164
rect 24728 12152 24734 12164
rect 25041 12155 25099 12161
rect 25041 12152 25053 12155
rect 24728 12124 25053 12152
rect 24728 12112 24734 12124
rect 25041 12121 25053 12124
rect 25087 12121 25099 12155
rect 25041 12115 25099 12121
rect 22557 12087 22615 12093
rect 22557 12084 22569 12087
rect 22244 12056 22569 12084
rect 22244 12044 22250 12056
rect 22557 12053 22569 12056
rect 22603 12053 22615 12087
rect 22557 12047 22615 12053
rect 24486 12044 24492 12096
rect 24544 12084 24550 12096
rect 25516 12084 25544 12192
rect 24544 12056 25544 12084
rect 24544 12044 24550 12056
rect 25590 12044 25596 12096
rect 25648 12044 25654 12096
rect 552 11994 31372 12016
rect 552 11942 4250 11994
rect 4302 11942 4314 11994
rect 4366 11942 4378 11994
rect 4430 11942 4442 11994
rect 4494 11942 4506 11994
rect 4558 11942 11955 11994
rect 12007 11942 12019 11994
rect 12071 11942 12083 11994
rect 12135 11942 12147 11994
rect 12199 11942 12211 11994
rect 12263 11942 19660 11994
rect 19712 11942 19724 11994
rect 19776 11942 19788 11994
rect 19840 11942 19852 11994
rect 19904 11942 19916 11994
rect 19968 11942 27365 11994
rect 27417 11942 27429 11994
rect 27481 11942 27493 11994
rect 27545 11942 27557 11994
rect 27609 11942 27621 11994
rect 27673 11942 31372 11994
rect 552 11920 31372 11942
rect 7607 11883 7665 11889
rect 7607 11849 7619 11883
rect 7653 11880 7665 11883
rect 9214 11880 9220 11892
rect 7653 11852 8892 11880
rect 7653 11849 7665 11852
rect 7607 11843 7665 11849
rect 8435 11815 8493 11821
rect 8435 11812 8447 11815
rect 7668 11784 8447 11812
rect 7536 11679 7594 11685
rect 7536 11645 7548 11679
rect 7582 11676 7594 11679
rect 7668 11676 7696 11784
rect 8435 11781 8447 11784
rect 8481 11781 8493 11815
rect 8435 11775 8493 11781
rect 8711 11747 8769 11753
rect 8711 11744 8723 11747
rect 8404 11716 8723 11744
rect 7582 11648 7696 11676
rect 7582 11645 7594 11648
rect 7536 11639 7594 11645
rect 7742 11636 7748 11688
rect 7800 11685 7806 11688
rect 7800 11679 7838 11685
rect 7826 11645 7838 11679
rect 7800 11639 7838 11645
rect 8088 11679 8146 11685
rect 8088 11645 8100 11679
rect 8134 11676 8146 11679
rect 8404 11676 8432 11716
rect 8711 11713 8723 11716
rect 8757 11713 8769 11747
rect 8711 11707 8769 11713
rect 8864 11685 8892 11852
rect 8956 11852 9220 11880
rect 8956 11685 8984 11852
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 10744 11852 11100 11880
rect 10744 11840 10750 11852
rect 9033 11815 9091 11821
rect 9033 11781 9045 11815
rect 9079 11812 9091 11815
rect 9079 11784 9628 11812
rect 9079 11781 9091 11784
rect 9033 11775 9091 11781
rect 9398 11704 9404 11756
rect 9456 11704 9462 11756
rect 8506 11679 8564 11685
rect 8506 11676 8518 11679
rect 8134 11648 8432 11676
rect 8134 11645 8146 11648
rect 8088 11639 8146 11645
rect 8496 11645 8518 11676
rect 8552 11645 8564 11679
rect 8496 11639 8564 11645
rect 8814 11679 8892 11685
rect 8814 11645 8826 11679
rect 8860 11648 8892 11679
rect 8941 11679 8999 11685
rect 8860 11645 8872 11648
rect 8814 11639 8872 11645
rect 8941 11645 8953 11679
rect 8987 11645 8999 11679
rect 8941 11639 8999 11645
rect 7800 11636 7806 11639
rect 7883 11611 7941 11617
rect 7883 11577 7895 11611
rect 7929 11608 7941 11611
rect 8496 11608 8524 11639
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 9252 11687 9310 11693
rect 9252 11684 9264 11687
rect 9232 11676 9264 11684
rect 9088 11653 9264 11676
rect 9298 11653 9310 11687
rect 9088 11648 9310 11653
rect 9088 11636 9094 11648
rect 9252 11647 9310 11648
rect 9416 11608 9444 11704
rect 7929 11580 8524 11608
rect 8772 11580 9444 11608
rect 9600 11608 9628 11784
rect 9674 11636 9680 11688
rect 9732 11636 9738 11688
rect 9950 11636 9956 11688
rect 10008 11636 10014 11688
rect 10042 11636 10048 11688
rect 10100 11636 10106 11688
rect 10290 11611 10348 11617
rect 10290 11608 10302 11611
rect 9600 11580 10302 11608
rect 7929 11577 7941 11580
rect 7883 11571 7941 11577
rect 8159 11543 8217 11549
rect 8159 11509 8171 11543
rect 8205 11540 8217 11543
rect 8772 11540 8800 11580
rect 10290 11577 10302 11580
rect 10336 11577 10348 11611
rect 11072 11608 11100 11852
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 11425 11883 11483 11889
rect 11425 11880 11437 11883
rect 11388 11852 11437 11880
rect 11388 11840 11394 11852
rect 11425 11849 11437 11852
rect 11471 11849 11483 11883
rect 11425 11843 11483 11849
rect 11698 11840 11704 11892
rect 11756 11840 11762 11892
rect 13725 11883 13783 11889
rect 13725 11849 13737 11883
rect 13771 11880 13783 11883
rect 13906 11880 13912 11892
rect 13771 11852 13912 11880
rect 13771 11849 13783 11852
rect 13725 11843 13783 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 14001 11883 14059 11889
rect 14001 11849 14013 11883
rect 14047 11849 14059 11883
rect 14001 11843 14059 11849
rect 14277 11883 14335 11889
rect 14277 11849 14289 11883
rect 14323 11880 14335 11883
rect 15194 11880 15200 11892
rect 14323 11852 15200 11880
rect 14323 11849 14335 11852
rect 14277 11843 14335 11849
rect 14016 11812 14044 11843
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 15381 11883 15439 11889
rect 15381 11849 15393 11883
rect 15427 11880 15439 11883
rect 15470 11880 15476 11892
rect 15427 11852 15476 11880
rect 15427 11849 15439 11852
rect 15381 11843 15439 11849
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 15654 11840 15660 11892
rect 15712 11880 15718 11892
rect 16301 11883 16359 11889
rect 16301 11880 16313 11883
rect 15712 11852 16313 11880
rect 15712 11840 15718 11852
rect 16301 11849 16313 11852
rect 16347 11849 16359 11883
rect 17218 11880 17224 11892
rect 16301 11843 16359 11849
rect 16408 11852 17224 11880
rect 14553 11815 14611 11821
rect 14016 11784 14504 11812
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13998 11744 14004 11756
rect 13127 11716 14004 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14090 11704 14096 11756
rect 14148 11704 14154 11756
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 13265 11679 13323 11685
rect 13265 11645 13277 11679
rect 13311 11676 13323 11679
rect 13633 11679 13691 11685
rect 13633 11676 13645 11679
rect 13311 11648 13645 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 13633 11645 13645 11648
rect 13679 11645 13691 11679
rect 13633 11639 13691 11645
rect 12814 11611 12872 11617
rect 12814 11608 12826 11611
rect 11072 11580 12826 11608
rect 10290 11571 10348 11577
rect 12814 11577 12826 11580
rect 12860 11577 12872 11611
rect 13188 11608 13216 11639
rect 13814 11636 13820 11688
rect 13872 11636 13878 11688
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14108 11676 14136 11704
rect 14476 11685 14504 11784
rect 14553 11781 14565 11815
rect 14599 11812 14611 11815
rect 14918 11812 14924 11824
rect 14599 11784 14924 11812
rect 14599 11781 14611 11784
rect 14553 11775 14611 11781
rect 14918 11772 14924 11784
rect 14976 11772 14982 11824
rect 16408 11812 16436 11852
rect 17218 11840 17224 11852
rect 17276 11840 17282 11892
rect 18417 11883 18475 11889
rect 18417 11849 18429 11883
rect 18463 11880 18475 11883
rect 18506 11880 18512 11892
rect 18463 11852 18512 11880
rect 18463 11849 18475 11852
rect 18417 11843 18475 11849
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 20257 11883 20315 11889
rect 20257 11849 20269 11883
rect 20303 11880 20315 11883
rect 20346 11880 20352 11892
rect 20303 11852 20352 11880
rect 20303 11849 20315 11852
rect 20257 11843 20315 11849
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 20530 11840 20536 11892
rect 20588 11840 20594 11892
rect 20622 11840 20628 11892
rect 20680 11880 20686 11892
rect 20809 11883 20867 11889
rect 20809 11880 20821 11883
rect 20680 11852 20821 11880
rect 20680 11840 20686 11852
rect 20809 11849 20821 11852
rect 20855 11849 20867 11883
rect 20809 11843 20867 11849
rect 21082 11840 21088 11892
rect 21140 11840 21146 11892
rect 24489 11883 24547 11889
rect 24489 11880 24501 11883
rect 21192 11852 24501 11880
rect 15212 11784 16436 11812
rect 13955 11648 14136 11676
rect 14185 11679 14243 11685
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 14185 11645 14197 11679
rect 14231 11645 14243 11679
rect 14185 11639 14243 11645
rect 14461 11679 14519 11685
rect 14461 11645 14473 11679
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 13538 11608 13544 11620
rect 13188 11580 13544 11608
rect 12814 11571 12872 11577
rect 13538 11568 13544 11580
rect 13596 11608 13602 11620
rect 14200 11608 14228 11639
rect 14918 11636 14924 11688
rect 14976 11636 14982 11688
rect 15010 11636 15016 11688
rect 15068 11670 15074 11688
rect 15212 11670 15240 11784
rect 15654 11704 15660 11756
rect 15712 11704 15718 11756
rect 15068 11642 15240 11670
rect 15068 11636 15074 11642
rect 15470 11636 15476 11688
rect 15528 11636 15534 11688
rect 15565 11679 15623 11685
rect 15565 11645 15577 11679
rect 15611 11676 15623 11679
rect 15764 11676 15792 11784
rect 15856 11716 16160 11744
rect 15856 11688 15884 11716
rect 15611 11648 15792 11676
rect 15611 11645 15623 11648
rect 15565 11639 15623 11645
rect 15838 11636 15844 11688
rect 15896 11636 15902 11688
rect 16025 11679 16083 11685
rect 16025 11645 16037 11679
rect 16071 11645 16083 11679
rect 16025 11639 16083 11645
rect 15286 11608 15292 11620
rect 13596 11580 15292 11608
rect 13596 11568 13602 11580
rect 15286 11568 15292 11580
rect 15344 11568 15350 11620
rect 15933 11611 15991 11617
rect 15933 11577 15945 11611
rect 15979 11577 15991 11611
rect 15933 11571 15991 11577
rect 8205 11512 8800 11540
rect 9355 11543 9413 11549
rect 8205 11509 8217 11512
rect 8159 11503 8217 11509
rect 9355 11509 9367 11543
rect 9401 11540 9413 11543
rect 9490 11540 9496 11552
rect 9401 11512 9496 11540
rect 9401 11509 9413 11512
rect 9355 11503 9413 11509
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 9582 11500 9588 11552
rect 9640 11500 9646 11552
rect 9858 11500 9864 11552
rect 9916 11500 9922 11552
rect 14826 11500 14832 11552
rect 14884 11500 14890 11552
rect 15102 11500 15108 11552
rect 15160 11500 15166 11552
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 15948 11540 15976 11571
rect 15528 11512 15976 11540
rect 16040 11540 16068 11639
rect 16132 11608 16160 11716
rect 16408 11685 16436 11784
rect 16577 11815 16635 11821
rect 16577 11781 16589 11815
rect 16623 11812 16635 11815
rect 16666 11812 16672 11824
rect 16623 11784 16672 11812
rect 16623 11781 16635 11784
rect 16577 11775 16635 11781
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11744 16911 11747
rect 17034 11744 17040 11756
rect 16899 11716 17040 11744
rect 16899 11713 16911 11716
rect 16853 11707 16911 11713
rect 17034 11704 17040 11716
rect 17092 11744 17098 11756
rect 18693 11747 18751 11753
rect 18693 11744 18705 11747
rect 17092 11716 18705 11744
rect 17092 11704 17098 11716
rect 18693 11713 18705 11716
rect 18739 11713 18751 11747
rect 18693 11707 18751 11713
rect 18874 11704 18880 11756
rect 18932 11704 18938 11756
rect 21192 11744 21220 11852
rect 24489 11849 24501 11852
rect 24535 11849 24547 11883
rect 24489 11843 24547 11849
rect 24762 11840 24768 11892
rect 24820 11840 24826 11892
rect 25498 11880 25504 11892
rect 25332 11852 25504 11880
rect 21266 11772 21272 11824
rect 21324 11812 21330 11824
rect 21637 11815 21695 11821
rect 21637 11812 21649 11815
rect 21324 11784 21649 11812
rect 21324 11772 21330 11784
rect 21637 11781 21649 11784
rect 21683 11781 21695 11815
rect 25332 11812 25360 11852
rect 25498 11840 25504 11852
rect 25556 11840 25562 11892
rect 25590 11840 25596 11892
rect 25648 11880 25654 11892
rect 25648 11852 26096 11880
rect 25648 11840 25654 11852
rect 25869 11815 25927 11821
rect 25869 11812 25881 11815
rect 21637 11775 21695 11781
rect 23952 11784 25360 11812
rect 25424 11784 25881 11812
rect 21913 11747 21971 11753
rect 21913 11744 21925 11747
rect 19996 11716 21220 11744
rect 21376 11716 21925 11744
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 16669 11679 16727 11685
rect 16669 11645 16681 11679
rect 16715 11645 16727 11679
rect 16669 11639 16727 11645
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 18892 11676 18920 11704
rect 17175 11648 18920 11676
rect 18969 11679 19027 11685
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 18969 11645 18981 11679
rect 19015 11676 19027 11679
rect 19702 11676 19708 11688
rect 19015 11648 19708 11676
rect 19015 11645 19027 11648
rect 18969 11639 19027 11645
rect 16684 11608 16712 11639
rect 19702 11636 19708 11648
rect 19760 11636 19766 11688
rect 16132 11580 16712 11608
rect 19996 11552 20024 11716
rect 20625 11679 20683 11685
rect 20625 11645 20637 11679
rect 20671 11645 20683 11679
rect 20625 11639 20683 11645
rect 20901 11679 20959 11685
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 20990 11676 20996 11688
rect 20947 11648 20996 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 20640 11608 20668 11639
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 21177 11679 21235 11685
rect 21177 11645 21189 11679
rect 21223 11676 21235 11679
rect 21376 11676 21404 11716
rect 21913 11713 21925 11716
rect 21959 11713 21971 11747
rect 21913 11707 21971 11713
rect 21223 11648 21404 11676
rect 21453 11679 21511 11685
rect 21223 11645 21235 11648
rect 21177 11639 21235 11645
rect 21453 11645 21465 11679
rect 21499 11676 21511 11679
rect 21542 11676 21548 11688
rect 21499 11648 21548 11676
rect 21499 11645 21511 11648
rect 21453 11639 21511 11645
rect 21542 11636 21548 11648
rect 21600 11636 21606 11688
rect 21634 11636 21640 11688
rect 21692 11676 21698 11688
rect 21729 11679 21787 11685
rect 21729 11676 21741 11679
rect 21692 11648 21741 11676
rect 21692 11636 21698 11648
rect 21729 11645 21741 11648
rect 21775 11645 21787 11679
rect 21729 11639 21787 11645
rect 21818 11636 21824 11688
rect 21876 11636 21882 11688
rect 22186 11636 22192 11688
rect 22244 11636 22250 11688
rect 22456 11679 22514 11685
rect 22456 11645 22468 11679
rect 22502 11676 22514 11679
rect 23952 11676 23980 11784
rect 22502 11648 23980 11676
rect 24029 11689 24087 11695
rect 24029 11655 24041 11689
rect 24075 11655 24087 11689
rect 24029 11649 24087 11655
rect 22502 11645 22514 11648
rect 22456 11639 22514 11645
rect 24044 11620 24072 11649
rect 24302 11636 24308 11688
rect 24360 11676 24366 11688
rect 24486 11676 24492 11688
rect 24360 11648 24492 11676
rect 24360 11636 24366 11648
rect 24486 11636 24492 11648
rect 24544 11636 24550 11688
rect 24581 11679 24639 11685
rect 24581 11645 24593 11679
rect 24627 11645 24639 11679
rect 24581 11639 24639 11645
rect 21361 11611 21419 11617
rect 21361 11608 21373 11611
rect 20640 11580 21373 11608
rect 21361 11577 21373 11580
rect 21407 11577 21419 11611
rect 23937 11611 23995 11617
rect 23937 11608 23949 11611
rect 21361 11571 21419 11577
rect 21560 11580 22094 11608
rect 21560 11552 21588 11580
rect 16666 11540 16672 11552
rect 16040 11512 16672 11540
rect 15528 11500 15534 11512
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 19978 11500 19984 11552
rect 20036 11500 20042 11552
rect 21542 11500 21548 11552
rect 21600 11500 21606 11552
rect 22066 11540 22094 11580
rect 22572 11580 23949 11608
rect 22572 11540 22600 11580
rect 23937 11577 23949 11580
rect 23983 11577 23995 11611
rect 23937 11571 23995 11577
rect 24026 11568 24032 11620
rect 24084 11568 24090 11620
rect 22066 11512 22600 11540
rect 23569 11543 23627 11549
rect 23569 11509 23581 11543
rect 23615 11540 23627 11543
rect 24118 11540 24124 11552
rect 23615 11512 24124 11540
rect 23615 11509 23627 11512
rect 23569 11503 23627 11509
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 24210 11500 24216 11552
rect 24268 11500 24274 11552
rect 24596 11540 24624 11639
rect 24670 11636 24676 11688
rect 24728 11636 24734 11688
rect 24857 11679 24915 11685
rect 24857 11645 24869 11679
rect 24903 11645 24915 11679
rect 24857 11639 24915 11645
rect 24872 11608 24900 11639
rect 25038 11636 25044 11688
rect 25096 11676 25102 11688
rect 25424 11685 25452 11784
rect 25869 11781 25881 11784
rect 25915 11781 25927 11815
rect 25869 11775 25927 11781
rect 25700 11716 26004 11744
rect 25700 11685 25728 11716
rect 25976 11688 26004 11716
rect 25133 11679 25191 11685
rect 25133 11676 25145 11679
rect 25096 11648 25145 11676
rect 25096 11636 25102 11648
rect 25133 11645 25145 11648
rect 25179 11645 25191 11679
rect 25133 11639 25191 11645
rect 25409 11679 25467 11685
rect 25409 11645 25421 11679
rect 25455 11645 25467 11679
rect 25409 11639 25467 11645
rect 25685 11679 25743 11685
rect 25685 11645 25697 11679
rect 25731 11645 25743 11679
rect 25685 11639 25743 11645
rect 25777 11679 25835 11685
rect 25777 11645 25789 11679
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 25593 11611 25651 11617
rect 25593 11608 25605 11611
rect 24872 11580 25605 11608
rect 25593 11577 25605 11580
rect 25639 11577 25651 11611
rect 25792 11608 25820 11639
rect 25958 11636 25964 11688
rect 26016 11636 26022 11688
rect 26068 11685 26096 11852
rect 26053 11679 26111 11685
rect 26053 11645 26065 11679
rect 26099 11645 26111 11679
rect 26053 11639 26111 11645
rect 25593 11571 25651 11577
rect 25700 11580 25820 11608
rect 25041 11543 25099 11549
rect 25041 11540 25053 11543
rect 24596 11512 25053 11540
rect 25041 11509 25053 11512
rect 25087 11509 25099 11543
rect 25041 11503 25099 11509
rect 25130 11500 25136 11552
rect 25188 11540 25194 11552
rect 25317 11543 25375 11549
rect 25317 11540 25329 11543
rect 25188 11512 25329 11540
rect 25188 11500 25194 11512
rect 25317 11509 25329 11512
rect 25363 11509 25375 11543
rect 25317 11503 25375 11509
rect 25406 11500 25412 11552
rect 25464 11540 25470 11552
rect 25700 11540 25728 11580
rect 25866 11568 25872 11620
rect 25924 11608 25930 11620
rect 26145 11611 26203 11617
rect 26145 11608 26157 11611
rect 25924 11580 26157 11608
rect 25924 11568 25930 11580
rect 26145 11577 26157 11580
rect 26191 11577 26203 11611
rect 26145 11571 26203 11577
rect 25464 11512 25728 11540
rect 25464 11500 25470 11512
rect 552 11450 31531 11472
rect 552 11398 8102 11450
rect 8154 11398 8166 11450
rect 8218 11398 8230 11450
rect 8282 11398 8294 11450
rect 8346 11398 8358 11450
rect 8410 11398 15807 11450
rect 15859 11398 15871 11450
rect 15923 11398 15935 11450
rect 15987 11398 15999 11450
rect 16051 11398 16063 11450
rect 16115 11398 23512 11450
rect 23564 11398 23576 11450
rect 23628 11398 23640 11450
rect 23692 11398 23704 11450
rect 23756 11398 23768 11450
rect 23820 11398 31217 11450
rect 31269 11398 31281 11450
rect 31333 11398 31345 11450
rect 31397 11398 31409 11450
rect 31461 11398 31473 11450
rect 31525 11398 31531 11450
rect 552 11376 31531 11398
rect 7742 11296 7748 11348
rect 7800 11336 7806 11348
rect 10042 11336 10048 11348
rect 7800 11308 10048 11336
rect 7800 11296 7806 11308
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10336 11308 11468 11336
rect 10134 11268 10140 11280
rect 8864 11240 10140 11268
rect 8110 11160 8116 11212
rect 8168 11160 8174 11212
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 6178 11092 6184 11144
rect 6236 11132 6242 11144
rect 8404 11132 8432 11163
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 8864 11209 8892 11240
rect 9692 11209 9720 11240
rect 10134 11228 10140 11240
rect 10192 11228 10198 11280
rect 10336 11209 10364 11308
rect 10413 11271 10471 11277
rect 10413 11237 10425 11271
rect 10459 11268 10471 11271
rect 10459 11240 11008 11268
rect 10459 11237 10471 11240
rect 10413 11231 10471 11237
rect 10980 11209 11008 11240
rect 11440 11209 11468 11308
rect 11606 11296 11612 11348
rect 11664 11296 11670 11348
rect 12434 11336 12440 11348
rect 11992 11308 12440 11336
rect 11992 11268 12020 11308
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 14366 11296 14372 11348
rect 14424 11336 14430 11348
rect 14553 11339 14611 11345
rect 14553 11336 14565 11339
rect 14424 11308 14565 11336
rect 14424 11296 14430 11308
rect 14553 11305 14565 11308
rect 14599 11305 14611 11339
rect 14553 11299 14611 11305
rect 15562 11296 15568 11348
rect 15620 11296 15626 11348
rect 15657 11339 15715 11345
rect 15657 11305 15669 11339
rect 15703 11336 15715 11339
rect 16298 11336 16304 11348
rect 15703 11308 16304 11336
rect 15703 11305 15715 11308
rect 15657 11299 15715 11305
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 16482 11296 16488 11348
rect 16540 11296 16546 11348
rect 17218 11296 17224 11348
rect 17276 11296 17282 11348
rect 18046 11296 18052 11348
rect 18104 11296 18110 11348
rect 18230 11296 18236 11348
rect 18288 11296 18294 11348
rect 19426 11296 19432 11348
rect 19484 11296 19490 11348
rect 19518 11296 19524 11348
rect 19576 11296 19582 11348
rect 19702 11296 19708 11348
rect 19760 11296 19766 11348
rect 20070 11296 20076 11348
rect 20128 11296 20134 11348
rect 24210 11336 24216 11348
rect 20180 11308 24216 11336
rect 11532 11240 12020 11268
rect 12176 11240 12388 11268
rect 11532 11209 11560 11240
rect 8849 11203 8907 11209
rect 8849 11200 8861 11203
rect 8536 11172 8861 11200
rect 8536 11160 8542 11172
rect 8849 11169 8861 11172
rect 8895 11169 8907 11203
rect 8849 11163 8907 11169
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11200 9183 11203
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 9171 11172 9321 11200
rect 9171 11169 9183 11172
rect 9125 11163 9183 11169
rect 9309 11169 9321 11172
rect 9355 11169 9367 11203
rect 9309 11163 9367 11169
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 9953 11203 10011 11209
rect 9953 11169 9965 11203
rect 9999 11200 10011 11203
rect 10229 11203 10287 11209
rect 9999 11172 10088 11200
rect 9999 11169 10011 11172
rect 9953 11163 10011 11169
rect 6236 11104 8432 11132
rect 6236 11092 6242 11104
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 9033 11135 9091 11141
rect 9033 11132 9045 11135
rect 8628 11104 9045 11132
rect 8628 11092 8634 11104
rect 9033 11101 9045 11104
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9416 11132 9444 11163
rect 10060 11132 10088 11172
rect 10229 11169 10241 11203
rect 10275 11200 10287 11203
rect 10321 11203 10379 11209
rect 10321 11200 10333 11203
rect 10275 11172 10333 11200
rect 10275 11169 10287 11172
rect 10229 11163 10287 11169
rect 10321 11169 10333 11172
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11169 11483 11203
rect 11425 11163 11483 11169
rect 11517 11203 11575 11209
rect 11517 11169 11529 11203
rect 11563 11169 11575 11203
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11517 11163 11575 11169
rect 11716 11172 11989 11200
rect 10410 11132 10416 11144
rect 9272 11104 9996 11132
rect 10060 11104 10416 11132
rect 9272 11092 9278 11104
rect 9968 11076 9996 11104
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 8205 11067 8263 11073
rect 8205 11033 8217 11067
rect 8251 11064 8263 11067
rect 8481 11067 8539 11073
rect 8481 11064 8493 11067
rect 8251 11036 8493 11064
rect 8251 11033 8263 11036
rect 8205 11027 8263 11033
rect 8481 11033 8493 11036
rect 8527 11033 8539 11067
rect 8481 11027 8539 11033
rect 8938 11024 8944 11076
rect 8996 11064 9002 11076
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 8996 11036 9873 11064
rect 8996 11024 9002 11036
rect 9861 11033 9873 11036
rect 9907 11033 9919 11067
rect 9861 11027 9919 11033
rect 9950 11024 9956 11076
rect 10008 11064 10014 11076
rect 10612 11064 10640 11163
rect 11440 11132 11468 11163
rect 11440 11104 11652 11132
rect 11624 11076 11652 11104
rect 11716 11076 11744 11172
rect 11977 11169 11989 11172
rect 12023 11200 12035 11203
rect 12176 11200 12204 11240
rect 12360 11209 12388 11240
rect 13188 11240 14044 11268
rect 13188 11209 13216 11240
rect 14016 11212 14044 11240
rect 13446 11209 13452 11212
rect 12023 11172 12204 11200
rect 12253 11203 12311 11209
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 12253 11169 12265 11203
rect 12299 11169 12311 11203
rect 12253 11163 12311 11169
rect 12345 11203 12403 11209
rect 12345 11169 12357 11203
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11200 12495 11203
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 12483 11172 12633 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 12621 11169 12633 11172
rect 12667 11169 12679 11203
rect 12621 11163 12679 11169
rect 12897 11203 12955 11209
rect 12897 11169 12909 11203
rect 12943 11200 12955 11203
rect 13173 11203 13231 11209
rect 12943 11172 13124 11200
rect 12943 11169 12955 11172
rect 12897 11163 12955 11169
rect 12268 11132 12296 11163
rect 12526 11132 12532 11144
rect 12268 11104 12532 11132
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 10008 11036 10640 11064
rect 10008 11024 10014 11036
rect 10336 11008 10364 11036
rect 11330 11024 11336 11076
rect 11388 11024 11394 11076
rect 11606 11024 11612 11076
rect 11664 11024 11670 11076
rect 11698 11024 11704 11076
rect 11756 11064 11762 11076
rect 12161 11067 12219 11073
rect 11756 11036 12112 11064
rect 11756 11024 11762 11036
rect 8754 10956 8760 11008
rect 8812 10956 8818 11008
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9585 10999 9643 11005
rect 9585 10996 9597 10999
rect 9180 10968 9597 10996
rect 9180 10956 9186 10968
rect 9585 10965 9597 10968
rect 9631 10965 9643 10999
rect 9585 10959 9643 10965
rect 10134 10956 10140 11008
rect 10192 10956 10198 11008
rect 10318 10956 10324 11008
rect 10376 10956 10382 11008
rect 10686 10956 10692 11008
rect 10744 10956 10750 11008
rect 11054 10956 11060 11008
rect 11112 10956 11118 11008
rect 11238 10956 11244 11008
rect 11296 10996 11302 11008
rect 11885 10999 11943 11005
rect 11885 10996 11897 10999
rect 11296 10968 11897 10996
rect 11296 10956 11302 10968
rect 11885 10965 11897 10968
rect 11931 10965 11943 10999
rect 12084 10996 12112 11036
rect 12161 11033 12173 11067
rect 12207 11064 12219 11067
rect 12713 11067 12771 11073
rect 12713 11064 12725 11067
rect 12207 11036 12725 11064
rect 12207 11033 12219 11036
rect 12161 11027 12219 11033
rect 12713 11033 12725 11036
rect 12759 11033 12771 11067
rect 13096 11064 13124 11172
rect 13173 11169 13185 11203
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 13429 11203 13452 11209
rect 13429 11169 13441 11203
rect 13429 11163 13452 11169
rect 13446 11160 13452 11163
rect 13504 11160 13510 11212
rect 13998 11160 14004 11212
rect 14056 11160 14062 11212
rect 15105 11203 15163 11209
rect 15105 11169 15117 11203
rect 15151 11200 15163 11203
rect 15286 11200 15292 11212
rect 15151 11172 15292 11200
rect 15151 11169 15163 11172
rect 15105 11163 15163 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15378 11160 15384 11212
rect 15436 11160 15442 11212
rect 15473 11203 15531 11209
rect 15473 11169 15485 11203
rect 15519 11200 15531 11203
rect 15580 11200 15608 11296
rect 16500 11268 16528 11296
rect 15672 11240 16528 11268
rect 17236 11268 17264 11296
rect 17236 11240 18000 11268
rect 15672 11209 15700 11240
rect 15519 11172 15608 11200
rect 15657 11203 15715 11209
rect 15519 11169 15531 11172
rect 15473 11163 15531 11169
rect 15657 11169 15669 11203
rect 15703 11169 15715 11203
rect 15657 11163 15715 11169
rect 15933 11203 15991 11209
rect 15933 11169 15945 11203
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 15948 11132 15976 11163
rect 16114 11160 16120 11212
rect 16172 11160 16178 11212
rect 16482 11160 16488 11212
rect 16540 11200 16546 11212
rect 17972 11209 18000 11240
rect 17957 11203 18015 11209
rect 16540 11172 17908 11200
rect 16540 11160 16546 11172
rect 16850 11132 16856 11144
rect 15948 11104 16856 11132
rect 16850 11092 16856 11104
rect 16908 11092 16914 11144
rect 17880 11132 17908 11172
rect 17957 11169 17969 11203
rect 18003 11169 18015 11203
rect 18064 11200 18092 11296
rect 19536 11268 19564 11296
rect 20088 11268 20116 11296
rect 18616 11240 18828 11268
rect 18233 11203 18291 11209
rect 18233 11200 18245 11203
rect 18064 11172 18245 11200
rect 17957 11163 18015 11169
rect 18233 11169 18245 11172
rect 18279 11169 18291 11203
rect 18233 11163 18291 11169
rect 18417 11203 18475 11209
rect 18417 11169 18429 11203
rect 18463 11169 18475 11203
rect 18417 11163 18475 11169
rect 18432 11132 18460 11163
rect 17880 11104 18460 11132
rect 12713 11027 12771 11033
rect 12912 11036 13124 11064
rect 12912 10996 12940 11036
rect 12084 10968 12940 10996
rect 11885 10959 11943 10965
rect 12986 10956 12992 11008
rect 13044 10956 13050 11008
rect 13096 10996 13124 11036
rect 15013 11067 15071 11073
rect 15013 11033 15025 11067
rect 15059 11064 15071 11067
rect 15470 11064 15476 11076
rect 15059 11036 15476 11064
rect 15059 11033 15071 11036
rect 15013 11027 15071 11033
rect 15470 11024 15476 11036
rect 15528 11024 15534 11076
rect 15764 11036 16068 11064
rect 14090 10996 14096 11008
rect 13096 10968 14096 10996
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 15289 10999 15347 11005
rect 15289 10965 15301 10999
rect 15335 10996 15347 10999
rect 15764 10996 15792 11036
rect 15335 10968 15792 10996
rect 15335 10965 15347 10968
rect 15289 10959 15347 10965
rect 15838 10956 15844 11008
rect 15896 10956 15902 11008
rect 16040 10996 16068 11036
rect 16942 11024 16948 11076
rect 17000 11064 17006 11076
rect 17589 11067 17647 11073
rect 17589 11064 17601 11067
rect 17000 11036 17601 11064
rect 17000 11024 17006 11036
rect 17589 11033 17601 11036
rect 17635 11064 17647 11067
rect 17770 11064 17776 11076
rect 17635 11036 17776 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 17770 11024 17776 11036
rect 17828 11024 17834 11076
rect 18616 11064 18644 11240
rect 18800 11209 18828 11240
rect 19260 11240 19564 11268
rect 19812 11240 20116 11268
rect 19260 11209 19288 11240
rect 19812 11209 19840 11240
rect 18693 11203 18751 11209
rect 18693 11169 18705 11203
rect 18739 11169 18751 11203
rect 18693 11163 18751 11169
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11200 18843 11203
rect 19153 11203 19211 11209
rect 19153 11200 19165 11203
rect 18831 11172 19165 11200
rect 18831 11169 18843 11172
rect 18785 11163 18843 11169
rect 19153 11169 19165 11172
rect 19199 11169 19211 11203
rect 19153 11163 19211 11169
rect 19245 11203 19303 11209
rect 19245 11169 19257 11203
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 19337 11203 19395 11209
rect 19337 11169 19349 11203
rect 19383 11169 19395 11203
rect 19337 11163 19395 11169
rect 19797 11203 19855 11209
rect 19797 11169 19809 11203
rect 19843 11169 19855 11203
rect 19797 11163 19855 11169
rect 17972 11036 18644 11064
rect 18708 11064 18736 11163
rect 19168 11132 19196 11163
rect 19352 11132 19380 11163
rect 19978 11160 19984 11212
rect 20036 11160 20042 11212
rect 20180 11209 20208 11308
rect 24210 11296 24216 11308
rect 24268 11296 24274 11348
rect 24394 11296 24400 11348
rect 24452 11336 24458 11348
rect 25038 11336 25044 11348
rect 24452 11308 25044 11336
rect 24452 11296 24458 11308
rect 25038 11296 25044 11308
rect 25096 11336 25102 11348
rect 25406 11336 25412 11348
rect 25096 11308 25412 11336
rect 25096 11296 25102 11308
rect 25406 11296 25412 11308
rect 25464 11296 25470 11348
rect 20349 11271 20407 11277
rect 20349 11237 20361 11271
rect 20395 11268 20407 11271
rect 20395 11240 20944 11268
rect 20395 11237 20407 11240
rect 20349 11231 20407 11237
rect 20165 11203 20223 11209
rect 20165 11169 20177 11203
rect 20211 11169 20223 11203
rect 20165 11163 20223 11169
rect 20254 11160 20260 11212
rect 20312 11200 20318 11212
rect 20916 11209 20944 11240
rect 20990 11228 20996 11280
rect 21048 11268 21054 11280
rect 21726 11268 21732 11280
rect 21048 11240 21732 11268
rect 21048 11228 21054 11240
rect 21726 11228 21732 11240
rect 21784 11228 21790 11280
rect 23290 11228 23296 11280
rect 23348 11228 23354 11280
rect 23842 11268 23848 11280
rect 23676 11240 23848 11268
rect 20533 11203 20591 11209
rect 20533 11200 20545 11203
rect 20312 11172 20545 11200
rect 20312 11160 20318 11172
rect 20533 11169 20545 11172
rect 20579 11200 20591 11203
rect 20901 11203 20959 11209
rect 20579 11172 20852 11200
rect 20579 11169 20591 11172
rect 20533 11163 20591 11169
rect 19168 11104 19380 11132
rect 20625 11135 20683 11141
rect 20625 11101 20637 11135
rect 20671 11132 20683 11135
rect 20714 11132 20720 11144
rect 20671 11104 20720 11132
rect 20671 11101 20683 11104
rect 20625 11095 20683 11101
rect 20714 11092 20720 11104
rect 20772 11092 20778 11144
rect 20824 11132 20852 11172
rect 20901 11169 20913 11203
rect 20947 11169 20959 11203
rect 20901 11163 20959 11169
rect 21453 11203 21511 11209
rect 21453 11169 21465 11203
rect 21499 11200 21511 11203
rect 21542 11200 21548 11212
rect 21499 11172 21548 11200
rect 21499 11169 21511 11172
rect 21453 11163 21511 11169
rect 21542 11160 21548 11172
rect 21600 11160 21606 11212
rect 21637 11203 21695 11209
rect 21637 11169 21649 11203
rect 21683 11200 21695 11203
rect 22186 11200 22192 11212
rect 21683 11172 22192 11200
rect 21683 11169 21695 11172
rect 21637 11163 21695 11169
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 23385 11203 23443 11209
rect 23385 11169 23397 11203
rect 23431 11200 23443 11203
rect 23566 11200 23572 11212
rect 23431 11172 23572 11200
rect 23431 11169 23443 11172
rect 23385 11163 23443 11169
rect 23566 11160 23572 11172
rect 23624 11160 23630 11212
rect 23676 11209 23704 11240
rect 23842 11228 23848 11240
rect 23900 11228 23906 11280
rect 24118 11228 24124 11280
rect 24176 11268 24182 11280
rect 28258 11268 28264 11280
rect 24176 11240 28264 11268
rect 24176 11228 24182 11240
rect 28258 11228 28264 11240
rect 28316 11228 28322 11280
rect 23661 11203 23719 11209
rect 23661 11169 23673 11203
rect 23707 11169 23719 11203
rect 23661 11163 23719 11169
rect 23753 11203 23811 11209
rect 23753 11169 23765 11203
rect 23799 11200 23811 11203
rect 23937 11203 23995 11209
rect 23937 11200 23949 11203
rect 23799 11172 23949 11200
rect 23799 11169 23811 11172
rect 23753 11163 23811 11169
rect 23937 11169 23949 11172
rect 23983 11169 23995 11203
rect 23937 11163 23995 11169
rect 24210 11160 24216 11212
rect 24268 11200 24274 11212
rect 24397 11203 24455 11209
rect 24397 11200 24409 11203
rect 24268 11172 24409 11200
rect 24268 11160 24274 11172
rect 24397 11169 24409 11172
rect 24443 11169 24455 11203
rect 24397 11163 24455 11169
rect 24486 11160 24492 11212
rect 24544 11160 24550 11212
rect 24670 11160 24676 11212
rect 24728 11200 24734 11212
rect 24765 11203 24823 11209
rect 24765 11200 24777 11203
rect 24728 11172 24777 11200
rect 24728 11160 24734 11172
rect 24765 11169 24777 11172
rect 24811 11169 24823 11203
rect 24765 11163 24823 11169
rect 25222 11160 25228 11212
rect 25280 11160 25286 11212
rect 25317 11203 25375 11209
rect 25317 11169 25329 11203
rect 25363 11169 25375 11203
rect 25317 11163 25375 11169
rect 21913 11135 21971 11141
rect 20824 11104 21588 11132
rect 21560 11076 21588 11104
rect 21913 11101 21925 11135
rect 21959 11132 21971 11135
rect 25130 11132 25136 11144
rect 21959 11104 25136 11132
rect 21959 11101 21971 11104
rect 21913 11095 21971 11101
rect 25130 11092 25136 11104
rect 25188 11092 25194 11144
rect 19334 11064 19340 11076
rect 18708 11036 19340 11064
rect 16758 10996 16764 11008
rect 16040 10968 16764 10996
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 17126 10956 17132 11008
rect 17184 10996 17190 11008
rect 17972 10996 18000 11036
rect 19334 11024 19340 11036
rect 19392 11024 19398 11076
rect 20073 11067 20131 11073
rect 20073 11033 20085 11067
rect 20119 11064 20131 11067
rect 21450 11064 21456 11076
rect 20119 11036 21456 11064
rect 20119 11033 20131 11036
rect 20073 11027 20131 11033
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 21542 11024 21548 11076
rect 21600 11024 21606 11076
rect 23934 11024 23940 11076
rect 23992 11064 23998 11076
rect 25332 11064 25360 11163
rect 23992 11036 25360 11064
rect 23992 11024 23998 11036
rect 17184 10968 18000 10996
rect 17184 10956 17190 10968
rect 18046 10956 18052 11008
rect 18104 10956 18110 11008
rect 18598 10956 18604 11008
rect 18656 10956 18662 11008
rect 18874 10956 18880 11008
rect 18932 10956 18938 11008
rect 21174 10956 21180 11008
rect 21232 10996 21238 11008
rect 21361 10999 21419 11005
rect 21361 10996 21373 10999
rect 21232 10968 21373 10996
rect 21232 10956 21238 10968
rect 21361 10965 21373 10968
rect 21407 10996 21419 10999
rect 21634 10996 21640 11008
rect 21407 10968 21640 10996
rect 21407 10965 21419 10968
rect 21361 10959 21419 10965
rect 21634 10956 21640 10968
rect 21692 10956 21698 11008
rect 23474 10956 23480 11008
rect 23532 10956 23538 11008
rect 24026 10956 24032 11008
rect 24084 10956 24090 11008
rect 24302 10956 24308 11008
rect 24360 10956 24366 11008
rect 24578 10956 24584 11008
rect 24636 10956 24642 11008
rect 24854 10956 24860 11008
rect 24912 10956 24918 11008
rect 24946 10956 24952 11008
rect 25004 10996 25010 11008
rect 25133 10999 25191 11005
rect 25133 10996 25145 10999
rect 25004 10968 25145 10996
rect 25004 10956 25010 10968
rect 25133 10965 25145 10968
rect 25179 10965 25191 10999
rect 25133 10959 25191 10965
rect 25314 10956 25320 11008
rect 25372 10996 25378 11008
rect 25409 10999 25467 11005
rect 25409 10996 25421 10999
rect 25372 10968 25421 10996
rect 25372 10956 25378 10968
rect 25409 10965 25421 10968
rect 25455 10965 25467 10999
rect 25409 10959 25467 10965
rect 552 10906 31372 10928
rect 552 10854 4250 10906
rect 4302 10854 4314 10906
rect 4366 10854 4378 10906
rect 4430 10854 4442 10906
rect 4494 10854 4506 10906
rect 4558 10854 11955 10906
rect 12007 10854 12019 10906
rect 12071 10854 12083 10906
rect 12135 10854 12147 10906
rect 12199 10854 12211 10906
rect 12263 10854 19660 10906
rect 19712 10854 19724 10906
rect 19776 10854 19788 10906
rect 19840 10854 19852 10906
rect 19904 10854 19916 10906
rect 19968 10854 27365 10906
rect 27417 10854 27429 10906
rect 27481 10854 27493 10906
rect 27545 10854 27557 10906
rect 27609 10854 27621 10906
rect 27673 10854 31372 10906
rect 552 10832 31372 10854
rect 7561 10795 7619 10801
rect 7561 10761 7573 10795
rect 7607 10792 7619 10795
rect 8110 10792 8116 10804
rect 7607 10764 8116 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 8481 10795 8539 10801
rect 8481 10761 8493 10795
rect 8527 10792 8539 10795
rect 8938 10792 8944 10804
rect 8527 10764 8944 10792
rect 8527 10761 8539 10764
rect 8481 10755 8539 10761
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9122 10752 9128 10804
rect 9180 10752 9186 10804
rect 9585 10795 9643 10801
rect 9585 10761 9597 10795
rect 9631 10792 9643 10795
rect 11514 10792 11520 10804
rect 9631 10764 11520 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 13262 10752 13268 10804
rect 13320 10752 13326 10804
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16025 10795 16083 10801
rect 16025 10792 16037 10795
rect 15896 10764 16037 10792
rect 15896 10752 15902 10764
rect 16025 10761 16037 10764
rect 16071 10761 16083 10795
rect 16025 10755 16083 10761
rect 16206 10752 16212 10804
rect 16264 10752 16270 10804
rect 16574 10752 16580 10804
rect 16632 10752 16638 10804
rect 16850 10752 16856 10804
rect 16908 10752 16914 10804
rect 19334 10752 19340 10804
rect 19392 10752 19398 10804
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 21913 10795 21971 10801
rect 21913 10792 21925 10795
rect 20956 10764 21925 10792
rect 20956 10752 20962 10764
rect 21913 10761 21925 10764
rect 21959 10761 21971 10795
rect 21913 10755 21971 10761
rect 24026 10752 24032 10804
rect 24084 10792 24090 10804
rect 24213 10795 24271 10801
rect 24213 10792 24225 10795
rect 24084 10764 24225 10792
rect 24084 10752 24090 10764
rect 24213 10761 24225 10764
rect 24259 10761 24271 10795
rect 24213 10755 24271 10761
rect 24489 10795 24547 10801
rect 24489 10761 24501 10795
rect 24535 10792 24547 10795
rect 24670 10792 24676 10804
rect 24535 10764 24676 10792
rect 24535 10761 24547 10764
rect 24489 10755 24547 10761
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 24765 10795 24823 10801
rect 24765 10761 24777 10795
rect 24811 10792 24823 10795
rect 24854 10792 24860 10804
rect 24811 10764 24860 10792
rect 24811 10761 24823 10764
rect 24765 10755 24823 10761
rect 24854 10752 24860 10764
rect 24912 10752 24918 10804
rect 25222 10752 25228 10804
rect 25280 10792 25286 10804
rect 25317 10795 25375 10801
rect 25317 10792 25329 10795
rect 25280 10764 25329 10792
rect 25280 10752 25286 10764
rect 25317 10761 25329 10764
rect 25363 10761 25375 10795
rect 25317 10755 25375 10761
rect 9140 10724 9168 10752
rect 8588 10696 9168 10724
rect 8478 10656 8484 10668
rect 8220 10628 8484 10656
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 7650 10588 7656 10600
rect 7515 10560 7656 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 7929 10591 7987 10597
rect 7929 10557 7941 10591
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 7944 10520 7972 10551
rect 8018 10548 8024 10600
rect 8076 10588 8082 10600
rect 8220 10597 8248 10628
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 8588 10597 8616 10696
rect 9674 10684 9680 10736
rect 9732 10684 9738 10736
rect 10686 10724 10692 10736
rect 9968 10696 10692 10724
rect 9692 10656 9720 10684
rect 8680 10628 9720 10656
rect 8680 10597 8708 10628
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 8076 10560 8217 10588
rect 8076 10548 8082 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10557 8723 10591
rect 8665 10551 8723 10557
rect 8754 10548 8760 10600
rect 8812 10548 8818 10600
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9214 10588 9220 10600
rect 9171 10560 9220 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 9858 10588 9864 10600
rect 9723 10560 9864 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 8772 10520 8800 10548
rect 7944 10492 8800 10520
rect 9416 10520 9444 10551
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 9968 10597 9996 10696
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 15289 10727 15347 10733
rect 15289 10693 15301 10727
rect 15335 10724 15347 10727
rect 16224 10724 16252 10752
rect 15335 10696 16252 10724
rect 15335 10693 15347 10696
rect 15289 10687 15347 10693
rect 16592 10656 16620 10752
rect 18417 10727 18475 10733
rect 18417 10693 18429 10727
rect 18463 10724 18475 10727
rect 19426 10724 19432 10736
rect 18463 10696 19432 10724
rect 18463 10693 18475 10696
rect 18417 10687 18475 10693
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 20257 10727 20315 10733
rect 20257 10693 20269 10727
rect 20303 10724 20315 10727
rect 23569 10727 23627 10733
rect 20303 10696 21956 10724
rect 20303 10693 20315 10696
rect 20257 10687 20315 10693
rect 16132 10628 16620 10656
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10588 10103 10591
rect 10134 10588 10140 10600
rect 10091 10560 10140 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11793 10591 11851 10597
rect 11793 10588 11805 10591
rect 11204 10560 11805 10588
rect 11204 10548 11210 10560
rect 11793 10557 11805 10560
rect 11839 10588 11851 10591
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 11839 10560 11897 10588
rect 11839 10557 11851 10560
rect 11793 10551 11851 10557
rect 11885 10557 11897 10560
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 13814 10548 13820 10600
rect 13872 10548 13878 10600
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10588 13967 10591
rect 13998 10588 14004 10600
rect 13955 10560 14004 10588
rect 13955 10557 13967 10560
rect 13909 10551 13967 10557
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 16132 10597 16160 10628
rect 17034 10616 17040 10668
rect 17092 10616 17098 10668
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10656 19671 10659
rect 21361 10659 21419 10665
rect 21361 10656 21373 10659
rect 19659 10628 19840 10656
rect 19659 10625 19671 10628
rect 19613 10619 19671 10625
rect 15841 10591 15899 10597
rect 15841 10588 15853 10591
rect 15712 10560 15853 10588
rect 15712 10548 15718 10560
rect 15841 10557 15853 10560
rect 15887 10557 15899 10591
rect 15841 10551 15899 10557
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10588 16451 10591
rect 16577 10591 16635 10597
rect 16577 10588 16589 10591
rect 16439 10560 16589 10588
rect 16439 10557 16451 10560
rect 16393 10551 16451 10557
rect 16577 10557 16589 10560
rect 16623 10557 16635 10591
rect 16577 10551 16635 10557
rect 16669 10591 16727 10597
rect 16669 10557 16681 10591
rect 16715 10588 16727 10591
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16715 10560 16957 10588
rect 16715 10557 16727 10560
rect 16669 10551 16727 10557
rect 16945 10557 16957 10560
rect 16991 10588 17003 10591
rect 17126 10588 17132 10600
rect 16991 10560 17132 10588
rect 16991 10557 17003 10560
rect 16945 10551 17003 10557
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 18046 10548 18052 10600
rect 18104 10588 18110 10600
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 18104 10560 18705 10588
rect 18104 10548 18110 10560
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 18874 10548 18880 10600
rect 18932 10588 18938 10600
rect 19812 10597 19840 10628
rect 20640 10628 21373 10656
rect 18969 10591 19027 10597
rect 18969 10588 18981 10591
rect 18932 10560 18981 10588
rect 18932 10548 18938 10560
rect 18969 10557 18981 10560
rect 19015 10557 19027 10591
rect 18969 10551 19027 10557
rect 19245 10591 19303 10597
rect 19245 10557 19257 10591
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10557 19763 10591
rect 19705 10551 19763 10557
rect 19797 10591 19855 10597
rect 19797 10557 19809 10591
rect 19843 10557 19855 10591
rect 19797 10551 19855 10557
rect 9766 10520 9772 10532
rect 9416 10492 9772 10520
rect 9766 10480 9772 10492
rect 9824 10480 9830 10532
rect 10152 10492 11468 10520
rect 7834 10412 7840 10464
rect 7892 10412 7898 10464
rect 8018 10412 8024 10464
rect 8076 10452 8082 10464
rect 8113 10455 8171 10461
rect 8113 10452 8125 10455
rect 8076 10424 8125 10452
rect 8076 10412 8082 10424
rect 8113 10421 8125 10424
rect 8159 10421 8171 10455
rect 8113 10415 8171 10421
rect 8754 10412 8760 10464
rect 8812 10412 8818 10464
rect 9030 10412 9036 10464
rect 9088 10412 9094 10464
rect 9306 10412 9312 10464
rect 9364 10412 9370 10464
rect 9858 10412 9864 10464
rect 9916 10412 9922 10464
rect 10152 10461 10180 10492
rect 10137 10455 10195 10461
rect 10137 10421 10149 10455
rect 10183 10421 10195 10455
rect 10137 10415 10195 10421
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 10413 10455 10471 10461
rect 10413 10452 10425 10455
rect 10284 10424 10425 10452
rect 10284 10412 10290 10424
rect 10413 10421 10425 10424
rect 10459 10421 10471 10455
rect 11440 10452 11468 10492
rect 11514 10480 11520 10532
rect 11572 10529 11578 10532
rect 11572 10520 11584 10529
rect 12130 10523 12188 10529
rect 12130 10520 12142 10523
rect 11572 10492 11617 10520
rect 11716 10492 12142 10520
rect 11572 10483 11584 10492
rect 11572 10480 11578 10483
rect 11716 10452 11744 10492
rect 12130 10489 12142 10492
rect 12176 10489 12188 10523
rect 12130 10483 12188 10489
rect 13354 10480 13360 10532
rect 13412 10520 13418 10532
rect 14154 10523 14212 10529
rect 14154 10520 14166 10523
rect 13412 10492 14166 10520
rect 13412 10480 13418 10492
rect 14154 10489 14166 10492
rect 14200 10489 14212 10523
rect 14154 10483 14212 10489
rect 15102 10480 15108 10532
rect 15160 10520 15166 10532
rect 17304 10523 17362 10529
rect 15160 10492 16344 10520
rect 15160 10480 15166 10492
rect 11440 10424 11744 10452
rect 10413 10415 10471 10421
rect 13722 10412 13728 10464
rect 13780 10412 13786 10464
rect 15749 10455 15807 10461
rect 15749 10421 15761 10455
rect 15795 10452 15807 10455
rect 16206 10452 16212 10464
rect 15795 10424 16212 10452
rect 15795 10421 15807 10424
rect 15749 10415 15807 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16316 10461 16344 10492
rect 17304 10489 17316 10523
rect 17350 10520 17362 10523
rect 19061 10523 19119 10529
rect 19061 10520 19073 10523
rect 17350 10492 19073 10520
rect 17350 10489 17362 10492
rect 17304 10483 17362 10489
rect 19061 10489 19073 10492
rect 19107 10489 19119 10523
rect 19061 10483 19119 10489
rect 16301 10455 16359 10461
rect 16301 10421 16313 10455
rect 16347 10452 16359 10455
rect 16666 10452 16672 10464
rect 16347 10424 16672 10452
rect 16347 10421 16359 10424
rect 16301 10415 16359 10421
rect 16666 10412 16672 10424
rect 16724 10452 16730 10464
rect 17126 10452 17132 10464
rect 16724 10424 17132 10452
rect 16724 10412 16730 10424
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 18785 10455 18843 10461
rect 18785 10452 18797 10455
rect 18196 10424 18797 10452
rect 18196 10412 18202 10424
rect 18785 10421 18797 10424
rect 18831 10452 18843 10455
rect 19260 10452 19288 10551
rect 19720 10520 19748 10551
rect 20254 10548 20260 10600
rect 20312 10548 20318 10600
rect 20346 10548 20352 10600
rect 20404 10548 20410 10600
rect 20640 10597 20668 10628
rect 21361 10625 21373 10628
rect 21407 10625 21419 10659
rect 21361 10619 21419 10625
rect 20441 10591 20499 10597
rect 20441 10557 20453 10591
rect 20487 10557 20499 10591
rect 20441 10551 20499 10557
rect 20625 10591 20683 10597
rect 20625 10557 20637 10591
rect 20671 10557 20683 10591
rect 20625 10551 20683 10557
rect 20272 10520 20300 10548
rect 19720 10492 20300 10520
rect 18831 10424 19288 10452
rect 18831 10421 18843 10424
rect 18785 10415 18843 10421
rect 19886 10412 19892 10464
rect 19944 10412 19950 10464
rect 20456 10452 20484 10551
rect 20714 10548 20720 10600
rect 20772 10548 20778 10600
rect 21174 10548 21180 10600
rect 21232 10548 21238 10600
rect 21453 10591 21511 10597
rect 21453 10557 21465 10591
rect 21499 10557 21511 10591
rect 21453 10551 21511 10557
rect 20533 10523 20591 10529
rect 20533 10489 20545 10523
rect 20579 10520 20591 10523
rect 21085 10523 21143 10529
rect 21085 10520 21097 10523
rect 20579 10492 21097 10520
rect 20579 10489 20591 10492
rect 20533 10483 20591 10489
rect 21085 10489 21097 10492
rect 21131 10489 21143 10523
rect 21085 10483 21143 10489
rect 21358 10480 21364 10532
rect 21416 10520 21422 10532
rect 21468 10520 21496 10551
rect 21542 10548 21548 10600
rect 21600 10588 21606 10600
rect 21729 10591 21787 10597
rect 21729 10588 21741 10591
rect 21600 10560 21741 10588
rect 21600 10548 21606 10560
rect 21729 10557 21741 10560
rect 21775 10557 21787 10591
rect 21729 10551 21787 10557
rect 21821 10591 21879 10597
rect 21821 10557 21833 10591
rect 21867 10588 21879 10591
rect 21928 10588 21956 10696
rect 23569 10693 23581 10727
rect 23615 10724 23627 10727
rect 28258 10724 28264 10736
rect 23615 10696 28264 10724
rect 23615 10693 23627 10696
rect 23569 10687 23627 10693
rect 28258 10684 28264 10696
rect 28316 10684 28322 10736
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 23216 10628 23949 10656
rect 21867 10560 21956 10588
rect 21867 10557 21879 10560
rect 21821 10551 21879 10557
rect 21416 10492 21496 10520
rect 21744 10520 21772 10551
rect 22094 10548 22100 10600
rect 22152 10588 22158 10600
rect 22189 10591 22247 10597
rect 22189 10588 22201 10591
rect 22152 10560 22201 10588
rect 22152 10548 22158 10560
rect 22189 10557 22201 10560
rect 22235 10557 22247 10591
rect 23216 10588 23244 10628
rect 23937 10625 23949 10628
rect 23983 10656 23995 10659
rect 23983 10628 24440 10656
rect 23983 10625 23995 10628
rect 23937 10619 23995 10625
rect 22189 10551 22247 10557
rect 22287 10560 23244 10588
rect 21910 10520 21916 10532
rect 21744 10492 21916 10520
rect 21416 10480 21422 10492
rect 21910 10480 21916 10492
rect 21968 10520 21974 10532
rect 22287 10520 22315 10560
rect 23474 10548 23480 10600
rect 23532 10588 23538 10600
rect 23845 10591 23903 10597
rect 23845 10588 23857 10591
rect 23532 10560 23857 10588
rect 23532 10548 23538 10560
rect 23845 10557 23857 10560
rect 23891 10557 23903 10591
rect 23845 10551 23903 10557
rect 24302 10548 24308 10600
rect 24360 10548 24366 10600
rect 24412 10597 24440 10628
rect 24486 10616 24492 10668
rect 24544 10656 24550 10668
rect 24544 10628 25452 10656
rect 24544 10616 24550 10628
rect 24397 10591 24455 10597
rect 24397 10557 24409 10591
rect 24443 10557 24455 10591
rect 24397 10551 24455 10557
rect 24578 10548 24584 10600
rect 24636 10588 24642 10600
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 24636 10560 24685 10588
rect 24636 10548 24642 10560
rect 24673 10557 24685 10560
rect 24719 10557 24731 10591
rect 24673 10551 24731 10557
rect 25133 10591 25191 10597
rect 25133 10557 25145 10591
rect 25179 10588 25191 10591
rect 25314 10588 25320 10600
rect 25179 10560 25320 10588
rect 25179 10557 25191 10560
rect 25133 10551 25191 10557
rect 25314 10548 25320 10560
rect 25372 10548 25378 10600
rect 25424 10597 25452 10628
rect 25409 10591 25467 10597
rect 25409 10557 25421 10591
rect 25455 10588 25467 10591
rect 25593 10591 25651 10597
rect 25593 10588 25605 10591
rect 25455 10560 25605 10588
rect 25455 10557 25467 10560
rect 25409 10551 25467 10557
rect 25593 10557 25605 10560
rect 25639 10557 25651 10591
rect 25593 10551 25651 10557
rect 25682 10548 25688 10600
rect 25740 10548 25746 10600
rect 21968 10492 22315 10520
rect 22456 10523 22514 10529
rect 21968 10480 21974 10492
rect 22456 10489 22468 10523
rect 22502 10520 22514 10523
rect 25041 10523 25099 10529
rect 25041 10520 25053 10523
rect 22502 10492 25053 10520
rect 22502 10489 22514 10492
rect 22456 10483 22514 10489
rect 25041 10489 25053 10492
rect 25087 10489 25099 10523
rect 25041 10483 25099 10489
rect 20809 10455 20867 10461
rect 20809 10452 20821 10455
rect 20456 10424 20821 10452
rect 20809 10421 20821 10424
rect 20855 10421 20867 10455
rect 20809 10415 20867 10421
rect 21266 10412 21272 10464
rect 21324 10452 21330 10464
rect 21637 10455 21695 10461
rect 21637 10452 21649 10455
rect 21324 10424 21649 10452
rect 21324 10412 21330 10424
rect 21637 10421 21649 10424
rect 21683 10421 21695 10455
rect 21637 10415 21695 10421
rect 23566 10412 23572 10464
rect 23624 10452 23630 10464
rect 24026 10452 24032 10464
rect 23624 10424 24032 10452
rect 23624 10412 23630 10424
rect 24026 10412 24032 10424
rect 24084 10412 24090 10464
rect 24210 10412 24216 10464
rect 24268 10452 24274 10464
rect 31662 10452 31668 10464
rect 24268 10424 31668 10452
rect 24268 10412 24274 10424
rect 31662 10412 31668 10424
rect 31720 10412 31726 10464
rect 552 10362 31531 10384
rect 552 10310 8102 10362
rect 8154 10310 8166 10362
rect 8218 10310 8230 10362
rect 8282 10310 8294 10362
rect 8346 10310 8358 10362
rect 8410 10310 15807 10362
rect 15859 10310 15871 10362
rect 15923 10310 15935 10362
rect 15987 10310 15999 10362
rect 16051 10310 16063 10362
rect 16115 10310 23512 10362
rect 23564 10310 23576 10362
rect 23628 10310 23640 10362
rect 23692 10310 23704 10362
rect 23756 10310 23768 10362
rect 23820 10310 31217 10362
rect 31269 10310 31281 10362
rect 31333 10310 31345 10362
rect 31397 10310 31409 10362
rect 31461 10310 31473 10362
rect 31525 10310 31531 10362
rect 552 10288 31531 10310
rect 7926 10208 7932 10260
rect 7984 10208 7990 10260
rect 8018 10208 8024 10260
rect 8076 10208 8082 10260
rect 8570 10208 8576 10260
rect 8628 10208 8634 10260
rect 8754 10208 8760 10260
rect 8812 10208 8818 10260
rect 8849 10251 8907 10257
rect 8849 10217 8861 10251
rect 8895 10248 8907 10251
rect 9030 10248 9036 10260
rect 8895 10220 9036 10248
rect 8895 10217 8907 10220
rect 8849 10211 8907 10217
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9122 10208 9128 10260
rect 9180 10208 9186 10260
rect 9582 10208 9588 10260
rect 9640 10208 9646 10260
rect 9858 10208 9864 10260
rect 9916 10248 9922 10260
rect 11054 10248 11060 10260
rect 9916 10220 11060 10248
rect 9916 10208 9922 10220
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 12526 10208 12532 10260
rect 12584 10208 12590 10260
rect 12986 10208 12992 10260
rect 13044 10208 13050 10260
rect 13354 10208 13360 10260
rect 13412 10208 13418 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 13722 10248 13728 10260
rect 13679 10220 13728 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13872 10220 13921 10248
rect 13872 10208 13878 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 13909 10211 13967 10217
rect 15194 10208 15200 10260
rect 15252 10208 15258 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15565 10251 15623 10257
rect 15565 10248 15577 10251
rect 15344 10220 15577 10248
rect 15344 10208 15350 10220
rect 15565 10217 15577 10220
rect 15611 10217 15623 10251
rect 15565 10211 15623 10217
rect 16206 10208 16212 10260
rect 16264 10208 16270 10260
rect 16758 10208 16764 10260
rect 16816 10208 16822 10260
rect 18601 10251 18659 10257
rect 18601 10217 18613 10251
rect 18647 10248 18659 10251
rect 18690 10248 18696 10260
rect 18647 10220 18696 10248
rect 18647 10217 18659 10220
rect 18601 10211 18659 10217
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 19886 10208 19892 10260
rect 19944 10208 19950 10260
rect 20346 10208 20352 10260
rect 20404 10208 20410 10260
rect 20717 10251 20775 10257
rect 20717 10217 20729 10251
rect 20763 10248 20775 10251
rect 22005 10251 22063 10257
rect 22005 10248 22017 10251
rect 20763 10220 22017 10248
rect 20763 10217 20775 10220
rect 20717 10211 20775 10217
rect 22005 10217 22017 10220
rect 22051 10217 22063 10251
rect 22005 10211 22063 10217
rect 23845 10251 23903 10257
rect 23845 10217 23857 10251
rect 23891 10248 23903 10251
rect 28258 10248 28264 10260
rect 23891 10220 28264 10248
rect 23891 10217 23903 10220
rect 23845 10211 23903 10217
rect 28258 10208 28264 10220
rect 28316 10208 28322 10260
rect 7944 10180 7972 10208
rect 8588 10180 8616 10208
rect 7852 10152 7972 10180
rect 8036 10152 8616 10180
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10081 7067 10115
rect 7009 10075 7067 10081
rect 7024 10044 7052 10075
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7285 10115 7343 10121
rect 7285 10112 7297 10115
rect 7248 10084 7297 10112
rect 7248 10072 7254 10084
rect 7285 10081 7297 10084
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 7374 10072 7380 10124
rect 7432 10072 7438 10124
rect 7558 10072 7564 10124
rect 7616 10072 7622 10124
rect 7852 10121 7880 10152
rect 7837 10115 7895 10121
rect 7837 10081 7849 10115
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10112 7987 10115
rect 8036 10112 8064 10152
rect 7975 10084 8064 10112
rect 8113 10115 8171 10121
rect 7975 10081 7987 10084
rect 7929 10075 7987 10081
rect 8113 10081 8125 10115
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 8478 10112 8484 10124
rect 8435 10084 8484 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 8128 10044 8156 10075
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 8662 10072 8668 10124
rect 8720 10072 8726 10124
rect 8772 10121 8800 10208
rect 9600 10180 9628 10208
rect 11425 10183 11483 10189
rect 11425 10180 11437 10183
rect 8864 10152 9628 10180
rect 10796 10152 11437 10180
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10081 8815 10115
rect 8757 10075 8815 10081
rect 8864 10044 8892 10152
rect 8941 10115 8999 10121
rect 8941 10081 8953 10115
rect 8987 10112 8999 10115
rect 9306 10112 9312 10124
rect 8987 10084 9312 10112
rect 8987 10081 8999 10084
rect 8941 10075 8999 10081
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 10796 10121 10824 10152
rect 11425 10149 11437 10152
rect 11471 10149 11483 10183
rect 11425 10143 11483 10149
rect 11606 10140 11612 10192
rect 11664 10180 11670 10192
rect 13004 10180 13032 10208
rect 15212 10180 15240 10208
rect 16224 10180 16252 10208
rect 19052 10183 19110 10189
rect 11664 10152 12480 10180
rect 13004 10152 13308 10180
rect 11664 10140 11670 10152
rect 10238 10115 10296 10121
rect 10238 10112 10250 10115
rect 9416 10084 10250 10112
rect 7024 10016 7328 10044
rect 8128 10016 8892 10044
rect 6730 9936 6736 9988
rect 6788 9976 6794 9988
rect 7193 9979 7251 9985
rect 7193 9976 7205 9979
rect 6788 9948 7205 9976
rect 6788 9936 6794 9948
rect 7193 9945 7205 9948
rect 7239 9945 7251 9979
rect 7193 9939 7251 9945
rect 7300 9920 7328 10016
rect 7834 9936 7840 9988
rect 7892 9976 7898 9988
rect 9416 9976 9444 10084
rect 10238 10081 10250 10084
rect 10284 10081 10296 10115
rect 10238 10075 10296 10081
rect 10781 10115 10839 10121
rect 10781 10081 10793 10115
rect 10827 10081 10839 10115
rect 10781 10075 10839 10081
rect 11146 10072 11152 10124
rect 11204 10072 11210 10124
rect 11238 10072 11244 10124
rect 11296 10072 11302 10124
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 11698 10112 11704 10124
rect 11563 10084 11704 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 12069 10115 12127 10121
rect 12069 10081 12081 10115
rect 12115 10112 12127 10115
rect 12161 10115 12219 10121
rect 12161 10112 12173 10115
rect 12115 10084 12173 10112
rect 12115 10081 12127 10084
rect 12069 10075 12127 10081
rect 12161 10081 12173 10084
rect 12207 10112 12219 10115
rect 12342 10112 12348 10124
rect 12207 10084 12348 10112
rect 12207 10081 12219 10084
rect 12161 10075 12219 10081
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10044 10563 10047
rect 11164 10044 11192 10072
rect 10551 10016 11192 10044
rect 11808 10044 11836 10075
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12452 10121 12480 10152
rect 13280 10121 13308 10152
rect 13372 10152 13952 10180
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10081 12495 10115
rect 12437 10075 12495 10081
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10112 12955 10115
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 12943 10084 13185 10112
rect 12943 10081 12955 10084
rect 12897 10075 12955 10081
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 13078 10044 13084 10056
rect 11808 10016 13084 10044
rect 10551 10013 10563 10016
rect 10505 10007 10563 10013
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 13188 10044 13216 10075
rect 13372 10044 13400 10152
rect 13924 10124 13952 10152
rect 14016 10152 14688 10180
rect 15212 10152 16160 10180
rect 16224 10152 16436 10180
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10081 13783 10115
rect 13725 10075 13783 10081
rect 13188 10016 13400 10044
rect 13740 10044 13768 10075
rect 13906 10072 13912 10124
rect 13964 10072 13970 10124
rect 14016 10121 14044 10152
rect 14660 10124 14688 10152
rect 14001 10115 14059 10121
rect 14001 10081 14013 10115
rect 14047 10081 14059 10115
rect 14001 10075 14059 10081
rect 14090 10072 14096 10124
rect 14148 10072 14154 10124
rect 14366 10072 14372 10124
rect 14424 10072 14430 10124
rect 14642 10072 14648 10124
rect 14700 10072 14706 10124
rect 14829 10115 14887 10121
rect 14829 10081 14841 10115
rect 14875 10112 14887 10115
rect 14921 10115 14979 10121
rect 14921 10112 14933 10115
rect 14875 10084 14933 10112
rect 14875 10081 14887 10084
rect 14829 10075 14887 10081
rect 14921 10081 14933 10084
rect 14967 10112 14979 10115
rect 15102 10112 15108 10124
rect 14967 10084 15108 10112
rect 14967 10081 14979 10084
rect 14921 10075 14979 10081
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15197 10115 15255 10121
rect 15197 10081 15209 10115
rect 15243 10081 15255 10115
rect 15197 10075 15255 10081
rect 14185 10047 14243 10053
rect 14185 10044 14197 10047
rect 13740 10016 14197 10044
rect 14185 10013 14197 10016
rect 14231 10013 14243 10047
rect 14185 10007 14243 10013
rect 15010 10004 15016 10056
rect 15068 10044 15074 10056
rect 15212 10044 15240 10075
rect 15562 10072 15568 10124
rect 15620 10102 15626 10124
rect 15657 10115 15715 10121
rect 15657 10102 15669 10115
rect 15620 10081 15669 10102
rect 15703 10081 15715 10115
rect 15620 10075 15715 10081
rect 15749 10115 15807 10121
rect 15749 10081 15761 10115
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 15620 10074 15700 10075
rect 15620 10072 15626 10074
rect 15764 10044 15792 10075
rect 15068 10016 15240 10044
rect 15672 10016 15792 10044
rect 15068 10004 15074 10016
rect 7892 9948 9444 9976
rect 12805 9979 12863 9985
rect 7892 9936 7898 9948
rect 12805 9945 12817 9979
rect 12851 9976 12863 9979
rect 13814 9976 13820 9988
rect 12851 9948 13820 9976
rect 12851 9945 12863 9948
rect 12805 9939 12863 9945
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 15672 9976 15700 10016
rect 15838 10004 15844 10056
rect 15896 10004 15902 10056
rect 16132 10044 16160 10152
rect 16298 10072 16304 10124
rect 16356 10072 16362 10124
rect 16408 10121 16436 10152
rect 17052 10152 18828 10180
rect 17052 10124 17080 10152
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10081 16451 10115
rect 16393 10075 16451 10081
rect 16669 10115 16727 10121
rect 16669 10081 16681 10115
rect 16715 10081 16727 10115
rect 16669 10075 16727 10081
rect 16684 10044 16712 10075
rect 17034 10072 17040 10124
rect 17092 10072 17098 10124
rect 17126 10072 17132 10124
rect 17184 10112 17190 10124
rect 17310 10112 17316 10124
rect 17184 10084 17316 10112
rect 17184 10072 17190 10084
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 17488 10115 17546 10121
rect 17488 10081 17500 10115
rect 17534 10112 17546 10115
rect 18598 10112 18604 10124
rect 17534 10084 18604 10112
rect 17534 10081 17546 10084
rect 17488 10075 17546 10081
rect 18598 10072 18604 10084
rect 18656 10072 18662 10124
rect 18800 10121 18828 10152
rect 19052 10149 19064 10183
rect 19098 10180 19110 10183
rect 19904 10180 19932 10208
rect 19098 10152 19932 10180
rect 19098 10149 19110 10152
rect 19052 10143 19110 10149
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10081 18843 10115
rect 18785 10075 18843 10081
rect 16132 10016 16712 10044
rect 17052 10044 17080 10072
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 17052 10016 17233 10044
rect 17221 10013 17233 10016
rect 17267 10013 17279 10047
rect 17221 10007 17279 10013
rect 15028 9948 15700 9976
rect 6638 9868 6644 9920
rect 6696 9908 6702 9920
rect 6917 9911 6975 9917
rect 6917 9908 6929 9911
rect 6696 9880 6929 9908
rect 6696 9868 6702 9880
rect 6917 9877 6929 9880
rect 6963 9877 6975 9911
rect 6917 9871 6975 9877
rect 7282 9868 7288 9920
rect 7340 9868 7346 9920
rect 7466 9868 7472 9920
rect 7524 9868 7530 9920
rect 7742 9868 7748 9920
rect 7800 9868 7806 9920
rect 8294 9868 8300 9920
rect 8352 9868 8358 9920
rect 8570 9868 8576 9920
rect 8628 9868 8634 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 9858 9908 9864 9920
rect 8720 9880 9864 9908
rect 8720 9868 8726 9880
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 10318 9868 10324 9920
rect 10376 9908 10382 9920
rect 10689 9911 10747 9917
rect 10689 9908 10701 9911
rect 10376 9880 10701 9908
rect 10376 9868 10382 9880
rect 10689 9877 10701 9880
rect 10735 9877 10747 9911
rect 10689 9871 10747 9877
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 11149 9911 11207 9917
rect 11149 9908 11161 9911
rect 11112 9880 11161 9908
rect 11112 9868 11118 9880
rect 11149 9877 11161 9880
rect 11195 9877 11207 9911
rect 11149 9871 11207 9877
rect 11698 9868 11704 9920
rect 11756 9868 11762 9920
rect 11790 9868 11796 9920
rect 11848 9908 11854 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11848 9880 11989 9908
rect 11848 9868 11854 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 11977 9871 12035 9877
rect 12253 9911 12311 9917
rect 12253 9877 12265 9911
rect 12299 9908 12311 9911
rect 12894 9908 12900 9920
rect 12299 9880 12900 9908
rect 12299 9877 12311 9880
rect 12253 9871 12311 9877
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 12986 9868 12992 9920
rect 13044 9908 13050 9920
rect 13081 9911 13139 9917
rect 13081 9908 13093 9911
rect 13044 9880 13093 9908
rect 13044 9868 13050 9880
rect 13081 9877 13093 9880
rect 13127 9877 13139 9911
rect 13081 9871 13139 9877
rect 13906 9868 13912 9920
rect 13964 9908 13970 9920
rect 14461 9911 14519 9917
rect 14461 9908 14473 9911
rect 13964 9880 14473 9908
rect 13964 9868 13970 9880
rect 14461 9877 14473 9880
rect 14507 9877 14519 9911
rect 14461 9871 14519 9877
rect 14734 9868 14740 9920
rect 14792 9868 14798 9920
rect 15028 9917 15056 9948
rect 15746 9936 15752 9988
rect 15804 9976 15810 9988
rect 17037 9979 17095 9985
rect 17037 9976 17049 9979
rect 15804 9948 17049 9976
rect 15804 9936 15810 9948
rect 17037 9945 17049 9948
rect 17083 9945 17095 9979
rect 17037 9939 17095 9945
rect 15013 9911 15071 9917
rect 15013 9877 15025 9911
rect 15059 9877 15071 9911
rect 15013 9871 15071 9877
rect 15286 9868 15292 9920
rect 15344 9868 15350 9920
rect 15378 9868 15384 9920
rect 15436 9908 15442 9920
rect 16209 9911 16267 9917
rect 16209 9908 16221 9911
rect 15436 9880 16221 9908
rect 15436 9868 15442 9880
rect 16209 9877 16221 9880
rect 16255 9877 16267 9911
rect 16209 9871 16267 9877
rect 16482 9868 16488 9920
rect 16540 9868 16546 9920
rect 20162 9868 20168 9920
rect 20220 9868 20226 9920
rect 20364 9908 20392 10208
rect 20898 10140 20904 10192
rect 20956 10140 20962 10192
rect 21266 10140 21272 10192
rect 21324 10140 21330 10192
rect 21744 10152 22416 10180
rect 20533 10115 20591 10121
rect 20533 10081 20545 10115
rect 20579 10081 20591 10115
rect 20533 10075 20591 10081
rect 20717 10115 20775 10121
rect 20717 10081 20729 10115
rect 20763 10081 20775 10115
rect 20717 10075 20775 10081
rect 20993 10115 21051 10121
rect 20993 10081 21005 10115
rect 21039 10112 21051 10115
rect 21284 10112 21312 10140
rect 21744 10124 21772 10152
rect 21039 10084 21312 10112
rect 21039 10081 21051 10084
rect 20993 10075 21051 10081
rect 20548 9976 20576 10075
rect 20732 10044 20760 10075
rect 21358 10072 21364 10124
rect 21416 10072 21422 10124
rect 21453 10115 21511 10121
rect 21453 10081 21465 10115
rect 21499 10112 21511 10115
rect 21637 10115 21695 10121
rect 21637 10112 21649 10115
rect 21499 10084 21649 10112
rect 21499 10081 21511 10084
rect 21453 10075 21511 10081
rect 21637 10081 21649 10084
rect 21683 10081 21695 10115
rect 21637 10075 21695 10081
rect 21726 10072 21732 10124
rect 21784 10072 21790 10124
rect 21910 10072 21916 10124
rect 21968 10112 21974 10124
rect 22388 10121 22416 10152
rect 23382 10140 23388 10192
rect 23440 10180 23446 10192
rect 24946 10180 24952 10192
rect 23440 10152 24348 10180
rect 23440 10140 23446 10152
rect 22097 10115 22155 10121
rect 22097 10112 22109 10115
rect 21968 10084 22109 10112
rect 21968 10072 21974 10084
rect 22097 10081 22109 10084
rect 22143 10081 22155 10115
rect 22097 10075 22155 10081
rect 22373 10115 22431 10121
rect 22373 10081 22385 10115
rect 22419 10081 22431 10115
rect 22373 10075 22431 10081
rect 22732 10115 22790 10121
rect 22732 10081 22744 10115
rect 22778 10112 22790 10115
rect 22778 10084 23980 10112
rect 22778 10081 22790 10084
rect 22732 10075 22790 10081
rect 22281 10047 22339 10053
rect 22281 10044 22293 10047
rect 20732 10016 22293 10044
rect 22281 10013 22293 10016
rect 22327 10013 22339 10047
rect 22281 10007 22339 10013
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10013 22523 10047
rect 23952 10044 23980 10084
rect 24026 10072 24032 10124
rect 24084 10072 24090 10124
rect 24320 10121 24348 10152
rect 24412 10152 24952 10180
rect 24305 10115 24363 10121
rect 24305 10081 24317 10115
rect 24351 10081 24363 10115
rect 24305 10075 24363 10081
rect 24412 10044 24440 10152
rect 24946 10140 24952 10152
rect 25004 10140 25010 10192
rect 26142 10180 26148 10192
rect 25056 10152 26148 10180
rect 25056 10124 25084 10152
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10112 24639 10115
rect 24762 10112 24768 10124
rect 24627 10084 24768 10112
rect 24627 10081 24639 10084
rect 24581 10075 24639 10081
rect 24762 10072 24768 10084
rect 24820 10072 24826 10124
rect 24857 10115 24915 10121
rect 24857 10081 24869 10115
rect 24903 10112 24915 10115
rect 25038 10112 25044 10124
rect 24903 10084 25044 10112
rect 24903 10081 24915 10084
rect 24857 10075 24915 10081
rect 25038 10072 25044 10084
rect 25096 10072 25102 10124
rect 25130 10072 25136 10124
rect 25188 10072 25194 10124
rect 25314 10072 25320 10124
rect 25372 10072 25378 10124
rect 25884 10121 25912 10152
rect 26142 10140 26148 10152
rect 26200 10140 26206 10192
rect 25593 10115 25651 10121
rect 25593 10081 25605 10115
rect 25639 10112 25651 10115
rect 25777 10115 25835 10121
rect 25777 10112 25789 10115
rect 25639 10084 25789 10112
rect 25639 10081 25651 10084
rect 25593 10075 25651 10081
rect 25777 10081 25789 10084
rect 25823 10081 25835 10115
rect 25777 10075 25835 10081
rect 25869 10115 25927 10121
rect 25869 10081 25881 10115
rect 25915 10081 25927 10115
rect 25869 10075 25927 10081
rect 25961 10115 26019 10121
rect 25961 10081 25973 10115
rect 26007 10081 26019 10115
rect 25961 10075 26019 10081
rect 25976 10044 26004 10075
rect 26050 10044 26056 10056
rect 23952 10016 24440 10044
rect 24872 10016 26056 10044
rect 22465 10007 22523 10013
rect 21729 9979 21787 9985
rect 21729 9976 21741 9979
rect 20548 9948 21741 9976
rect 21729 9945 21741 9948
rect 21775 9945 21787 9979
rect 21729 9939 21787 9945
rect 22094 9936 22100 9988
rect 22152 9976 22158 9988
rect 22480 9976 22508 10007
rect 24872 9988 24900 10016
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 22152 9948 22508 9976
rect 22152 9936 22158 9948
rect 24854 9936 24860 9988
rect 24912 9936 24918 9988
rect 24949 9979 25007 9985
rect 24949 9945 24961 9979
rect 24995 9976 25007 9979
rect 25958 9976 25964 9988
rect 24995 9948 25964 9976
rect 24995 9945 25007 9948
rect 24949 9939 25007 9945
rect 25958 9936 25964 9948
rect 26016 9936 26022 9988
rect 21358 9908 21364 9920
rect 20364 9880 21364 9908
rect 21358 9868 21364 9880
rect 21416 9908 21422 9920
rect 21910 9908 21916 9920
rect 21416 9880 21916 9908
rect 21416 9868 21422 9880
rect 21910 9868 21916 9880
rect 21968 9868 21974 9920
rect 24121 9911 24179 9917
rect 24121 9877 24133 9911
rect 24167 9908 24179 9911
rect 24302 9908 24308 9920
rect 24167 9880 24308 9908
rect 24167 9877 24179 9880
rect 24121 9871 24179 9877
rect 24302 9868 24308 9880
rect 24360 9868 24366 9920
rect 24394 9868 24400 9920
rect 24452 9868 24458 9920
rect 24670 9868 24676 9920
rect 24728 9868 24734 9920
rect 25222 9868 25228 9920
rect 25280 9868 25286 9920
rect 25498 9868 25504 9920
rect 25556 9868 25562 9920
rect 26053 9911 26111 9917
rect 26053 9877 26065 9911
rect 26099 9908 26111 9911
rect 26234 9908 26240 9920
rect 26099 9880 26240 9908
rect 26099 9877 26111 9880
rect 26053 9871 26111 9877
rect 26234 9868 26240 9880
rect 26292 9868 26298 9920
rect 552 9818 31372 9840
rect 552 9766 4250 9818
rect 4302 9766 4314 9818
rect 4366 9766 4378 9818
rect 4430 9766 4442 9818
rect 4494 9766 4506 9818
rect 4558 9766 11955 9818
rect 12007 9766 12019 9818
rect 12071 9766 12083 9818
rect 12135 9766 12147 9818
rect 12199 9766 12211 9818
rect 12263 9766 19660 9818
rect 19712 9766 19724 9818
rect 19776 9766 19788 9818
rect 19840 9766 19852 9818
rect 19904 9766 19916 9818
rect 19968 9766 27365 9818
rect 27417 9766 27429 9818
rect 27481 9766 27493 9818
rect 27545 9766 27557 9818
rect 27609 9766 27621 9818
rect 27673 9766 31372 9818
rect 552 9744 31372 9766
rect 7190 9704 7196 9716
rect 6932 9676 7196 9704
rect 6178 9596 6184 9648
rect 6236 9596 6242 9648
rect 6273 9503 6331 9509
rect 6273 9469 6285 9503
rect 6319 9469 6331 9503
rect 6273 9463 6331 9469
rect 6288 9432 6316 9463
rect 6454 9460 6460 9512
rect 6512 9460 6518 9512
rect 6549 9503 6607 9509
rect 6549 9469 6561 9503
rect 6595 9500 6607 9503
rect 6730 9500 6736 9512
rect 6595 9472 6736 9500
rect 6595 9469 6607 9472
rect 6549 9463 6607 9469
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 6932 9500 6960 9676
rect 7190 9664 7196 9676
rect 7248 9664 7254 9716
rect 7285 9707 7343 9713
rect 7285 9673 7297 9707
rect 7331 9704 7343 9707
rect 7466 9704 7472 9716
rect 7331 9676 7472 9704
rect 7331 9673 7343 9676
rect 7285 9667 7343 9673
rect 7466 9664 7472 9676
rect 7524 9664 7530 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7837 9707 7895 9713
rect 7837 9704 7849 9707
rect 7616 9676 7849 9704
rect 7616 9664 7622 9676
rect 7837 9673 7849 9676
rect 7883 9673 7895 9707
rect 9674 9704 9680 9716
rect 7837 9667 7895 9673
rect 8220 9676 9680 9704
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 7374 9636 7380 9648
rect 7055 9608 7380 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 8220 9636 8248 9676
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 11606 9704 11612 9716
rect 9824 9676 10824 9704
rect 9824 9664 9830 9676
rect 7484 9608 8248 9636
rect 7484 9568 7512 9608
rect 8294 9596 8300 9648
rect 8352 9596 8358 9648
rect 8662 9596 8668 9648
rect 8720 9596 8726 9648
rect 10686 9636 10692 9648
rect 10060 9608 10692 9636
rect 7116 9540 7512 9568
rect 7116 9512 7144 9540
rect 8213 9513 8271 9519
rect 6871 9472 6960 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 7190 9460 7196 9512
rect 7248 9500 7254 9512
rect 7300 9500 7385 9510
rect 7469 9503 7527 9509
rect 7469 9500 7481 9503
rect 7248 9482 7481 9500
rect 7248 9472 7328 9482
rect 7357 9472 7481 9482
rect 7248 9460 7254 9472
rect 7469 9469 7481 9472
rect 7515 9469 7527 9503
rect 7469 9463 7527 9469
rect 7282 9432 7288 9444
rect 6288 9404 7288 9432
rect 7282 9392 7288 9404
rect 7340 9392 7346 9444
rect 7484 9432 7512 9463
rect 7926 9460 7932 9512
rect 7984 9509 7990 9512
rect 7984 9463 7995 9509
rect 8213 9479 8225 9513
rect 8259 9510 8271 9513
rect 8312 9510 8340 9596
rect 10060 9568 10088 9608
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 10796 9645 10824 9676
rect 10980 9676 11612 9704
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9605 10839 9639
rect 10781 9599 10839 9605
rect 10980 9568 11008 9676
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 11698 9664 11704 9716
rect 11756 9664 11762 9716
rect 11790 9664 11796 9716
rect 11848 9664 11854 9716
rect 13265 9707 13323 9713
rect 13265 9704 13277 9707
rect 12820 9676 13277 9704
rect 11057 9639 11115 9645
rect 11057 9605 11069 9639
rect 11103 9636 11115 9639
rect 11330 9636 11336 9648
rect 11103 9608 11336 9636
rect 11103 9605 11115 9608
rect 11057 9599 11115 9605
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 11716 9568 11744 9664
rect 9968 9540 10088 9568
rect 10336 9540 11008 9568
rect 11164 9540 11744 9568
rect 11808 9568 11836 9664
rect 11882 9596 11888 9648
rect 11940 9596 11946 9648
rect 12342 9636 12348 9648
rect 12268 9608 12348 9636
rect 11808 9540 12020 9568
rect 8259 9482 8340 9510
rect 8259 9479 8271 9482
rect 8213 9473 8271 9479
rect 7984 9460 7990 9463
rect 8478 9460 8484 9512
rect 8536 9500 8542 9512
rect 9968 9500 9996 9540
rect 8536 9472 9168 9500
rect 8536 9460 8542 9472
rect 8018 9432 8024 9444
rect 7484 9404 8024 9432
rect 8018 9392 8024 9404
rect 8076 9392 8082 9444
rect 8113 9435 8171 9441
rect 8113 9401 8125 9435
rect 8159 9432 8171 9435
rect 8570 9432 8576 9444
rect 8159 9404 8576 9432
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 8570 9392 8576 9404
rect 8628 9392 8634 9444
rect 9140 9376 9168 9472
rect 9646 9472 9996 9500
rect 6730 9324 6736 9376
rect 6788 9324 6794 9376
rect 7561 9367 7619 9373
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 8754 9364 8760 9376
rect 7607 9336 8760 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 9646 9364 9674 9472
rect 10042 9460 10048 9512
rect 10100 9460 10106 9512
rect 10336 9509 10364 9540
rect 10888 9509 10916 9540
rect 10321 9503 10379 9509
rect 10321 9469 10333 9503
rect 10367 9469 10379 9503
rect 10321 9463 10379 9469
rect 10413 9503 10471 9509
rect 10413 9469 10425 9503
rect 10459 9469 10471 9503
rect 10413 9463 10471 9469
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9500 11023 9503
rect 11054 9500 11060 9512
rect 11011 9472 11060 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 9766 9392 9772 9444
rect 9824 9441 9830 9444
rect 9824 9432 9836 9441
rect 10428 9432 10456 9463
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 11164 9509 11192 9540
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9469 11207 9503
rect 11149 9463 11207 9469
rect 11425 9503 11483 9509
rect 11425 9469 11437 9503
rect 11471 9469 11483 9503
rect 11425 9463 11483 9469
rect 9824 9404 9869 9432
rect 10336 9404 10456 9432
rect 11440 9432 11468 9463
rect 11514 9460 11520 9512
rect 11572 9460 11578 9512
rect 11701 9503 11759 9509
rect 11701 9469 11713 9503
rect 11747 9500 11759 9503
rect 11882 9500 11888 9512
rect 11747 9472 11888 9500
rect 11747 9469 11759 9472
rect 11701 9463 11759 9469
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 11992 9509 12020 9540
rect 12268 9509 12296 9608
rect 12342 9596 12348 9608
rect 12400 9636 12406 9648
rect 12820 9636 12848 9676
rect 13265 9673 13277 9676
rect 13311 9704 13323 9707
rect 13311 9676 13492 9704
rect 13311 9673 13323 9676
rect 13265 9667 13323 9673
rect 12400 9608 12848 9636
rect 12400 9596 12406 9608
rect 12713 9571 12771 9577
rect 12713 9568 12725 9571
rect 12360 9540 12725 9568
rect 12360 9509 12388 9540
rect 12713 9537 12725 9540
rect 12759 9537 12771 9571
rect 12713 9531 12771 9537
rect 12986 9528 12992 9580
rect 13044 9528 13050 9580
rect 11977 9503 12035 9509
rect 11977 9469 11989 9503
rect 12023 9469 12035 9503
rect 11977 9463 12035 9469
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 12345 9503 12403 9509
rect 12345 9469 12357 9503
rect 12391 9469 12403 9503
rect 12345 9463 12403 9469
rect 12529 9503 12587 9509
rect 12529 9469 12541 9503
rect 12575 9500 12587 9503
rect 12618 9500 12624 9512
rect 12575 9472 12624 9500
rect 12575 9469 12587 9472
rect 12529 9463 12587 9469
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9500 12863 9503
rect 13004 9500 13032 9528
rect 12851 9472 13032 9500
rect 13081 9503 13139 9509
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 13081 9469 13093 9503
rect 13127 9500 13139 9503
rect 13280 9500 13308 9667
rect 13464 9636 13492 9676
rect 13906 9664 13912 9716
rect 13964 9664 13970 9716
rect 14185 9707 14243 9713
rect 14185 9673 14197 9707
rect 14231 9704 14243 9707
rect 14366 9704 14372 9716
rect 14231 9676 14372 9704
rect 14231 9673 14243 9676
rect 14185 9667 14243 9673
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 15289 9707 15347 9713
rect 15289 9704 15301 9707
rect 15247 9676 15301 9704
rect 15289 9673 15301 9676
rect 15335 9704 15347 9707
rect 15562 9704 15568 9716
rect 15335 9676 15568 9704
rect 15335 9673 15347 9676
rect 15289 9667 15347 9673
rect 14642 9636 14648 9648
rect 13464 9608 14648 9636
rect 14642 9596 14648 9608
rect 14700 9596 14706 9648
rect 14737 9639 14795 9645
rect 14737 9605 14749 9639
rect 14783 9605 14795 9639
rect 14737 9599 14795 9605
rect 13906 9568 13912 9580
rect 13372 9540 13912 9568
rect 13372 9509 13400 9540
rect 13906 9528 13912 9540
rect 13964 9528 13970 9580
rect 14752 9568 14780 9599
rect 14016 9540 14780 9568
rect 13127 9472 13308 9500
rect 13357 9503 13415 9509
rect 13127 9469 13139 9472
rect 13081 9463 13139 9469
rect 13357 9469 13369 9503
rect 13403 9469 13415 9503
rect 13357 9463 13415 9469
rect 13541 9503 13599 9509
rect 13541 9469 13553 9503
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 12161 9435 12219 9441
rect 12161 9432 12173 9435
rect 11440 9404 12173 9432
rect 9824 9395 9836 9404
rect 9824 9392 9830 9395
rect 10336 9376 10364 9404
rect 12161 9401 12173 9404
rect 12207 9401 12219 9435
rect 12161 9395 12219 9401
rect 12437 9435 12495 9441
rect 12437 9401 12449 9435
rect 12483 9432 12495 9435
rect 12989 9435 13047 9441
rect 12989 9432 13001 9435
rect 12483 9404 13001 9432
rect 12483 9401 12495 9404
rect 12437 9395 12495 9401
rect 12989 9401 13001 9404
rect 13035 9401 13047 9435
rect 12989 9395 13047 9401
rect 9180 9336 9674 9364
rect 9180 9324 9186 9336
rect 10226 9324 10232 9376
rect 10284 9324 10290 9376
rect 10318 9324 10324 9376
rect 10376 9324 10382 9376
rect 10502 9324 10508 9376
rect 10560 9324 10566 9376
rect 11330 9324 11336 9376
rect 11388 9324 11394 9376
rect 11698 9324 11704 9376
rect 11756 9324 11762 9376
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 13354 9364 13360 9376
rect 12952 9336 13360 9364
rect 12952 9324 12958 9336
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 13556 9364 13584 9463
rect 13722 9460 13728 9512
rect 13780 9460 13786 9512
rect 14016 9509 14044 9540
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 14148 9472 14565 9500
rect 14148 9460 14154 9472
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 13633 9435 13691 9441
rect 13633 9401 13645 9435
rect 13679 9432 13691 9435
rect 14461 9435 14519 9441
rect 14461 9432 14473 9435
rect 13679 9404 14473 9432
rect 13679 9401 13691 9404
rect 13633 9395 13691 9401
rect 14461 9401 14473 9404
rect 14507 9401 14519 9435
rect 14568 9432 14596 9463
rect 14642 9460 14648 9512
rect 14700 9460 14706 9512
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 14921 9503 14979 9509
rect 14921 9500 14933 9503
rect 14792 9472 14933 9500
rect 14792 9460 14798 9472
rect 14921 9469 14933 9472
rect 14967 9469 14979 9503
rect 15304 9500 15332 9667
rect 15562 9664 15568 9676
rect 15620 9704 15626 9716
rect 15620 9676 15976 9704
rect 15620 9664 15626 9676
rect 15841 9639 15899 9645
rect 15841 9636 15853 9639
rect 15396 9608 15853 9636
rect 15396 9509 15424 9608
rect 15841 9605 15853 9608
rect 15887 9605 15899 9639
rect 15948 9636 15976 9676
rect 20162 9664 20168 9716
rect 20220 9704 20226 9716
rect 24210 9704 24216 9716
rect 20220 9676 24216 9704
rect 20220 9664 20226 9676
rect 24210 9664 24216 9676
rect 24268 9664 24274 9716
rect 24394 9664 24400 9716
rect 24452 9704 24458 9716
rect 24489 9707 24547 9713
rect 24489 9704 24501 9707
rect 24452 9676 24501 9704
rect 24452 9664 24458 9676
rect 24489 9673 24501 9676
rect 24535 9673 24547 9707
rect 24489 9667 24547 9673
rect 24670 9664 24676 9716
rect 24728 9704 24734 9716
rect 25041 9707 25099 9713
rect 24728 9676 24992 9704
rect 24728 9664 24734 9676
rect 17497 9639 17555 9645
rect 15948 9608 17172 9636
rect 15841 9599 15899 9605
rect 15562 9528 15568 9580
rect 15620 9528 15626 9580
rect 14921 9463 14979 9469
rect 15028 9472 15332 9500
rect 15381 9503 15439 9509
rect 15028 9432 15056 9472
rect 15381 9469 15393 9503
rect 15427 9469 15439 9503
rect 15381 9463 15439 9469
rect 15657 9503 15715 9509
rect 15657 9469 15669 9503
rect 15703 9500 15715 9503
rect 15746 9500 15752 9512
rect 15703 9472 15752 9500
rect 15703 9469 15715 9472
rect 15657 9463 15715 9469
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 15930 9460 15936 9512
rect 15988 9500 15994 9512
rect 15988 9472 16896 9500
rect 15988 9460 15994 9472
rect 14568 9404 15056 9432
rect 14461 9395 14519 9401
rect 15194 9392 15200 9444
rect 15252 9432 15258 9444
rect 16025 9435 16083 9441
rect 16025 9432 16037 9435
rect 15252 9404 16037 9432
rect 15252 9392 15258 9404
rect 16025 9401 16037 9404
rect 16071 9401 16083 9435
rect 16868 9432 16896 9472
rect 16942 9432 16948 9444
rect 16868 9404 16948 9432
rect 16025 9395 16083 9401
rect 16942 9392 16948 9404
rect 17000 9392 17006 9444
rect 17144 9432 17172 9608
rect 17497 9605 17509 9639
rect 17543 9636 17555 9639
rect 17586 9636 17592 9648
rect 17543 9608 17592 9636
rect 17543 9605 17555 9608
rect 17497 9599 17555 9605
rect 17586 9596 17592 9608
rect 17644 9596 17650 9648
rect 17954 9596 17960 9648
rect 18012 9596 18018 9648
rect 20901 9639 20959 9645
rect 20901 9605 20913 9639
rect 20947 9636 20959 9639
rect 20947 9608 21772 9636
rect 20947 9605 20959 9608
rect 20901 9599 20959 9605
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 18693 9571 18751 9577
rect 18693 9568 18705 9571
rect 17920 9540 18705 9568
rect 17920 9528 17926 9540
rect 18693 9537 18705 9540
rect 18739 9537 18751 9571
rect 18693 9531 18751 9537
rect 21744 9512 21772 9608
rect 23290 9596 23296 9648
rect 23348 9636 23354 9648
rect 23385 9639 23443 9645
rect 23385 9636 23397 9639
rect 23348 9608 23397 9636
rect 23348 9596 23354 9608
rect 23385 9605 23397 9608
rect 23431 9605 23443 9639
rect 23385 9599 23443 9605
rect 24765 9639 24823 9645
rect 24765 9605 24777 9639
rect 24811 9605 24823 9639
rect 24964 9636 24992 9676
rect 25041 9673 25053 9707
rect 25087 9704 25099 9707
rect 25130 9704 25136 9716
rect 25087 9676 25136 9704
rect 25087 9673 25099 9676
rect 25041 9667 25099 9673
rect 25130 9664 25136 9676
rect 25188 9664 25194 9716
rect 25314 9664 25320 9716
rect 25372 9704 25378 9716
rect 25593 9707 25651 9713
rect 25593 9704 25605 9707
rect 25372 9676 25605 9704
rect 25372 9664 25378 9676
rect 25593 9673 25605 9676
rect 25639 9673 25651 9707
rect 25593 9667 25651 9673
rect 25682 9664 25688 9716
rect 25740 9704 25746 9716
rect 26697 9707 26755 9713
rect 26697 9704 26709 9707
rect 25740 9676 26709 9704
rect 25740 9664 25746 9676
rect 26697 9673 26709 9676
rect 26743 9673 26755 9707
rect 26697 9667 26755 9673
rect 24964 9608 25544 9636
rect 24765 9599 24823 9605
rect 24780 9568 24808 9599
rect 23768 9540 24523 9568
rect 24780 9540 25268 9568
rect 18046 9460 18052 9512
rect 18104 9460 18110 9512
rect 18141 9503 18199 9509
rect 18141 9469 18153 9503
rect 18187 9469 18199 9503
rect 18141 9463 18199 9469
rect 18156 9432 18184 9463
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 18949 9503 19007 9509
rect 18949 9500 18961 9503
rect 18288 9472 18961 9500
rect 18288 9460 18294 9472
rect 18949 9469 18961 9472
rect 18995 9469 19007 9503
rect 18949 9463 19007 9469
rect 19426 9460 19432 9512
rect 19484 9500 19490 9512
rect 20349 9503 20407 9509
rect 20349 9500 20361 9503
rect 19484 9472 20361 9500
rect 19484 9460 19490 9472
rect 20349 9469 20361 9472
rect 20395 9469 20407 9503
rect 20349 9463 20407 9469
rect 20441 9503 20499 9509
rect 20441 9469 20453 9503
rect 20487 9500 20499 9503
rect 20533 9503 20591 9509
rect 20533 9500 20545 9503
rect 20487 9472 20545 9500
rect 20487 9469 20499 9472
rect 20441 9463 20499 9469
rect 20533 9469 20545 9472
rect 20579 9469 20591 9503
rect 20533 9463 20591 9469
rect 20625 9503 20683 9509
rect 20625 9469 20637 9503
rect 20671 9500 20683 9503
rect 20809 9503 20867 9509
rect 20809 9500 20821 9503
rect 20671 9472 20821 9500
rect 20671 9469 20683 9472
rect 20625 9463 20683 9469
rect 20809 9469 20821 9472
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 17144 9404 18184 9432
rect 20548 9432 20576 9463
rect 21358 9460 21364 9512
rect 21416 9460 21422 9512
rect 21634 9460 21640 9512
rect 21692 9460 21698 9512
rect 21726 9460 21732 9512
rect 21784 9460 21790 9512
rect 21910 9460 21916 9512
rect 21968 9460 21974 9512
rect 22005 9503 22063 9509
rect 22005 9469 22017 9503
rect 22051 9469 22063 9503
rect 22005 9463 22063 9469
rect 22272 9503 22330 9509
rect 22272 9469 22284 9503
rect 22318 9500 22330 9503
rect 23768 9500 23796 9540
rect 22318 9472 23796 9500
rect 22318 9469 22330 9472
rect 22272 9463 22330 9469
rect 20548 9404 20760 9432
rect 20732 9376 20760 9404
rect 21082 9392 21088 9444
rect 21140 9432 21146 9444
rect 21821 9435 21879 9441
rect 21821 9432 21833 9435
rect 21140 9404 21833 9432
rect 21140 9392 21146 9404
rect 21821 9401 21833 9404
rect 21867 9401 21879 9435
rect 21821 9395 21879 9401
rect 15013 9367 15071 9373
rect 15013 9364 15025 9367
rect 13556 9336 15025 9364
rect 15013 9333 15025 9336
rect 15059 9333 15071 9367
rect 15013 9327 15071 9333
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 18233 9367 18291 9373
rect 18233 9364 18245 9367
rect 15620 9336 18245 9364
rect 15620 9324 15626 9336
rect 18233 9333 18245 9336
rect 18279 9333 18291 9367
rect 18233 9327 18291 9333
rect 20070 9324 20076 9376
rect 20128 9324 20134 9376
rect 20714 9324 20720 9376
rect 20772 9324 20778 9376
rect 21266 9324 21272 9376
rect 21324 9324 21330 9376
rect 21542 9324 21548 9376
rect 21600 9324 21606 9376
rect 21928 9364 21956 9460
rect 22020 9432 22048 9463
rect 23842 9460 23848 9512
rect 23900 9460 23906 9512
rect 24121 9503 24179 9509
rect 24121 9469 24133 9503
rect 24167 9469 24179 9503
rect 24121 9463 24179 9469
rect 22094 9432 22100 9444
rect 22020 9404 22100 9432
rect 22094 9392 22100 9404
rect 22152 9392 22158 9444
rect 22186 9392 22192 9444
rect 22244 9432 22250 9444
rect 24136 9432 24164 9463
rect 24302 9460 24308 9512
rect 24360 9500 24366 9512
rect 24397 9503 24455 9509
rect 24397 9500 24409 9503
rect 24360 9472 24409 9500
rect 24360 9460 24366 9472
rect 24397 9469 24409 9472
rect 24443 9469 24455 9503
rect 24397 9463 24455 9469
rect 22244 9404 24164 9432
rect 22244 9392 22250 9404
rect 23934 9364 23940 9376
rect 21928 9336 23940 9364
rect 23934 9324 23940 9336
rect 23992 9324 23998 9376
rect 24026 9324 24032 9376
rect 24084 9364 24090 9376
rect 24213 9367 24271 9373
rect 24213 9364 24225 9367
rect 24084 9336 24225 9364
rect 24084 9324 24090 9336
rect 24213 9333 24225 9336
rect 24259 9333 24271 9367
rect 24495 9364 24523 9540
rect 24578 9460 24584 9512
rect 24636 9500 24642 9512
rect 25240 9509 25268 9540
rect 24673 9503 24731 9509
rect 24673 9500 24685 9503
rect 24636 9472 24685 9500
rect 24636 9460 24642 9472
rect 24673 9469 24685 9472
rect 24719 9469 24731 9503
rect 24949 9503 25007 9509
rect 24949 9500 24961 9503
rect 24673 9463 24731 9469
rect 24780 9472 24961 9500
rect 24780 9444 24808 9472
rect 24949 9469 24961 9472
rect 24995 9469 25007 9503
rect 24949 9463 25007 9469
rect 25225 9503 25283 9509
rect 25225 9469 25237 9503
rect 25271 9469 25283 9503
rect 25225 9463 25283 9469
rect 25314 9460 25320 9512
rect 25372 9460 25378 9512
rect 25516 9509 25544 9608
rect 26050 9596 26056 9648
rect 26108 9596 26114 9648
rect 26142 9596 26148 9648
rect 26200 9596 26206 9648
rect 25501 9503 25559 9509
rect 25501 9469 25513 9503
rect 25547 9469 25559 9503
rect 25777 9503 25835 9509
rect 25777 9500 25789 9503
rect 25501 9463 25559 9469
rect 25608 9472 25789 9500
rect 24762 9392 24768 9444
rect 24820 9432 24826 9444
rect 25608 9432 25636 9472
rect 25777 9469 25789 9472
rect 25823 9469 25835 9503
rect 25777 9463 25835 9469
rect 25866 9460 25872 9512
rect 25924 9460 25930 9512
rect 26068 9509 26096 9596
rect 26160 9568 26188 9596
rect 26160 9540 26832 9568
rect 26053 9503 26111 9509
rect 26053 9469 26065 9503
rect 26099 9469 26111 9503
rect 26053 9463 26111 9469
rect 26234 9460 26240 9512
rect 26292 9500 26298 9512
rect 26804 9509 26832 9540
rect 26329 9503 26387 9509
rect 26329 9500 26341 9503
rect 26292 9472 26341 9500
rect 26292 9460 26298 9472
rect 26329 9469 26341 9472
rect 26375 9469 26387 9503
rect 26329 9463 26387 9469
rect 26789 9503 26847 9509
rect 26789 9469 26801 9503
rect 26835 9500 26847 9503
rect 26881 9503 26939 9509
rect 26881 9500 26893 9503
rect 26835 9472 26893 9500
rect 26835 9469 26847 9472
rect 26789 9463 26847 9469
rect 26881 9469 26893 9472
rect 26927 9469 26939 9503
rect 26881 9463 26939 9469
rect 24820 9404 25636 9432
rect 25884 9404 26464 9432
rect 24820 9392 24826 9404
rect 25884 9364 25912 9404
rect 24495 9336 25912 9364
rect 26145 9367 26203 9373
rect 24213 9327 24271 9333
rect 26145 9333 26157 9367
rect 26191 9364 26203 9367
rect 26234 9364 26240 9376
rect 26191 9336 26240 9364
rect 26191 9333 26203 9336
rect 26145 9327 26203 9333
rect 26234 9324 26240 9336
rect 26292 9324 26298 9376
rect 26436 9373 26464 9404
rect 26421 9367 26479 9373
rect 26421 9333 26433 9367
rect 26467 9333 26479 9367
rect 26421 9327 26479 9333
rect 26970 9324 26976 9376
rect 27028 9324 27034 9376
rect 552 9274 31531 9296
rect 552 9222 8102 9274
rect 8154 9222 8166 9274
rect 8218 9222 8230 9274
rect 8282 9222 8294 9274
rect 8346 9222 8358 9274
rect 8410 9222 15807 9274
rect 15859 9222 15871 9274
rect 15923 9222 15935 9274
rect 15987 9222 15999 9274
rect 16051 9222 16063 9274
rect 16115 9222 23512 9274
rect 23564 9222 23576 9274
rect 23628 9222 23640 9274
rect 23692 9222 23704 9274
rect 23756 9222 23768 9274
rect 23820 9222 31217 9274
rect 31269 9222 31281 9274
rect 31333 9222 31345 9274
rect 31397 9222 31409 9274
rect 31461 9222 31473 9274
rect 31525 9222 31531 9274
rect 552 9200 31531 9222
rect 6638 9120 6644 9172
rect 6696 9120 6702 9172
rect 6730 9120 6736 9172
rect 6788 9120 6794 9172
rect 7742 9120 7748 9172
rect 7800 9120 7806 9172
rect 7929 9163 7987 9169
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8386 9160 8392 9172
rect 7975 9132 8392 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 9309 9163 9367 9169
rect 9309 9160 9321 9163
rect 8649 9132 9321 9160
rect 6748 9033 6776 9120
rect 7098 9052 7104 9104
rect 7156 9052 7162 9104
rect 7760 9092 7788 9120
rect 8649 9092 8677 9132
rect 9309 9129 9321 9132
rect 9355 9129 9367 9163
rect 9309 9123 9367 9129
rect 10226 9120 10232 9172
rect 10284 9120 10290 9172
rect 10410 9120 10416 9172
rect 10468 9120 10474 9172
rect 10502 9120 10508 9172
rect 10560 9120 10566 9172
rect 10686 9120 10692 9172
rect 10744 9120 10750 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 11756 9132 13185 9160
rect 11756 9120 11762 9132
rect 13173 9129 13185 9132
rect 13219 9129 13231 9163
rect 13173 9123 13231 9129
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 13320 9132 13492 9160
rect 13320 9120 13326 9132
rect 7484 9064 7788 9092
rect 7944 9064 8677 9092
rect 6457 9027 6515 9033
rect 6457 8993 6469 9027
rect 6503 9024 6515 9027
rect 6641 9027 6699 9033
rect 6503 8996 6592 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 6564 8888 6592 8996
rect 6641 8993 6653 9027
rect 6687 8993 6699 9027
rect 6641 8987 6699 8993
rect 6733 9027 6791 9033
rect 6733 8993 6745 9027
rect 6779 8993 6791 9027
rect 7116 9024 7144 9052
rect 7484 9033 7512 9064
rect 7944 9036 7972 9064
rect 8754 9052 8760 9104
rect 8812 9052 8818 9104
rect 9861 9095 9919 9101
rect 9416 9064 9812 9092
rect 7193 9027 7251 9033
rect 7193 9024 7205 9027
rect 7116 8996 7205 9024
rect 6733 8987 6791 8993
rect 7193 8993 7205 8996
rect 7239 8993 7251 9027
rect 7193 8987 7251 8993
rect 7469 9027 7527 9033
rect 7469 8993 7481 9027
rect 7515 8993 7527 9027
rect 7469 8987 7527 8993
rect 7561 9027 7619 9033
rect 7561 8993 7573 9027
rect 7607 9024 7619 9027
rect 7837 9027 7895 9033
rect 7837 9024 7849 9027
rect 7607 8996 7849 9024
rect 7607 8993 7619 8996
rect 7561 8987 7619 8993
rect 7837 8993 7849 8996
rect 7883 8993 7895 9027
rect 7837 8987 7895 8993
rect 6656 8956 6684 8987
rect 7101 8959 7159 8965
rect 7101 8956 7113 8959
rect 6656 8928 7113 8956
rect 7101 8925 7113 8928
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 7374 8916 7380 8968
rect 7432 8956 7438 8968
rect 7576 8956 7604 8987
rect 7432 8928 7604 8956
rect 7852 8956 7880 8987
rect 7926 8984 7932 9036
rect 7984 8984 7990 9036
rect 8110 8984 8116 9036
rect 8168 8984 8174 9036
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 8220 8996 8401 9024
rect 8220 8956 8248 8996
rect 8389 8993 8401 8996
rect 8435 9024 8447 9027
rect 8570 9024 8576 9036
rect 8435 8996 8576 9024
rect 8435 8993 8447 8996
rect 8389 8987 8447 8993
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 8665 9027 8723 9033
rect 8665 8993 8677 9027
rect 8711 8993 8723 9027
rect 8772 9024 8800 9052
rect 9416 9033 9444 9064
rect 9784 9036 9812 9064
rect 9861 9061 9873 9095
rect 9907 9092 9919 9095
rect 10134 9092 10140 9104
rect 9907 9064 10140 9092
rect 9907 9061 9919 9064
rect 9861 9055 9919 9061
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 8941 9027 8999 9033
rect 8941 9024 8953 9027
rect 8772 8996 8953 9024
rect 8665 8987 8723 8993
rect 8941 8993 8953 8996
rect 8987 8993 8999 9027
rect 8941 8987 8999 8993
rect 9401 9027 9459 9033
rect 9401 8993 9413 9027
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 7852 8928 8248 8956
rect 7432 8916 7438 8928
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8680 8956 8708 8987
rect 9508 8956 9536 8987
rect 9766 8984 9772 9036
rect 9824 8984 9830 9036
rect 10244 9033 10272 9120
rect 10520 9092 10548 9120
rect 10520 9064 10640 9092
rect 9953 9027 10011 9033
rect 9953 8993 9965 9027
rect 9999 8993 10011 9027
rect 9953 8987 10011 8993
rect 10229 9027 10287 9033
rect 10229 8993 10241 9027
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 8352 8928 8708 8956
rect 8956 8928 9536 8956
rect 9968 8956 9996 8987
rect 10318 8984 10324 9036
rect 10376 9024 10382 9036
rect 10612 9033 10640 9064
rect 11882 9052 11888 9104
rect 11940 9092 11946 9104
rect 12897 9095 12955 9101
rect 12897 9092 12909 9095
rect 11940 9064 12909 9092
rect 11940 9052 11946 9064
rect 12897 9061 12909 9064
rect 12943 9061 12955 9095
rect 12897 9055 12955 9061
rect 10505 9027 10563 9033
rect 10505 9024 10517 9027
rect 10376 8996 10517 9024
rect 10376 8984 10382 8996
rect 10505 8993 10517 8996
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 8993 10655 9027
rect 10597 8987 10655 8993
rect 12710 8984 12716 9036
rect 12768 8984 12774 9036
rect 12989 9027 13047 9033
rect 12989 8993 13001 9027
rect 13035 9024 13047 9027
rect 13078 9024 13084 9036
rect 13035 8996 13084 9024
rect 13035 8993 13047 8996
rect 12989 8987 13047 8993
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 8993 13323 9027
rect 13265 8987 13323 8993
rect 10870 8956 10876 8968
rect 9968 8928 10876 8956
rect 8352 8916 8358 8928
rect 6825 8891 6883 8897
rect 6825 8888 6837 8891
rect 6564 8860 6837 8888
rect 6825 8857 6837 8860
rect 6871 8857 6883 8891
rect 6825 8851 6883 8857
rect 7653 8891 7711 8897
rect 7653 8857 7665 8891
rect 7699 8888 7711 8891
rect 8570 8888 8576 8900
rect 7699 8860 8576 8888
rect 7699 8857 7711 8860
rect 7653 8851 7711 8857
rect 8570 8848 8576 8860
rect 8628 8848 8634 8900
rect 8956 8832 8984 8928
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 11241 8891 11299 8897
rect 11241 8888 11253 8891
rect 9732 8860 11253 8888
rect 9732 8848 9738 8860
rect 11241 8857 11253 8860
rect 11287 8857 11299 8891
rect 11241 8851 11299 8857
rect 11514 8848 11520 8900
rect 11572 8888 11578 8900
rect 13280 8888 13308 8987
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 13464 8956 13492 9132
rect 13538 9120 13544 9172
rect 13596 9120 13602 9172
rect 13722 9120 13728 9172
rect 13780 9120 13786 9172
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 15013 9163 15071 9169
rect 15013 9160 15025 9163
rect 13964 9132 15025 9160
rect 13964 9120 13970 9132
rect 15013 9129 15025 9132
rect 15059 9129 15071 9163
rect 15013 9123 15071 9129
rect 15286 9120 15292 9172
rect 15344 9120 15350 9172
rect 15654 9120 15660 9172
rect 15712 9160 15718 9172
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 15712 9132 15761 9160
rect 15712 9120 15718 9132
rect 15749 9129 15761 9132
rect 15795 9129 15807 9163
rect 15749 9123 15807 9129
rect 16482 9120 16488 9172
rect 16540 9120 16546 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 17368 9132 18000 9160
rect 17368 9120 17374 9132
rect 13556 9024 13584 9120
rect 13740 9092 13768 9120
rect 15304 9092 15332 9120
rect 13740 9064 15240 9092
rect 15304 9064 15792 9092
rect 13613 9027 13671 9033
rect 13613 9024 13625 9027
rect 13556 8996 13625 9024
rect 13613 8993 13625 8996
rect 13659 8993 13671 9027
rect 13613 8987 13671 8993
rect 15102 8984 15108 9036
rect 15160 8984 15166 9036
rect 15212 9024 15240 9064
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 15212 8996 15301 9024
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 15381 9027 15439 9033
rect 15381 8993 15393 9027
rect 15427 8993 15439 9027
rect 15381 8987 15439 8993
rect 15010 8956 15016 8968
rect 13403 8928 13492 8956
rect 14476 8928 15016 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 11572 8860 12434 8888
rect 13280 8860 13400 8888
rect 11572 8848 11578 8860
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 8205 8823 8263 8829
rect 8205 8820 8217 8823
rect 8076 8792 8217 8820
rect 8076 8780 8082 8792
rect 8205 8789 8217 8792
rect 8251 8789 8263 8823
rect 8205 8783 8263 8789
rect 8478 8780 8484 8832
rect 8536 8780 8542 8832
rect 8754 8780 8760 8832
rect 8812 8780 8818 8832
rect 8938 8780 8944 8832
rect 8996 8780 9002 8832
rect 9030 8780 9036 8832
rect 9088 8780 9094 8832
rect 9582 8780 9588 8832
rect 9640 8780 9646 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 9950 8820 9956 8832
rect 9824 8792 9956 8820
rect 9824 8780 9830 8792
rect 9950 8780 9956 8792
rect 10008 8820 10014 8832
rect 10137 8823 10195 8829
rect 10137 8820 10149 8823
rect 10008 8792 10149 8820
rect 10008 8780 10014 8792
rect 10137 8789 10149 8792
rect 10183 8820 10195 8823
rect 10318 8820 10324 8832
rect 10183 8792 10324 8820
rect 10183 8789 10195 8792
rect 10137 8783 10195 8789
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 12406 8820 12434 8860
rect 13170 8820 13176 8832
rect 12406 8792 13176 8820
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13372 8820 13400 8860
rect 14476 8832 14504 8928
rect 15010 8916 15016 8928
rect 15068 8956 15074 8968
rect 15396 8956 15424 8987
rect 15562 8984 15568 9036
rect 15620 9024 15626 9036
rect 15764 9033 15792 9064
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15620 8996 15669 9024
rect 15620 8984 15626 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 15749 9027 15807 9033
rect 15749 8993 15761 9027
rect 15795 8993 15807 9027
rect 15749 8987 15807 8993
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16500 9024 16528 9120
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 17865 9095 17923 9101
rect 17865 9092 17877 9095
rect 17828 9064 17877 9092
rect 17828 9052 17834 9064
rect 17865 9061 17877 9064
rect 17911 9061 17923 9095
rect 17972 9092 18000 9132
rect 18046 9120 18052 9172
rect 18104 9120 18110 9172
rect 21082 9120 21088 9172
rect 21140 9120 21146 9172
rect 21542 9120 21548 9172
rect 21600 9120 21606 9172
rect 21913 9163 21971 9169
rect 21913 9129 21925 9163
rect 21959 9160 21971 9163
rect 22186 9160 22192 9172
rect 21959 9132 22192 9160
rect 21959 9129 21971 9132
rect 21913 9123 21971 9129
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 23842 9160 23848 9172
rect 22296 9132 23848 9160
rect 20990 9092 20996 9104
rect 17972 9064 18276 9092
rect 17865 9055 17923 9061
rect 15979 8996 16528 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16942 8984 16948 9036
rect 17000 9024 17006 9036
rect 18138 9024 18144 9036
rect 17000 8996 18144 9024
rect 17000 8984 17006 8996
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 18248 9033 18276 9064
rect 20548 9064 20996 9092
rect 20548 9033 20576 9064
rect 20990 9052 20996 9064
rect 21048 9052 21054 9104
rect 21560 9092 21588 9120
rect 21108 9064 21588 9092
rect 21637 9095 21695 9101
rect 21108 9033 21136 9064
rect 21637 9061 21649 9095
rect 21683 9092 21695 9095
rect 22296 9092 22324 9132
rect 23842 9120 23848 9132
rect 23900 9120 23906 9172
rect 23934 9120 23940 9172
rect 23992 9160 23998 9172
rect 25038 9160 25044 9172
rect 23992 9132 25044 9160
rect 23992 9120 23998 9132
rect 25038 9120 25044 9132
rect 25096 9120 25102 9172
rect 25314 9120 25320 9172
rect 25372 9120 25378 9172
rect 25866 9120 25872 9172
rect 25924 9120 25930 9172
rect 25958 9120 25964 9172
rect 26016 9120 26022 9172
rect 26970 9120 26976 9172
rect 27028 9120 27034 9172
rect 21683 9064 22324 9092
rect 21683 9061 21695 9064
rect 21637 9055 21695 9061
rect 22370 9052 22376 9104
rect 22428 9052 22434 9104
rect 23474 9052 23480 9104
rect 23532 9092 23538 9104
rect 24854 9092 24860 9104
rect 23532 9064 24860 9092
rect 23532 9052 23538 9064
rect 24854 9052 24860 9064
rect 24912 9052 24918 9104
rect 18233 9027 18291 9033
rect 18233 8993 18245 9027
rect 18279 8993 18291 9027
rect 18233 8987 18291 8993
rect 18509 9027 18567 9033
rect 18509 8993 18521 9027
rect 18555 9024 18567 9027
rect 20441 9027 20499 9033
rect 18555 8996 19334 9024
rect 18555 8993 18567 8996
rect 18509 8987 18567 8993
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 15068 8928 16129 8956
rect 15068 8916 15074 8928
rect 16117 8925 16129 8928
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 18782 8916 18788 8968
rect 18840 8916 18846 8968
rect 19306 8956 19334 8996
rect 20441 8993 20453 9027
rect 20487 9024 20499 9027
rect 20533 9027 20591 9033
rect 20533 9024 20545 9027
rect 20487 8996 20545 9024
rect 20487 8993 20499 8996
rect 20441 8987 20499 8993
rect 20533 8993 20545 8996
rect 20579 8993 20591 9027
rect 20533 8987 20591 8993
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 9024 20959 9027
rect 21085 9027 21143 9033
rect 20947 8996 21036 9024
rect 20947 8993 20959 8996
rect 20901 8987 20959 8993
rect 20806 8956 20812 8968
rect 19306 8928 20812 8956
rect 20806 8916 20812 8928
rect 20864 8916 20870 8968
rect 21008 8956 21036 8996
rect 21085 8993 21097 9027
rect 21131 8993 21143 9027
rect 21085 8987 21143 8993
rect 21266 8984 21272 9036
rect 21324 8984 21330 9036
rect 21545 9027 21603 9033
rect 21545 8993 21557 9027
rect 21591 9024 21603 9027
rect 21726 9024 21732 9036
rect 21591 8996 21732 9024
rect 21591 8993 21603 8996
rect 21545 8987 21603 8993
rect 21726 8984 21732 8996
rect 21784 8984 21790 9036
rect 21821 9027 21879 9033
rect 21821 8993 21833 9027
rect 21867 8993 21879 9027
rect 21821 8987 21879 8993
rect 22097 9027 22155 9033
rect 22097 8993 22109 9027
rect 22143 8993 22155 9027
rect 22097 8987 22155 8993
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 21008 8928 21373 8956
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21836 8956 21864 8987
rect 21910 8956 21916 8968
rect 21836 8928 21916 8956
rect 21361 8919 21419 8925
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 20254 8848 20260 8900
rect 20312 8888 20318 8900
rect 21634 8888 21640 8900
rect 20312 8860 21640 8888
rect 20312 8848 20318 8860
rect 21634 8848 21640 8860
rect 21692 8888 21698 8900
rect 22112 8888 22140 8987
rect 22186 8984 22192 9036
rect 22244 9024 22250 9036
rect 23492 9024 23520 9052
rect 22244 8996 23520 9024
rect 24480 9027 24538 9033
rect 22244 8984 22250 8996
rect 24480 8993 24492 9027
rect 24526 9024 24538 9027
rect 25332 9024 25360 9120
rect 25777 9027 25835 9033
rect 25777 9024 25789 9027
rect 24526 8996 25268 9024
rect 25332 8996 25789 9024
rect 24526 8993 24538 8996
rect 24480 8987 24538 8993
rect 22922 8916 22928 8968
rect 22980 8956 22986 8968
rect 24213 8959 24271 8965
rect 24213 8956 24225 8959
rect 22980 8928 24225 8956
rect 22980 8916 22986 8928
rect 24213 8925 24225 8928
rect 24259 8925 24271 8959
rect 25240 8956 25268 8996
rect 25777 8993 25789 8996
rect 25823 8993 25835 9027
rect 25884 9024 25912 9120
rect 25961 9027 26019 9033
rect 25961 9024 25973 9027
rect 25884 8996 25973 9024
rect 25777 8987 25835 8993
rect 25961 8993 25973 8996
rect 26007 8993 26019 9027
rect 25961 8987 26019 8993
rect 26050 8984 26056 9036
rect 26108 8984 26114 9036
rect 26513 9027 26571 9033
rect 26513 8993 26525 9027
rect 26559 8993 26571 9027
rect 26513 8987 26571 8993
rect 26605 9027 26663 9033
rect 26605 8993 26617 9027
rect 26651 9024 26663 9027
rect 26988 9024 27016 9120
rect 26651 8996 27016 9024
rect 26651 8993 26663 8996
rect 26605 8987 26663 8993
rect 26528 8956 26556 8987
rect 25240 8928 26556 8956
rect 24213 8919 24271 8925
rect 21692 8860 23888 8888
rect 21692 8848 21698 8860
rect 23860 8832 23888 8860
rect 25406 8848 25412 8900
rect 25464 8888 25470 8900
rect 26234 8888 26240 8900
rect 25464 8860 26240 8888
rect 25464 8848 25470 8860
rect 26234 8848 26240 8860
rect 26292 8848 26298 8900
rect 14090 8820 14096 8832
rect 13372 8792 14096 8820
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 14458 8780 14464 8832
rect 14516 8780 14522 8832
rect 14734 8780 14740 8832
rect 14792 8780 14798 8832
rect 15562 8780 15568 8832
rect 15620 8780 15626 8832
rect 18322 8780 18328 8832
rect 18380 8780 18386 8832
rect 20073 8823 20131 8829
rect 20073 8789 20085 8823
rect 20119 8820 20131 8823
rect 20162 8820 20168 8832
rect 20119 8792 20168 8820
rect 20119 8789 20131 8792
rect 20073 8783 20131 8789
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 20346 8780 20352 8832
rect 20404 8780 20410 8832
rect 20625 8823 20683 8829
rect 20625 8789 20637 8823
rect 20671 8820 20683 8823
rect 21174 8820 21180 8832
rect 20671 8792 21180 8820
rect 20671 8789 20683 8792
rect 20625 8783 20683 8789
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 22189 8823 22247 8829
rect 22189 8789 22201 8823
rect 22235 8820 22247 8823
rect 23014 8820 23020 8832
rect 22235 8792 23020 8820
rect 22235 8789 22247 8792
rect 22189 8783 22247 8789
rect 23014 8780 23020 8792
rect 23072 8780 23078 8832
rect 23842 8780 23848 8832
rect 23900 8820 23906 8832
rect 24578 8820 24584 8832
rect 23900 8792 24584 8820
rect 23900 8780 23906 8792
rect 24578 8780 24584 8792
rect 24636 8780 24642 8832
rect 25590 8780 25596 8832
rect 25648 8780 25654 8832
rect 25958 8780 25964 8832
rect 26016 8820 26022 8832
rect 26145 8823 26203 8829
rect 26145 8820 26157 8823
rect 26016 8792 26157 8820
rect 26016 8780 26022 8792
rect 26145 8789 26157 8792
rect 26191 8789 26203 8823
rect 26145 8783 26203 8789
rect 552 8730 31372 8752
rect 552 8678 4250 8730
rect 4302 8678 4314 8730
rect 4366 8678 4378 8730
rect 4430 8678 4442 8730
rect 4494 8678 4506 8730
rect 4558 8678 11955 8730
rect 12007 8678 12019 8730
rect 12071 8678 12083 8730
rect 12135 8678 12147 8730
rect 12199 8678 12211 8730
rect 12263 8678 19660 8730
rect 19712 8678 19724 8730
rect 19776 8678 19788 8730
rect 19840 8678 19852 8730
rect 19904 8678 19916 8730
rect 19968 8678 27365 8730
rect 27417 8678 27429 8730
rect 27481 8678 27493 8730
rect 27545 8678 27557 8730
rect 27609 8678 27621 8730
rect 27673 8678 31372 8730
rect 552 8656 31372 8678
rect 7650 8616 7656 8628
rect 7116 8588 7656 8616
rect 6730 8372 6736 8424
rect 6788 8372 6794 8424
rect 7116 8421 7144 8588
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 8113 8619 8171 8625
rect 8113 8585 8125 8619
rect 8159 8616 8171 8619
rect 8294 8616 8300 8628
rect 8159 8588 8300 8616
rect 8159 8585 8171 8588
rect 8113 8579 8171 8585
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 9030 8616 9036 8628
rect 8619 8588 9036 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10686 8616 10692 8628
rect 10100 8588 10692 8616
rect 10100 8576 10106 8588
rect 7190 8508 7196 8560
rect 7248 8508 7254 8560
rect 7285 8551 7343 8557
rect 7285 8517 7297 8551
rect 7331 8548 7343 8551
rect 7834 8548 7840 8560
rect 7331 8520 7840 8548
rect 7331 8517 7343 8520
rect 7285 8511 7343 8517
rect 7834 8508 7840 8520
rect 7892 8508 7898 8560
rect 8404 8520 8616 8548
rect 7208 8480 7236 8508
rect 7561 8483 7619 8489
rect 7208 8452 7512 8480
rect 7484 8421 7512 8452
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 8404 8480 8432 8520
rect 7607 8452 8432 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8412 6883 8415
rect 7009 8415 7067 8421
rect 7009 8412 7021 8415
rect 6871 8384 7021 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 7009 8381 7021 8384
rect 7055 8381 7067 8415
rect 7009 8375 7067 8381
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 7377 8415 7435 8421
rect 7377 8381 7389 8415
rect 7423 8381 7435 8415
rect 7377 8375 7435 8381
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 7392 8344 7420 8375
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 7745 8415 7803 8421
rect 7745 8412 7757 8415
rect 7708 8384 7757 8412
rect 7708 8372 7714 8384
rect 7745 8381 7757 8384
rect 7791 8412 7803 8415
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7791 8384 8033 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 7837 8347 7895 8353
rect 7392 8316 7788 8344
rect 7760 8288 7788 8316
rect 7837 8313 7849 8347
rect 7883 8344 7895 8347
rect 7926 8344 7932 8356
rect 7883 8316 7932 8344
rect 7883 8313 7895 8316
rect 7837 8307 7895 8313
rect 7926 8304 7932 8316
rect 7984 8304 7990 8356
rect 8036 8344 8064 8375
rect 8478 8372 8484 8424
rect 8536 8372 8542 8424
rect 8588 8412 8616 8520
rect 8662 8508 8668 8560
rect 8720 8548 8726 8560
rect 8720 8520 8800 8548
rect 8720 8508 8726 8520
rect 8662 8412 8668 8424
rect 8588 8384 8668 8412
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8772 8412 8800 8520
rect 8846 8508 8852 8560
rect 8904 8508 8910 8560
rect 10244 8489 10272 8588
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10870 8576 10876 8628
rect 10928 8576 10934 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 11195 8588 12572 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 10778 8548 10784 8560
rect 10520 8520 10784 8548
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 10410 8412 10416 8424
rect 8772 8384 10416 8412
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 10520 8421 10548 8520
rect 10778 8508 10784 8520
rect 10836 8508 10842 8560
rect 12544 8548 12572 8588
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 12676 8588 14381 8616
rect 12676 8576 12682 8588
rect 14369 8585 14381 8588
rect 14415 8585 14427 8619
rect 14369 8579 14427 8585
rect 15562 8576 15568 8628
rect 15620 8576 15626 8628
rect 16758 8616 16764 8628
rect 15948 8588 16764 8616
rect 12544 8520 12940 8548
rect 12912 8492 12940 8520
rect 13170 8508 13176 8560
rect 13228 8548 13234 8560
rect 13817 8551 13875 8557
rect 13817 8548 13829 8551
rect 13228 8520 13829 8548
rect 13228 8508 13234 8520
rect 13817 8517 13829 8520
rect 13863 8517 13875 8551
rect 13817 8511 13875 8517
rect 14090 8508 14096 8560
rect 14148 8508 14154 8560
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8449 11667 8483
rect 11609 8443 11667 8449
rect 10505 8415 10563 8421
rect 10505 8381 10517 8415
rect 10551 8381 10563 8415
rect 10505 8375 10563 8381
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 10781 8415 10839 8421
rect 10781 8412 10793 8415
rect 10652 8384 10793 8412
rect 10652 8372 10658 8384
rect 10781 8381 10793 8384
rect 10827 8381 10839 8415
rect 10781 8375 10839 8381
rect 11057 8415 11115 8421
rect 11057 8381 11069 8415
rect 11103 8412 11115 8415
rect 11146 8412 11152 8424
rect 11103 8384 11152 8412
rect 11103 8381 11115 8384
rect 11057 8375 11115 8381
rect 11146 8372 11152 8384
rect 11204 8372 11210 8424
rect 11330 8372 11336 8424
rect 11388 8372 11394 8424
rect 11514 8372 11520 8424
rect 11572 8412 11578 8424
rect 11624 8412 11652 8443
rect 12894 8440 12900 8492
rect 12952 8440 12958 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 13280 8452 14565 8480
rect 13280 8424 13308 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 11572 8384 11652 8412
rect 11572 8372 11578 8384
rect 11698 8372 11704 8424
rect 11756 8412 11762 8424
rect 13173 8415 13231 8421
rect 13173 8412 13185 8415
rect 11756 8384 13185 8412
rect 11756 8372 11762 8384
rect 13173 8381 13185 8384
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 13262 8372 13268 8424
rect 13320 8372 13326 8424
rect 13354 8372 13360 8424
rect 13412 8412 13418 8424
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 13412 8384 13737 8412
rect 13412 8372 13418 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 13814 8372 13820 8424
rect 13872 8412 13878 8424
rect 14001 8415 14059 8421
rect 14001 8412 14013 8415
rect 13872 8384 14013 8412
rect 13872 8372 13878 8384
rect 14001 8381 14013 8384
rect 14047 8381 14059 8415
rect 14001 8375 14059 8381
rect 14458 8372 14464 8424
rect 14516 8372 14522 8424
rect 8938 8344 8944 8356
rect 8036 8316 8944 8344
rect 8938 8304 8944 8316
rect 8996 8304 9002 8356
rect 9766 8304 9772 8356
rect 9824 8344 9830 8356
rect 9962 8347 10020 8353
rect 9962 8344 9974 8347
rect 9824 8316 9974 8344
rect 9824 8304 9830 8316
rect 9962 8313 9974 8316
rect 10008 8313 10020 8347
rect 9962 8307 10020 8313
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 10192 8316 11376 8344
rect 10192 8304 10198 8316
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 8110 8276 8116 8288
rect 7800 8248 8116 8276
rect 7800 8236 7806 8248
rect 8110 8236 8116 8248
rect 8168 8276 8174 8288
rect 10042 8276 10048 8288
rect 8168 8248 10048 8276
rect 8168 8236 8174 8248
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 10594 8236 10600 8288
rect 10652 8236 10658 8288
rect 11348 8276 11376 8316
rect 11422 8304 11428 8356
rect 11480 8304 11486 8356
rect 11854 8347 11912 8353
rect 11854 8313 11866 8347
rect 11900 8313 11912 8347
rect 11854 8307 11912 8313
rect 11869 8276 11897 8307
rect 13078 8304 13084 8356
rect 13136 8344 13142 8356
rect 13906 8344 13912 8356
rect 13136 8316 13912 8344
rect 13136 8304 13142 8316
rect 13906 8304 13912 8316
rect 13964 8344 13970 8356
rect 14476 8344 14504 8372
rect 13964 8316 14504 8344
rect 14820 8347 14878 8353
rect 13964 8304 13970 8316
rect 14820 8313 14832 8347
rect 14866 8344 14878 8347
rect 15286 8344 15292 8356
rect 14866 8316 15292 8344
rect 14866 8313 14878 8316
rect 14820 8307 14878 8313
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 15580 8344 15608 8576
rect 15948 8557 15976 8588
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 17773 8619 17831 8625
rect 17773 8585 17785 8619
rect 17819 8616 17831 8619
rect 18230 8616 18236 8628
rect 17819 8588 18236 8616
rect 17819 8585 17831 8588
rect 17773 8579 17831 8585
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 18322 8576 18328 8628
rect 18380 8576 18386 8628
rect 18782 8576 18788 8628
rect 18840 8616 18846 8628
rect 19337 8619 19395 8625
rect 19337 8616 19349 8619
rect 18840 8588 19349 8616
rect 18840 8576 18846 8588
rect 19337 8585 19349 8588
rect 19383 8585 19395 8619
rect 19337 8579 19395 8585
rect 20165 8619 20223 8625
rect 20165 8585 20177 8619
rect 20211 8616 20223 8619
rect 21269 8619 21327 8625
rect 20211 8588 20852 8616
rect 20211 8585 20223 8588
rect 20165 8579 20223 8585
rect 15933 8551 15991 8557
rect 15933 8517 15945 8551
rect 15979 8517 15991 8551
rect 18340 8548 18368 8576
rect 15933 8511 15991 8517
rect 17880 8520 18368 8548
rect 16117 8415 16175 8421
rect 16117 8381 16129 8415
rect 16163 8412 16175 8415
rect 16850 8412 16856 8424
rect 16163 8384 16856 8412
rect 16163 8381 16175 8384
rect 16117 8375 16175 8381
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 17880 8421 17908 8520
rect 20346 8508 20352 8560
rect 20404 8508 20410 8560
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8480 18107 8483
rect 18095 8452 18736 8480
rect 18095 8449 18107 8452
rect 18049 8443 18107 8449
rect 17865 8415 17923 8421
rect 17865 8381 17877 8415
rect 17911 8381 17923 8415
rect 17865 8375 17923 8381
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18708 8421 18736 8452
rect 18874 8440 18880 8492
rect 18932 8480 18938 8492
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 18932 8452 19901 8480
rect 18932 8440 18938 8452
rect 19889 8449 19901 8452
rect 19935 8449 19947 8483
rect 20364 8480 20392 8508
rect 20364 8452 20760 8480
rect 19889 8443 19947 8449
rect 18417 8415 18475 8421
rect 18417 8412 18429 8415
rect 18012 8384 18429 8412
rect 18012 8372 18018 8384
rect 18417 8381 18429 8384
rect 18463 8381 18475 8415
rect 18417 8375 18475 8381
rect 18693 8415 18751 8421
rect 18693 8381 18705 8415
rect 18739 8381 18751 8415
rect 18693 8375 18751 8381
rect 18969 8415 19027 8421
rect 18969 8381 18981 8415
rect 19015 8381 19027 8415
rect 18969 8375 19027 8381
rect 16362 8347 16420 8353
rect 16362 8344 16374 8347
rect 15580 8316 16374 8344
rect 16362 8313 16374 8316
rect 16408 8313 16420 8347
rect 16362 8307 16420 8313
rect 17126 8304 17132 8356
rect 17184 8344 17190 8356
rect 18325 8347 18383 8353
rect 18325 8344 18337 8347
rect 17184 8316 18337 8344
rect 17184 8304 17190 8316
rect 18325 8313 18337 8316
rect 18371 8313 18383 8347
rect 18325 8307 18383 8313
rect 18506 8304 18512 8356
rect 18564 8344 18570 8356
rect 18785 8347 18843 8353
rect 18785 8344 18797 8347
rect 18564 8316 18797 8344
rect 18564 8304 18570 8316
rect 18785 8313 18797 8316
rect 18831 8313 18843 8347
rect 18785 8307 18843 8313
rect 11348 8248 11897 8276
rect 12986 8236 12992 8288
rect 13044 8236 13050 8288
rect 13265 8279 13323 8285
rect 13265 8245 13277 8279
rect 13311 8276 13323 8279
rect 13722 8276 13728 8288
rect 13311 8248 13728 8276
rect 13311 8245 13323 8248
rect 13265 8239 13323 8245
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 17494 8236 17500 8288
rect 17552 8236 17558 8288
rect 18984 8276 19012 8375
rect 19426 8372 19432 8424
rect 19484 8372 19490 8424
rect 19521 8415 19579 8421
rect 19521 8381 19533 8415
rect 19567 8381 19579 8415
rect 19521 8375 19579 8381
rect 19613 8415 19671 8421
rect 19613 8381 19625 8415
rect 19659 8412 19671 8415
rect 19797 8415 19855 8421
rect 19797 8412 19809 8415
rect 19659 8384 19809 8412
rect 19659 8381 19671 8384
rect 19613 8375 19671 8381
rect 19797 8381 19809 8384
rect 19843 8381 19855 8415
rect 19797 8375 19855 8381
rect 19061 8347 19119 8353
rect 19061 8313 19073 8347
rect 19107 8344 19119 8347
rect 19536 8344 19564 8375
rect 20254 8372 20260 8424
rect 20312 8372 20318 8424
rect 20530 8372 20536 8424
rect 20588 8372 20594 8424
rect 20633 8415 20691 8421
rect 20633 8381 20645 8415
rect 20679 8412 20691 8415
rect 20732 8412 20760 8452
rect 20679 8384 20760 8412
rect 20824 8412 20852 8588
rect 21269 8585 21281 8619
rect 21315 8616 21327 8619
rect 21818 8616 21824 8628
rect 21315 8588 21824 8616
rect 21315 8585 21327 8588
rect 21269 8579 21327 8585
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 24026 8616 24032 8628
rect 23216 8588 24032 8616
rect 20898 8508 20904 8560
rect 20956 8508 20962 8560
rect 22830 8508 22836 8560
rect 22888 8508 22894 8560
rect 20916 8480 20944 8508
rect 21450 8480 21456 8492
rect 20916 8452 21456 8480
rect 21450 8440 21456 8452
rect 21508 8440 21514 8492
rect 20901 8415 20959 8421
rect 20901 8412 20913 8415
rect 20824 8384 20913 8412
rect 20679 8381 20691 8384
rect 20633 8375 20691 8381
rect 20901 8381 20913 8384
rect 20947 8381 20959 8415
rect 20901 8375 20959 8381
rect 21085 8415 21143 8421
rect 21085 8381 21097 8415
rect 21131 8381 21143 8415
rect 21085 8375 21143 8381
rect 20441 8347 20499 8353
rect 19107 8316 19472 8344
rect 19536 8316 20300 8344
rect 19107 8313 19119 8316
rect 19061 8307 19119 8313
rect 19444 8288 19472 8316
rect 20272 8288 20300 8316
rect 20441 8313 20453 8347
rect 20487 8344 20499 8347
rect 20993 8347 21051 8353
rect 20993 8344 21005 8347
rect 20487 8316 21005 8344
rect 20487 8313 20499 8316
rect 20441 8307 20499 8313
rect 20993 8313 21005 8316
rect 21039 8313 21051 8347
rect 20993 8307 21051 8313
rect 19150 8276 19156 8288
rect 18984 8248 19156 8276
rect 19150 8236 19156 8248
rect 19208 8236 19214 8288
rect 19426 8236 19432 8288
rect 19484 8236 19490 8288
rect 20254 8236 20260 8288
rect 20312 8236 20318 8288
rect 20717 8279 20775 8285
rect 20717 8245 20729 8279
rect 20763 8276 20775 8279
rect 21100 8276 21128 8375
rect 21174 8372 21180 8424
rect 21232 8372 21238 8424
rect 23014 8372 23020 8424
rect 23072 8372 23078 8424
rect 23216 8421 23244 8588
rect 24026 8576 24032 8588
rect 24084 8576 24090 8628
rect 24213 8619 24271 8625
rect 24213 8585 24225 8619
rect 24259 8616 24271 8619
rect 25222 8616 25228 8628
rect 24259 8588 25228 8616
rect 24259 8585 24271 8588
rect 24213 8579 24271 8585
rect 25222 8576 25228 8588
rect 25280 8576 25286 8628
rect 25317 8619 25375 8625
rect 25317 8585 25329 8619
rect 25363 8616 25375 8619
rect 25498 8616 25504 8628
rect 25363 8588 25504 8616
rect 25363 8585 25375 8588
rect 25317 8579 25375 8585
rect 25498 8576 25504 8588
rect 25556 8576 25562 8628
rect 25682 8576 25688 8628
rect 25740 8616 25746 8628
rect 25740 8588 26740 8616
rect 25740 8576 25746 8588
rect 23382 8508 23388 8560
rect 23440 8508 23446 8560
rect 23474 8508 23480 8560
rect 23532 8508 23538 8560
rect 24504 8520 25176 8548
rect 23201 8415 23259 8421
rect 23201 8381 23213 8415
rect 23247 8381 23259 8415
rect 23201 8375 23259 8381
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 23492 8412 23520 8508
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8480 23995 8483
rect 23983 8452 24440 8480
rect 23983 8449 23995 8452
rect 23937 8443 23995 8449
rect 23339 8384 23520 8412
rect 23845 8415 23903 8421
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 23845 8381 23857 8415
rect 23891 8412 23903 8415
rect 24026 8412 24032 8424
rect 23891 8384 24032 8412
rect 23891 8381 23903 8384
rect 23845 8375 23903 8381
rect 24026 8372 24032 8384
rect 24084 8372 24090 8424
rect 24118 8372 24124 8424
rect 24176 8372 24182 8424
rect 24412 8421 24440 8452
rect 24397 8415 24455 8421
rect 24397 8381 24409 8415
rect 24443 8381 24455 8415
rect 24397 8375 24455 8381
rect 21720 8347 21778 8353
rect 21720 8313 21732 8347
rect 21766 8344 21778 8347
rect 21910 8344 21916 8356
rect 21766 8316 21916 8344
rect 21766 8313 21778 8316
rect 21720 8307 21778 8313
rect 21910 8304 21916 8316
rect 21968 8304 21974 8356
rect 24504 8353 24532 8520
rect 24578 8440 24584 8492
rect 24636 8480 24642 8492
rect 25148 8480 25176 8520
rect 26050 8508 26056 8560
rect 26108 8508 26114 8560
rect 26712 8557 26740 8588
rect 26697 8551 26755 8557
rect 26697 8517 26709 8551
rect 26743 8517 26755 8551
rect 26697 8511 26755 8517
rect 25222 8480 25228 8492
rect 24636 8452 24900 8480
rect 24636 8440 24642 8452
rect 24872 8421 24900 8452
rect 25148 8452 25228 8480
rect 25148 8421 25176 8452
rect 25222 8440 25228 8452
rect 25280 8480 25286 8492
rect 26068 8480 26096 8508
rect 25280 8452 25544 8480
rect 25280 8440 25286 8452
rect 24857 8415 24915 8421
rect 24857 8381 24869 8415
rect 24903 8381 24915 8415
rect 24857 8375 24915 8381
rect 25133 8415 25191 8421
rect 25133 8381 25145 8415
rect 25179 8381 25191 8415
rect 25133 8375 25191 8381
rect 25406 8372 25412 8424
rect 25464 8372 25470 8424
rect 25516 8412 25544 8452
rect 25700 8452 26096 8480
rect 25700 8421 25728 8452
rect 25685 8415 25743 8421
rect 25685 8412 25697 8415
rect 25516 8384 25697 8412
rect 25685 8381 25697 8384
rect 25731 8381 25743 8415
rect 25685 8375 25743 8381
rect 25777 8415 25835 8421
rect 25777 8381 25789 8415
rect 25823 8381 25835 8415
rect 25777 8375 25835 8381
rect 24489 8347 24547 8353
rect 24489 8344 24501 8347
rect 22940 8316 24501 8344
rect 20763 8248 21128 8276
rect 20763 8245 20775 8248
rect 20717 8239 20775 8245
rect 21174 8236 21180 8288
rect 21232 8276 21238 8288
rect 22940 8276 22968 8316
rect 24489 8313 24501 8316
rect 24535 8313 24547 8347
rect 24489 8307 24547 8313
rect 24578 8304 24584 8356
rect 24636 8344 24642 8356
rect 25792 8344 25820 8375
rect 25866 8372 25872 8424
rect 25924 8412 25930 8424
rect 26053 8415 26111 8421
rect 26053 8412 26065 8415
rect 25924 8384 26065 8412
rect 25924 8372 25930 8384
rect 26053 8381 26065 8384
rect 26099 8381 26111 8415
rect 26053 8375 26111 8381
rect 26326 8372 26332 8424
rect 26384 8372 26390 8424
rect 26421 8415 26479 8421
rect 26421 8381 26433 8415
rect 26467 8412 26479 8415
rect 26605 8415 26663 8421
rect 26605 8412 26617 8415
rect 26467 8384 26617 8412
rect 26467 8381 26479 8384
rect 26421 8375 26479 8381
rect 26605 8381 26617 8384
rect 26651 8381 26663 8415
rect 26605 8375 26663 8381
rect 24636 8316 25820 8344
rect 24636 8304 24642 8316
rect 21232 8248 22968 8276
rect 21232 8236 21238 8248
rect 23014 8236 23020 8288
rect 23072 8236 23078 8288
rect 24118 8236 24124 8288
rect 24176 8276 24182 8288
rect 24765 8279 24823 8285
rect 24765 8276 24777 8279
rect 24176 8248 24777 8276
rect 24176 8236 24182 8248
rect 24765 8245 24777 8248
rect 24811 8245 24823 8279
rect 24765 8239 24823 8245
rect 25038 8236 25044 8288
rect 25096 8236 25102 8288
rect 25590 8236 25596 8288
rect 25648 8236 25654 8288
rect 25869 8279 25927 8285
rect 25869 8245 25881 8279
rect 25915 8276 25927 8279
rect 26145 8279 26203 8285
rect 26145 8276 26157 8279
rect 25915 8248 26157 8276
rect 25915 8245 25927 8248
rect 25869 8239 25927 8245
rect 26145 8245 26157 8248
rect 26191 8245 26203 8279
rect 26145 8239 26203 8245
rect 552 8186 31531 8208
rect 552 8134 8102 8186
rect 8154 8134 8166 8186
rect 8218 8134 8230 8186
rect 8282 8134 8294 8186
rect 8346 8134 8358 8186
rect 8410 8134 15807 8186
rect 15859 8134 15871 8186
rect 15923 8134 15935 8186
rect 15987 8134 15999 8186
rect 16051 8134 16063 8186
rect 16115 8134 23512 8186
rect 23564 8134 23576 8186
rect 23628 8134 23640 8186
rect 23692 8134 23704 8186
rect 23756 8134 23768 8186
rect 23820 8134 31217 8186
rect 31269 8134 31281 8186
rect 31333 8134 31345 8186
rect 31397 8134 31409 8186
rect 31461 8134 31473 8186
rect 31525 8134 31531 8186
rect 552 8112 31531 8134
rect 7650 8032 7656 8084
rect 7708 8032 7714 8084
rect 7742 8032 7748 8084
rect 7800 8032 7806 8084
rect 8478 8032 8484 8084
rect 8536 8072 8542 8084
rect 8536 8044 8616 8072
rect 8536 8032 8542 8044
rect 7193 7939 7251 7945
rect 7193 7905 7205 7939
rect 7239 7936 7251 7939
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 7239 7908 7389 7936
rect 7239 7905 7251 7908
rect 7193 7899 7251 7905
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7936 7527 7939
rect 7668 7936 7696 8032
rect 7760 7945 7788 8032
rect 7515 7908 7696 7936
rect 7515 7905 7527 7908
rect 7469 7899 7527 7905
rect 7668 7800 7696 7908
rect 7745 7939 7803 7945
rect 7745 7905 7757 7939
rect 7791 7905 7803 7939
rect 7745 7899 7803 7905
rect 8018 7896 8024 7948
rect 8076 7896 8082 7948
rect 8294 7896 8300 7948
rect 8352 7896 8358 7948
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 8478 7936 8484 7948
rect 8435 7908 8484 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 8588 7936 8616 8044
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8812 8044 9045 8072
rect 8812 8032 8818 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 9582 8032 9588 8084
rect 9640 8032 9646 8084
rect 9674 8032 9680 8084
rect 9732 8032 9738 8084
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10413 8075 10471 8081
rect 10413 8072 10425 8075
rect 9916 8044 10425 8072
rect 9916 8032 9922 8044
rect 10413 8041 10425 8044
rect 10459 8041 10471 8075
rect 10413 8035 10471 8041
rect 10594 8032 10600 8084
rect 10652 8032 10658 8084
rect 10686 8032 10692 8084
rect 10744 8032 10750 8084
rect 17586 8072 17592 8084
rect 12728 8044 17592 8072
rect 8772 7976 9260 8004
rect 8665 7939 8723 7945
rect 8665 7936 8677 7939
rect 8588 7908 8677 7936
rect 8665 7905 8677 7908
rect 8711 7905 8723 7939
rect 8665 7899 8723 7905
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8570 7868 8576 7880
rect 7975 7840 8576 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 8772 7877 8800 7976
rect 8941 7939 8999 7945
rect 8941 7905 8953 7939
rect 8987 7936 8999 7939
rect 8987 7908 9076 7936
rect 8987 7905 8999 7908
rect 8941 7899 8999 7905
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 7668 7772 7788 7800
rect 7101 7735 7159 7741
rect 7101 7701 7113 7735
rect 7147 7732 7159 7735
rect 7190 7732 7196 7744
rect 7147 7704 7196 7732
rect 7147 7701 7159 7704
rect 7101 7695 7159 7701
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 7650 7692 7656 7744
rect 7708 7692 7714 7744
rect 7760 7732 7788 7772
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 8481 7803 8539 7809
rect 8168 7772 8432 7800
rect 8168 7760 8174 7772
rect 8205 7735 8263 7741
rect 8205 7732 8217 7735
rect 7760 7704 8217 7732
rect 8205 7701 8217 7704
rect 8251 7701 8263 7735
rect 8404 7732 8432 7772
rect 8481 7769 8493 7803
rect 8527 7800 8539 7803
rect 8846 7800 8852 7812
rect 8527 7772 8852 7800
rect 8527 7769 8539 7772
rect 8481 7763 8539 7769
rect 8846 7760 8852 7772
rect 8904 7760 8910 7812
rect 9048 7732 9076 7908
rect 9232 7868 9260 7976
rect 9401 7939 9459 7945
rect 9401 7905 9413 7939
rect 9447 7936 9459 7939
rect 9600 7936 9628 8032
rect 9692 8004 9720 8032
rect 9692 7976 9996 8004
rect 9968 7945 9996 7976
rect 9447 7908 9628 7936
rect 9677 7939 9735 7945
rect 9447 7905 9459 7908
rect 9401 7899 9459 7905
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 9953 7939 10011 7945
rect 9723 7908 9757 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 9953 7905 9965 7939
rect 9999 7905 10011 7939
rect 9953 7899 10011 7905
rect 9692 7868 9720 7899
rect 10226 7896 10232 7948
rect 10284 7896 10290 7948
rect 10318 7896 10324 7948
rect 10376 7896 10382 7948
rect 10612 7945 10640 8032
rect 10704 8004 10732 8032
rect 10965 8007 11023 8013
rect 10965 8004 10977 8007
rect 10704 7976 10977 8004
rect 10965 7973 10977 7976
rect 11011 8004 11023 8007
rect 11514 8004 11520 8016
rect 11011 7976 11520 8004
rect 11011 7973 11023 7976
rect 10965 7967 11023 7973
rect 11514 7964 11520 7976
rect 11572 7964 11578 8016
rect 12728 8013 12756 8044
rect 17586 8032 17592 8044
rect 17644 8072 17650 8084
rect 20901 8075 20959 8081
rect 17644 8044 20208 8072
rect 17644 8032 17650 8044
rect 12713 8007 12771 8013
rect 12713 7973 12725 8007
rect 12759 7973 12771 8007
rect 12713 7967 12771 7973
rect 12894 7964 12900 8016
rect 12952 8004 12958 8016
rect 13510 8007 13568 8013
rect 13510 8004 13522 8007
rect 12952 7976 13522 8004
rect 12952 7964 12958 7976
rect 13510 7973 13522 7976
rect 13556 7973 13568 8007
rect 13510 7967 13568 7973
rect 13722 7964 13728 8016
rect 13780 8004 13786 8016
rect 13780 7976 14964 8004
rect 13780 7964 13786 7976
rect 10597 7939 10655 7945
rect 10597 7905 10609 7939
rect 10643 7905 10655 7939
rect 10597 7899 10655 7905
rect 10778 7896 10784 7948
rect 10836 7896 10842 7948
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7905 13047 7939
rect 12989 7899 13047 7905
rect 10042 7868 10048 7880
rect 9232 7840 10048 7868
rect 10042 7828 10048 7840
rect 10100 7868 10106 7880
rect 10796 7868 10824 7896
rect 10100 7840 10824 7868
rect 10100 7828 10106 7840
rect 9490 7760 9496 7812
rect 9548 7800 9554 7812
rect 10137 7803 10195 7809
rect 10137 7800 10149 7803
rect 9548 7772 10149 7800
rect 9548 7760 9554 7772
rect 10137 7769 10149 7772
rect 10183 7769 10195 7803
rect 10137 7763 10195 7769
rect 11146 7760 11152 7812
rect 11204 7800 11210 7812
rect 11698 7800 11704 7812
rect 11204 7772 11704 7800
rect 11204 7760 11210 7772
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 8404 7704 9076 7732
rect 8205 7695 8263 7701
rect 9122 7692 9128 7744
rect 9180 7732 9186 7744
rect 9309 7735 9367 7741
rect 9309 7732 9321 7735
rect 9180 7704 9321 7732
rect 9180 7692 9186 7704
rect 9309 7701 9321 7704
rect 9355 7701 9367 7735
rect 9309 7695 9367 7701
rect 9582 7692 9588 7744
rect 9640 7692 9646 7744
rect 9858 7692 9864 7744
rect 9916 7692 9922 7744
rect 10689 7735 10747 7741
rect 10689 7701 10701 7735
rect 10735 7732 10747 7735
rect 12618 7732 12624 7744
rect 10735 7704 12624 7732
rect 10735 7701 10747 7704
rect 10689 7695 10747 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 13004 7732 13032 7899
rect 13262 7896 13268 7948
rect 13320 7896 13326 7948
rect 14826 7936 14832 7948
rect 13372 7908 14832 7936
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7868 13139 7871
rect 13372 7868 13400 7908
rect 14826 7896 14832 7908
rect 14884 7896 14890 7948
rect 14936 7945 14964 7976
rect 15286 7964 15292 8016
rect 15344 7964 15350 8016
rect 18325 8007 18383 8013
rect 18325 8004 18337 8007
rect 15672 7976 15884 8004
rect 15672 7945 15700 7976
rect 14921 7939 14979 7945
rect 14921 7905 14933 7939
rect 14967 7905 14979 7939
rect 14921 7899 14979 7905
rect 15389 7937 15447 7943
rect 15389 7903 15401 7937
rect 15435 7934 15447 7937
rect 15565 7939 15623 7945
rect 15565 7936 15577 7939
rect 15488 7934 15577 7936
rect 15435 7908 15577 7934
rect 15435 7906 15516 7908
rect 15435 7903 15447 7906
rect 13127 7840 13400 7868
rect 14936 7868 14964 7899
rect 15389 7897 15447 7903
rect 15565 7905 15577 7908
rect 15611 7905 15623 7939
rect 15565 7899 15623 7905
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 15749 7939 15807 7945
rect 15749 7905 15761 7939
rect 15795 7905 15807 7939
rect 15749 7899 15807 7905
rect 15672 7868 15700 7899
rect 14936 7840 15700 7868
rect 13127 7837 13139 7840
rect 13081 7831 13139 7837
rect 15580 7812 15608 7840
rect 15562 7760 15568 7812
rect 15620 7760 15626 7812
rect 13170 7732 13176 7744
rect 13004 7704 13176 7732
rect 13170 7692 13176 7704
rect 13228 7732 13234 7744
rect 14274 7732 14280 7744
rect 13228 7704 14280 7732
rect 13228 7692 13234 7704
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 14366 7692 14372 7744
rect 14424 7732 14430 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 14424 7704 14657 7732
rect 14424 7692 14430 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 14645 7695 14703 7701
rect 15013 7735 15071 7741
rect 15013 7701 15025 7735
rect 15059 7732 15071 7735
rect 15764 7732 15792 7899
rect 15856 7868 15884 7976
rect 16224 7976 18337 8004
rect 16224 7948 16252 7976
rect 18325 7973 18337 7976
rect 18371 8004 18383 8007
rect 18782 8004 18788 8016
rect 18371 7976 18788 8004
rect 18371 7973 18383 7976
rect 18325 7967 18383 7973
rect 18782 7964 18788 7976
rect 18840 7964 18846 8016
rect 19334 7964 19340 8016
rect 19392 8004 19398 8016
rect 20073 8007 20131 8013
rect 20073 8004 20085 8007
rect 19392 7976 20085 8004
rect 19392 7964 19398 7976
rect 20073 7973 20085 7976
rect 20119 7973 20131 8007
rect 20180 8004 20208 8044
rect 20901 8041 20913 8075
rect 20947 8072 20959 8075
rect 23014 8072 23020 8084
rect 20947 8044 23020 8072
rect 20947 8041 20959 8044
rect 20901 8035 20959 8041
rect 23014 8032 23020 8044
rect 23072 8032 23078 8084
rect 25590 8072 25596 8084
rect 23216 8044 25596 8072
rect 21269 8007 21327 8013
rect 21269 8004 21281 8007
rect 20180 7976 21281 8004
rect 20073 7967 20131 7973
rect 21269 7973 21281 7976
rect 21315 7973 21327 8007
rect 21269 7967 21327 7973
rect 21450 7964 21456 8016
rect 21508 8004 21514 8016
rect 21910 8004 21916 8016
rect 21508 7976 21916 8004
rect 21508 7964 21514 7976
rect 21910 7964 21916 7976
rect 21968 8004 21974 8016
rect 22833 8007 22891 8013
rect 22833 8004 22845 8007
rect 21968 7976 22845 8004
rect 21968 7964 21974 7976
rect 22833 7973 22845 7976
rect 22879 7973 22891 8007
rect 22833 7967 22891 7973
rect 16206 7896 16212 7948
rect 16264 7896 16270 7948
rect 16485 7939 16543 7945
rect 16485 7905 16497 7939
rect 16531 7905 16543 7939
rect 16485 7899 16543 7905
rect 16761 7939 16819 7945
rect 16761 7905 16773 7939
rect 16807 7936 16819 7939
rect 16850 7936 16856 7948
rect 16807 7908 16856 7936
rect 16807 7905 16819 7908
rect 16761 7899 16819 7905
rect 16500 7868 16528 7899
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 17028 7939 17086 7945
rect 17028 7905 17040 7939
rect 17074 7936 17086 7939
rect 18506 7936 18512 7948
rect 17074 7908 18512 7936
rect 17074 7905 17086 7908
rect 17028 7899 17086 7905
rect 18506 7896 18512 7908
rect 18564 7896 18570 7948
rect 20165 7939 20223 7945
rect 20165 7936 20177 7939
rect 19076 7908 20177 7936
rect 15856 7840 16528 7868
rect 19076 7812 19104 7908
rect 20165 7905 20177 7908
rect 20211 7905 20223 7939
rect 20165 7899 20223 7905
rect 20441 7939 20499 7945
rect 20441 7905 20453 7939
rect 20487 7905 20499 7939
rect 20441 7899 20499 7905
rect 20993 7939 21051 7945
rect 20993 7905 21005 7939
rect 21039 7936 21051 7939
rect 21726 7936 21732 7948
rect 21039 7908 21732 7936
rect 21039 7905 21051 7908
rect 20993 7899 21051 7905
rect 20254 7828 20260 7880
rect 20312 7868 20318 7880
rect 20456 7868 20484 7899
rect 21726 7896 21732 7908
rect 21784 7896 21790 7948
rect 22848 7936 22876 7967
rect 22922 7936 22928 7948
rect 22848 7908 22928 7936
rect 22922 7896 22928 7908
rect 22980 7936 22986 7948
rect 23098 7939 23156 7945
rect 23098 7936 23110 7939
rect 22980 7908 23110 7936
rect 22980 7896 22986 7908
rect 23098 7905 23110 7908
rect 23144 7905 23156 7939
rect 23098 7899 23156 7905
rect 20312 7840 20484 7868
rect 20312 7828 20318 7840
rect 22094 7828 22100 7880
rect 22152 7868 22158 7880
rect 23216 7868 23244 8044
rect 25590 8032 25596 8044
rect 25648 8032 25654 8084
rect 23376 8007 23434 8013
rect 23376 7973 23388 8007
rect 23422 8004 23434 8007
rect 25498 8004 25504 8016
rect 23422 7976 25504 8004
rect 23422 7973 23434 7976
rect 23376 7967 23434 7973
rect 25498 7964 25504 7976
rect 25556 7964 25562 8016
rect 25700 7976 26096 8004
rect 24673 7939 24731 7945
rect 24673 7905 24685 7939
rect 24719 7905 24731 7939
rect 24673 7899 24731 7905
rect 24949 7939 25007 7945
rect 24949 7905 24961 7939
rect 24995 7936 25007 7939
rect 25130 7936 25136 7948
rect 24995 7908 25136 7936
rect 24995 7905 25007 7908
rect 24949 7899 25007 7905
rect 22152 7840 23244 7868
rect 22152 7828 22158 7840
rect 19058 7800 19064 7812
rect 16500 7772 16804 7800
rect 16500 7744 16528 7772
rect 15059 7704 15792 7732
rect 15059 7701 15071 7704
rect 15013 7695 15071 7701
rect 15838 7692 15844 7744
rect 15896 7692 15902 7744
rect 16298 7692 16304 7744
rect 16356 7692 16362 7744
rect 16482 7692 16488 7744
rect 16540 7692 16546 7744
rect 16577 7735 16635 7741
rect 16577 7701 16589 7735
rect 16623 7732 16635 7735
rect 16666 7732 16672 7744
rect 16623 7704 16672 7732
rect 16623 7701 16635 7704
rect 16577 7695 16635 7701
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 16776 7732 16804 7772
rect 17972 7772 19064 7800
rect 17972 7744 18000 7772
rect 19058 7760 19064 7772
rect 19116 7760 19122 7812
rect 19518 7760 19524 7812
rect 19576 7800 19582 7812
rect 20533 7803 20591 7809
rect 20533 7800 20545 7803
rect 19576 7772 20545 7800
rect 19576 7760 19582 7772
rect 20533 7769 20545 7772
rect 20579 7769 20591 7803
rect 24688 7800 24716 7899
rect 25130 7896 25136 7908
rect 25188 7896 25194 7948
rect 25222 7896 25228 7948
rect 25280 7896 25286 7948
rect 25406 7896 25412 7948
rect 25464 7936 25470 7948
rect 25700 7945 25728 7976
rect 26068 7945 26096 7976
rect 25685 7939 25743 7945
rect 25685 7936 25697 7939
rect 25464 7908 25697 7936
rect 25464 7896 25470 7908
rect 25685 7905 25697 7908
rect 25731 7905 25743 7939
rect 26053 7939 26111 7945
rect 25685 7899 25743 7905
rect 25777 7929 25835 7935
rect 25777 7895 25789 7929
rect 25823 7895 25835 7929
rect 26053 7905 26065 7939
rect 26099 7905 26111 7939
rect 26053 7899 26111 7905
rect 25777 7889 25835 7895
rect 24762 7828 24768 7880
rect 24820 7828 24826 7880
rect 25317 7871 25375 7877
rect 25317 7837 25329 7871
rect 25363 7868 25375 7871
rect 25590 7868 25596 7880
rect 25363 7840 25596 7868
rect 25363 7837 25375 7840
rect 25317 7831 25375 7837
rect 25590 7828 25596 7840
rect 25648 7828 25654 7880
rect 25498 7800 25504 7812
rect 20533 7763 20591 7769
rect 24044 7772 24716 7800
rect 24780 7772 25504 7800
rect 17954 7732 17960 7744
rect 16776 7704 17960 7732
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18138 7692 18144 7744
rect 18196 7692 18202 7744
rect 19978 7692 19984 7744
rect 20036 7732 20042 7744
rect 20257 7735 20315 7741
rect 20257 7732 20269 7735
rect 20036 7704 20269 7732
rect 20036 7692 20042 7704
rect 20257 7701 20269 7704
rect 20303 7701 20315 7735
rect 20257 7695 20315 7701
rect 21726 7692 21732 7744
rect 21784 7732 21790 7744
rect 24044 7732 24072 7772
rect 21784 7704 24072 7732
rect 24489 7735 24547 7741
rect 21784 7692 21790 7704
rect 24489 7701 24501 7735
rect 24535 7732 24547 7735
rect 24780 7732 24808 7772
rect 25498 7760 25504 7772
rect 25556 7760 25562 7812
rect 25792 7744 25820 7889
rect 24535 7704 24808 7732
rect 24535 7701 24547 7704
rect 24489 7695 24547 7701
rect 24854 7692 24860 7744
rect 24912 7732 24918 7744
rect 25041 7735 25099 7741
rect 25041 7732 25053 7735
rect 24912 7704 25053 7732
rect 24912 7692 24918 7704
rect 25041 7701 25053 7704
rect 25087 7701 25099 7735
rect 25041 7695 25099 7701
rect 25593 7735 25651 7741
rect 25593 7701 25605 7735
rect 25639 7732 25651 7735
rect 25682 7732 25688 7744
rect 25639 7704 25688 7732
rect 25639 7701 25651 7704
rect 25593 7695 25651 7701
rect 25682 7692 25688 7704
rect 25740 7692 25746 7744
rect 25774 7692 25780 7744
rect 25832 7692 25838 7744
rect 25866 7692 25872 7744
rect 25924 7692 25930 7744
rect 26142 7692 26148 7744
rect 26200 7692 26206 7744
rect 552 7642 31372 7664
rect 552 7590 4250 7642
rect 4302 7590 4314 7642
rect 4366 7590 4378 7642
rect 4430 7590 4442 7642
rect 4494 7590 4506 7642
rect 4558 7590 11955 7642
rect 12007 7590 12019 7642
rect 12071 7590 12083 7642
rect 12135 7590 12147 7642
rect 12199 7590 12211 7642
rect 12263 7590 19660 7642
rect 19712 7590 19724 7642
rect 19776 7590 19788 7642
rect 19840 7590 19852 7642
rect 19904 7590 19916 7642
rect 19968 7590 27365 7642
rect 27417 7590 27429 7642
rect 27481 7590 27493 7642
rect 27545 7590 27557 7642
rect 27609 7590 27621 7642
rect 27673 7590 31372 7642
rect 552 7568 31372 7590
rect 7006 7488 7012 7540
rect 7064 7488 7070 7540
rect 7558 7528 7564 7540
rect 7208 7500 7564 7528
rect 6227 7463 6285 7469
rect 6227 7429 6239 7463
rect 6273 7460 6285 7463
rect 7208 7460 7236 7500
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 7834 7488 7840 7540
rect 7892 7528 7898 7540
rect 8110 7528 8116 7540
rect 7892 7500 8116 7528
rect 7892 7488 7898 7500
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 8352 7500 8861 7528
rect 8352 7488 8358 7500
rect 8849 7497 8861 7500
rect 8895 7497 8907 7531
rect 8849 7491 8907 7497
rect 9125 7531 9183 7537
rect 9125 7497 9137 7531
rect 9171 7528 9183 7531
rect 9582 7528 9588 7540
rect 9171 7500 9588 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 10689 7531 10747 7537
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 11330 7528 11336 7540
rect 10735 7500 11336 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 14369 7531 14427 7537
rect 12268 7500 14320 7528
rect 6273 7432 7236 7460
rect 7285 7463 7343 7469
rect 6273 7429 6285 7432
rect 6227 7423 6285 7429
rect 7285 7429 7297 7463
rect 7331 7460 7343 7463
rect 9214 7460 9220 7472
rect 7331 7432 9220 7460
rect 7331 7429 7343 7432
rect 7285 7423 7343 7429
rect 9214 7420 9220 7432
rect 9272 7420 9278 7472
rect 12268 7460 12296 7500
rect 9416 7432 10088 7460
rect 8754 7392 8760 7404
rect 8036 7364 8760 7392
rect 6156 7327 6214 7333
rect 6156 7293 6168 7327
rect 6202 7324 6214 7327
rect 6411 7327 6469 7333
rect 6411 7324 6423 7327
rect 6202 7296 6423 7324
rect 6202 7293 6214 7296
rect 6156 7287 6214 7293
rect 6411 7293 6423 7296
rect 6457 7293 6469 7327
rect 6411 7287 6469 7293
rect 6514 7327 6572 7333
rect 6514 7293 6526 7327
rect 6560 7324 6572 7327
rect 6708 7327 6766 7333
rect 6560 7293 6592 7324
rect 6514 7287 6592 7293
rect 6708 7293 6720 7327
rect 6754 7324 6766 7327
rect 7006 7324 7012 7336
rect 6754 7296 7012 7324
rect 6754 7293 6766 7296
rect 6708 7287 6766 7293
rect 6564 7256 6592 7287
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7098 7284 7104 7336
rect 7156 7284 7162 7336
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 7282 7324 7288 7336
rect 7239 7296 7288 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 7650 7333 7656 7336
rect 7645 7324 7656 7333
rect 7611 7296 7656 7324
rect 7645 7287 7656 7296
rect 7650 7284 7656 7287
rect 7708 7284 7714 7336
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7324 7987 7327
rect 8036 7324 8064 7364
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 9122 7392 9128 7404
rect 9048 7364 9128 7392
rect 7975 7296 8064 7324
rect 7975 7293 7987 7296
rect 7929 7287 7987 7293
rect 6564 7228 7144 7256
rect 7116 7200 7144 7228
rect 6779 7191 6837 7197
rect 6779 7157 6791 7191
rect 6825 7188 6837 7191
rect 6914 7188 6920 7200
rect 6825 7160 6920 7188
rect 6825 7157 6837 7160
rect 6779 7151 6837 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7098 7148 7104 7200
rect 7156 7148 7162 7200
rect 7561 7191 7619 7197
rect 7561 7157 7573 7191
rect 7607 7188 7619 7191
rect 7650 7188 7656 7200
rect 7607 7160 7656 7188
rect 7607 7157 7619 7160
rect 7561 7151 7619 7157
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 7760 7188 7788 7287
rect 8110 7284 8116 7336
rect 8168 7324 8174 7336
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 8168 7296 8217 7324
rect 8168 7284 8174 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 7837 7259 7895 7265
rect 7837 7225 7849 7259
rect 7883 7256 7895 7259
rect 8478 7256 8484 7268
rect 7883 7228 8484 7256
rect 7883 7225 7895 7228
rect 7837 7219 7895 7225
rect 8478 7216 8484 7228
rect 8536 7216 8542 7268
rect 8680 7256 8708 7287
rect 8938 7284 8944 7336
rect 8996 7284 9002 7336
rect 9048 7333 9076 7364
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 9416 7392 9444 7432
rect 9324 7364 9444 7392
rect 9324 7336 9352 7364
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 9858 7392 9864 7404
rect 9640 7364 9864 7392
rect 9640 7352 9646 7364
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 10060 7401 10088 7432
rect 10336 7432 12296 7460
rect 14292 7460 14320 7500
rect 14369 7497 14381 7531
rect 14415 7528 14427 7531
rect 15286 7528 15292 7540
rect 14415 7500 15292 7528
rect 14415 7497 14427 7500
rect 14369 7491 14427 7497
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15473 7531 15531 7537
rect 15473 7497 15485 7531
rect 15519 7497 15531 7531
rect 15473 7491 15531 7497
rect 15749 7531 15807 7537
rect 15749 7497 15761 7531
rect 15795 7528 15807 7531
rect 15838 7528 15844 7540
rect 15795 7500 15844 7528
rect 15795 7497 15807 7500
rect 15749 7491 15807 7497
rect 14458 7460 14464 7472
rect 14292 7432 14464 7460
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 9033 7327 9091 7333
rect 9033 7293 9045 7327
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 9214 7284 9220 7336
rect 9272 7284 9278 7336
rect 9306 7284 9312 7336
rect 9364 7284 9370 7336
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7324 9459 7327
rect 9490 7324 9496 7336
rect 9447 7296 9496 7324
rect 9447 7293 9459 7296
rect 9401 7287 9459 7293
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 9766 7284 9772 7336
rect 9824 7284 9830 7336
rect 10134 7284 10140 7336
rect 10192 7324 10198 7336
rect 10336 7333 10364 7432
rect 14458 7420 14464 7432
rect 14516 7420 14522 7472
rect 15488 7460 15516 7491
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 16850 7488 16856 7540
rect 16908 7528 16914 7540
rect 17770 7528 17776 7540
rect 16908 7500 17776 7528
rect 16908 7488 16914 7500
rect 16482 7460 16488 7472
rect 15120 7432 15516 7460
rect 16132 7432 16488 7460
rect 11238 7392 11244 7404
rect 10888 7364 11244 7392
rect 10888 7333 10916 7364
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 11698 7392 11704 7404
rect 11348 7364 11704 7392
rect 11348 7333 11376 7364
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 10321 7327 10379 7333
rect 10321 7324 10333 7327
rect 10192 7296 10333 7324
rect 10192 7284 10198 7296
rect 10321 7293 10333 7296
rect 10367 7293 10379 7327
rect 10321 7287 10379 7293
rect 10597 7327 10655 7333
rect 10597 7293 10609 7327
rect 10643 7293 10655 7327
rect 10597 7287 10655 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7293 10931 7327
rect 10873 7287 10931 7293
rect 11057 7327 11115 7333
rect 11057 7293 11069 7327
rect 11103 7293 11115 7327
rect 11057 7287 11115 7293
rect 11333 7327 11391 7333
rect 11333 7293 11345 7327
rect 11379 7293 11391 7327
rect 11333 7287 11391 7293
rect 11609 7327 11667 7333
rect 11609 7293 11621 7327
rect 11655 7324 11667 7327
rect 12526 7324 12532 7336
rect 11655 7296 12532 7324
rect 11655 7293 11667 7296
rect 11609 7287 11667 7293
rect 9858 7256 9864 7268
rect 8680 7228 9864 7256
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 10410 7216 10416 7268
rect 10468 7256 10474 7268
rect 10612 7256 10640 7287
rect 11072 7256 11100 7287
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 12618 7284 12624 7336
rect 12676 7324 12682 7336
rect 12906 7327 12964 7333
rect 12906 7324 12918 7327
rect 12676 7296 12918 7324
rect 12676 7284 12682 7296
rect 12906 7293 12918 7296
rect 12952 7293 12964 7327
rect 12906 7287 12964 7293
rect 13173 7327 13231 7333
rect 13173 7293 13185 7327
rect 13219 7324 13231 7327
rect 13262 7324 13268 7336
rect 13219 7296 13268 7324
rect 13219 7293 13231 7296
rect 13173 7287 13231 7293
rect 13262 7284 13268 7296
rect 13320 7324 13326 7336
rect 13630 7324 13636 7336
rect 13320 7296 13636 7324
rect 13320 7284 13326 7296
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 13722 7284 13728 7336
rect 13780 7284 13786 7336
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 13964 7296 14013 7324
rect 13964 7284 13970 7296
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 14274 7284 14280 7336
rect 14332 7284 14338 7336
rect 14550 7284 14556 7336
rect 14608 7284 14614 7336
rect 14737 7327 14795 7333
rect 14737 7293 14749 7327
rect 14783 7293 14795 7327
rect 14737 7287 14795 7293
rect 15013 7327 15071 7333
rect 15013 7293 15025 7327
rect 15059 7324 15071 7327
rect 15120 7324 15148 7432
rect 15059 7296 15148 7324
rect 15289 7327 15347 7333
rect 15059 7293 15071 7296
rect 15013 7287 15071 7293
rect 15289 7293 15301 7327
rect 15335 7324 15347 7327
rect 15335 7296 15516 7324
rect 15335 7293 15347 7296
rect 15289 7287 15347 7293
rect 12710 7256 12716 7268
rect 10468 7228 10916 7256
rect 11072 7228 12716 7256
rect 10468 7216 10474 7228
rect 10888 7200 10916 7228
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 13817 7259 13875 7265
rect 13817 7225 13829 7259
rect 13863 7256 13875 7259
rect 14642 7256 14648 7268
rect 13863 7228 14648 7256
rect 13863 7225 13875 7228
rect 13817 7219 13875 7225
rect 14642 7216 14648 7228
rect 14700 7216 14706 7268
rect 14752 7256 14780 7287
rect 15378 7256 15384 7268
rect 14752 7228 15384 7256
rect 15378 7216 15384 7228
rect 15436 7216 15442 7268
rect 8113 7191 8171 7197
rect 8113 7188 8125 7191
rect 7760 7160 8125 7188
rect 8113 7157 8125 7160
rect 8159 7157 8171 7191
rect 8113 7151 8171 7157
rect 8573 7191 8631 7197
rect 8573 7157 8585 7191
rect 8619 7188 8631 7191
rect 9214 7188 9220 7200
rect 8619 7160 9220 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 9677 7191 9735 7197
rect 9677 7157 9689 7191
rect 9723 7188 9735 7191
rect 10502 7188 10508 7200
rect 9723 7160 10508 7188
rect 9723 7157 9735 7160
rect 9677 7151 9735 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10870 7148 10876 7200
rect 10928 7148 10934 7200
rect 11054 7148 11060 7200
rect 11112 7148 11118 7200
rect 11241 7191 11299 7197
rect 11241 7157 11253 7191
rect 11287 7188 11299 7191
rect 11330 7188 11336 7200
rect 11287 7160 11336 7188
rect 11287 7157 11299 7160
rect 11241 7151 11299 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11514 7148 11520 7200
rect 11572 7148 11578 7200
rect 11790 7148 11796 7200
rect 11848 7148 11854 7200
rect 14090 7148 14096 7200
rect 14148 7148 14154 7200
rect 14737 7191 14795 7197
rect 14737 7157 14749 7191
rect 14783 7188 14795 7191
rect 14826 7188 14832 7200
rect 14783 7160 14832 7188
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 14826 7148 14832 7160
rect 14884 7148 14890 7200
rect 14918 7148 14924 7200
rect 14976 7148 14982 7200
rect 15194 7148 15200 7200
rect 15252 7148 15258 7200
rect 15488 7188 15516 7296
rect 15562 7284 15568 7336
rect 15620 7284 15626 7336
rect 16132 7333 16160 7432
rect 16482 7420 16488 7432
rect 16540 7460 16546 7472
rect 16540 7432 16988 7460
rect 16540 7420 16546 7432
rect 16298 7392 16304 7404
rect 16224 7364 16304 7392
rect 16224 7333 16252 7364
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 16577 7395 16635 7401
rect 16577 7392 16589 7395
rect 16408 7364 16589 7392
rect 16408 7333 16436 7364
rect 16577 7361 16589 7364
rect 16623 7361 16635 7395
rect 16577 7355 16635 7361
rect 16758 7352 16764 7404
rect 16816 7392 16822 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16816 7364 16865 7392
rect 16816 7352 16822 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 16666 7333 16672 7336
rect 15841 7327 15899 7333
rect 15841 7293 15853 7327
rect 15887 7324 15899 7327
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 15887 7296 16037 7324
rect 15887 7293 15899 7296
rect 15841 7287 15899 7293
rect 16025 7293 16037 7296
rect 16071 7293 16083 7327
rect 16025 7287 16083 7293
rect 16117 7327 16175 7333
rect 16117 7293 16129 7327
rect 16163 7293 16175 7327
rect 16117 7287 16175 7293
rect 16209 7327 16267 7333
rect 16209 7293 16221 7327
rect 16255 7293 16267 7327
rect 16209 7287 16267 7293
rect 16393 7327 16451 7333
rect 16393 7293 16405 7327
rect 16439 7293 16451 7327
rect 16393 7287 16451 7293
rect 16661 7287 16672 7333
rect 16724 7324 16730 7336
rect 16960 7333 16988 7432
rect 17052 7401 17080 7500
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 18782 7488 18788 7540
rect 18840 7528 18846 7540
rect 18840 7500 24164 7528
rect 18840 7488 18846 7500
rect 18598 7420 18604 7472
rect 18656 7460 18662 7472
rect 19337 7463 19395 7469
rect 19337 7460 19349 7463
rect 18656 7432 19349 7460
rect 18656 7420 18662 7432
rect 19337 7429 19349 7432
rect 19383 7429 19395 7463
rect 19337 7423 19395 7429
rect 19426 7420 19432 7472
rect 19484 7420 19490 7472
rect 19794 7420 19800 7472
rect 19852 7460 19858 7472
rect 19852 7432 20024 7460
rect 19852 7420 19858 7432
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7392 18843 7395
rect 18831 7364 19288 7392
rect 18831 7361 18843 7364
rect 18785 7355 18843 7361
rect 16945 7327 17003 7333
rect 16724 7296 16761 7324
rect 15654 7216 15660 7268
rect 15712 7256 15718 7268
rect 16132 7256 16160 7287
rect 16666 7284 16672 7287
rect 16724 7284 16730 7296
rect 16945 7293 16957 7327
rect 16991 7293 17003 7327
rect 16945 7287 17003 7293
rect 17126 7284 17132 7336
rect 17184 7284 17190 7336
rect 18690 7284 18696 7336
rect 18748 7284 18754 7336
rect 18874 7284 18880 7336
rect 18932 7284 18938 7336
rect 19058 7284 19064 7336
rect 19116 7324 19122 7336
rect 19260 7333 19288 7364
rect 19153 7327 19211 7333
rect 19153 7324 19165 7327
rect 19116 7296 19165 7324
rect 19116 7284 19122 7296
rect 19153 7293 19165 7296
rect 19199 7293 19211 7327
rect 19153 7287 19211 7293
rect 19245 7327 19303 7333
rect 19245 7293 19257 7327
rect 19291 7293 19303 7327
rect 19444 7324 19472 7420
rect 19610 7352 19616 7404
rect 19668 7352 19674 7404
rect 19996 7392 20024 7432
rect 23382 7420 23388 7472
rect 23440 7460 23446 7472
rect 23569 7463 23627 7469
rect 23569 7460 23581 7463
rect 23440 7432 23581 7460
rect 23440 7420 23446 7432
rect 23569 7429 23581 7432
rect 23615 7429 23627 7463
rect 23750 7460 23756 7472
rect 23569 7423 23627 7429
rect 23676 7432 23756 7460
rect 19996 7364 21220 7392
rect 19996 7333 20024 7364
rect 19521 7327 19579 7333
rect 19521 7324 19533 7327
rect 19444 7296 19533 7324
rect 19245 7287 19303 7293
rect 19521 7293 19533 7296
rect 19567 7293 19579 7327
rect 19521 7287 19579 7293
rect 19981 7327 20039 7333
rect 19981 7293 19993 7327
rect 20027 7293 20039 7327
rect 19981 7287 20039 7293
rect 20162 7284 20168 7336
rect 20220 7324 20226 7336
rect 20257 7329 20315 7335
rect 20640 7333 20668 7364
rect 21192 7333 21220 7364
rect 21910 7352 21916 7404
rect 21968 7352 21974 7404
rect 23676 7392 23704 7432
rect 23750 7420 23756 7432
rect 23808 7420 23814 7472
rect 24136 7460 24164 7500
rect 24486 7488 24492 7540
rect 24544 7488 24550 7540
rect 24578 7488 24584 7540
rect 24636 7528 24642 7540
rect 24765 7531 24823 7537
rect 24765 7528 24777 7531
rect 24636 7500 24777 7528
rect 24636 7488 24642 7500
rect 24765 7497 24777 7500
rect 24811 7497 24823 7531
rect 24765 7491 24823 7497
rect 25590 7488 25596 7540
rect 25648 7488 25654 7540
rect 25774 7488 25780 7540
rect 25832 7488 25838 7540
rect 25041 7463 25099 7469
rect 24136 7432 24716 7460
rect 23934 7392 23940 7404
rect 23584 7364 23704 7392
rect 23768 7364 23940 7392
rect 20257 7324 20269 7329
rect 20220 7296 20269 7324
rect 20220 7284 20226 7296
rect 20257 7295 20269 7296
rect 20303 7295 20315 7329
rect 20257 7289 20315 7295
rect 20349 7327 20407 7333
rect 20349 7293 20361 7327
rect 20395 7293 20407 7327
rect 20349 7287 20407 7293
rect 20625 7327 20683 7333
rect 20625 7293 20637 7327
rect 20671 7293 20683 7327
rect 20625 7287 20683 7293
rect 20717 7327 20775 7333
rect 20717 7293 20729 7327
rect 20763 7324 20775 7327
rect 20901 7327 20959 7333
rect 20901 7324 20913 7327
rect 20763 7296 20913 7324
rect 20763 7293 20775 7296
rect 20717 7287 20775 7293
rect 20901 7293 20913 7296
rect 20947 7293 20959 7327
rect 20901 7287 20959 7293
rect 21177 7327 21235 7333
rect 21177 7293 21189 7327
rect 21223 7293 21235 7327
rect 21177 7287 21235 7293
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 21453 7327 21511 7333
rect 21453 7324 21465 7327
rect 21315 7296 21465 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 21453 7293 21465 7296
rect 21499 7293 21511 7327
rect 21453 7287 21511 7293
rect 22180 7327 22238 7333
rect 22180 7293 22192 7327
rect 22226 7324 22238 7327
rect 23584 7324 23612 7364
rect 22226 7296 23612 7324
rect 23661 7327 23719 7333
rect 22226 7293 22238 7296
rect 22180 7287 22238 7293
rect 23661 7293 23673 7327
rect 23707 7324 23719 7327
rect 23768 7324 23796 7364
rect 23934 7352 23940 7364
rect 23992 7352 23998 7404
rect 23707 7296 23796 7324
rect 23845 7327 23903 7333
rect 23707 7293 23719 7296
rect 23661 7287 23719 7293
rect 23845 7293 23857 7327
rect 23891 7293 23903 7327
rect 23845 7287 23903 7293
rect 24029 7327 24087 7333
rect 24029 7293 24041 7327
rect 24075 7324 24087 7327
rect 24118 7324 24124 7336
rect 24075 7296 24124 7324
rect 24075 7293 24087 7296
rect 24029 7287 24087 7293
rect 15712 7228 16160 7256
rect 16301 7259 16359 7265
rect 15712 7216 15718 7228
rect 16301 7225 16313 7259
rect 16347 7256 16359 7259
rect 17144 7256 17172 7284
rect 16347 7228 17172 7256
rect 17304 7259 17362 7265
rect 16347 7225 16359 7228
rect 16301 7219 16359 7225
rect 17304 7225 17316 7259
rect 17350 7256 17362 7259
rect 18892 7256 18920 7284
rect 17350 7228 18920 7256
rect 17350 7225 17362 7228
rect 17304 7219 17362 7225
rect 18966 7216 18972 7268
rect 19024 7256 19030 7268
rect 20364 7256 20392 7287
rect 19024 7228 20392 7256
rect 19024 7216 19030 7228
rect 21358 7216 21364 7268
rect 21416 7256 21422 7268
rect 23860 7256 23888 7287
rect 24118 7284 24124 7296
rect 24176 7284 24182 7336
rect 24210 7284 24216 7336
rect 24268 7324 24274 7336
rect 24305 7327 24363 7333
rect 24305 7324 24317 7327
rect 24268 7296 24317 7324
rect 24268 7284 24274 7296
rect 24305 7293 24317 7296
rect 24351 7293 24363 7327
rect 24305 7287 24363 7293
rect 24486 7284 24492 7336
rect 24544 7324 24550 7336
rect 24688 7333 24716 7432
rect 25041 7429 25053 7463
rect 25087 7460 25099 7463
rect 25222 7460 25228 7472
rect 25087 7432 25228 7460
rect 25087 7429 25099 7432
rect 25041 7423 25099 7429
rect 25222 7420 25228 7432
rect 25280 7460 25286 7472
rect 25792 7460 25820 7488
rect 25280 7432 25820 7460
rect 25280 7420 25286 7432
rect 24581 7327 24639 7333
rect 24581 7324 24593 7327
rect 24544 7296 24593 7324
rect 24544 7284 24550 7296
rect 24581 7293 24593 7296
rect 24627 7293 24639 7327
rect 24581 7287 24639 7293
rect 24673 7327 24731 7333
rect 24673 7293 24685 7327
rect 24719 7293 24731 7327
rect 24673 7287 24731 7293
rect 24946 7284 24952 7336
rect 25004 7284 25010 7336
rect 25038 7284 25044 7336
rect 25096 7284 25102 7336
rect 25406 7324 25412 7336
rect 25240 7296 25412 7324
rect 21416 7228 23888 7256
rect 23937 7259 23995 7265
rect 21416 7216 21422 7228
rect 23937 7225 23949 7259
rect 23983 7256 23995 7259
rect 25056 7256 25084 7284
rect 23983 7228 25084 7256
rect 23983 7225 23995 7228
rect 23937 7219 23995 7225
rect 18322 7188 18328 7200
rect 15488 7160 18328 7188
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 18414 7148 18420 7200
rect 18472 7148 18478 7200
rect 18506 7148 18512 7200
rect 18564 7188 18570 7200
rect 19061 7191 19119 7197
rect 19061 7188 19073 7191
rect 18564 7160 19073 7188
rect 18564 7148 18570 7160
rect 19061 7157 19073 7160
rect 19107 7157 19119 7191
rect 19061 7151 19119 7157
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 19794 7188 19800 7200
rect 19208 7160 19800 7188
rect 19208 7148 19214 7160
rect 19794 7148 19800 7160
rect 19852 7148 19858 7200
rect 19886 7148 19892 7200
rect 19944 7148 19950 7200
rect 20162 7148 20168 7200
rect 20220 7148 20226 7200
rect 20346 7148 20352 7200
rect 20404 7188 20410 7200
rect 20441 7191 20499 7197
rect 20441 7188 20453 7191
rect 20404 7160 20453 7188
rect 20404 7148 20410 7160
rect 20441 7157 20453 7160
rect 20487 7157 20499 7191
rect 20441 7151 20499 7157
rect 20990 7148 20996 7200
rect 21048 7148 21054 7200
rect 21542 7148 21548 7200
rect 21600 7188 21606 7200
rect 23106 7188 23112 7200
rect 21600 7160 23112 7188
rect 21600 7148 21606 7160
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 23198 7148 23204 7200
rect 23256 7188 23262 7200
rect 23293 7191 23351 7197
rect 23293 7188 23305 7191
rect 23256 7160 23305 7188
rect 23256 7148 23262 7160
rect 23293 7157 23305 7160
rect 23339 7157 23351 7191
rect 23293 7151 23351 7157
rect 24118 7148 24124 7200
rect 24176 7188 24182 7200
rect 24213 7191 24271 7197
rect 24213 7188 24225 7191
rect 24176 7160 24225 7188
rect 24176 7148 24182 7160
rect 24213 7157 24225 7160
rect 24259 7157 24271 7191
rect 24213 7151 24271 7157
rect 25038 7148 25044 7200
rect 25096 7188 25102 7200
rect 25240 7188 25268 7296
rect 25406 7284 25412 7296
rect 25464 7284 25470 7336
rect 25498 7284 25504 7336
rect 25556 7284 25562 7336
rect 25096 7160 25268 7188
rect 25096 7148 25102 7160
rect 25314 7148 25320 7200
rect 25372 7148 25378 7200
rect 552 7098 31531 7120
rect 552 7046 8102 7098
rect 8154 7046 8166 7098
rect 8218 7046 8230 7098
rect 8282 7046 8294 7098
rect 8346 7046 8358 7098
rect 8410 7046 15807 7098
rect 15859 7046 15871 7098
rect 15923 7046 15935 7098
rect 15987 7046 15999 7098
rect 16051 7046 16063 7098
rect 16115 7046 23512 7098
rect 23564 7046 23576 7098
rect 23628 7046 23640 7098
rect 23692 7046 23704 7098
rect 23756 7046 23768 7098
rect 23820 7046 31217 7098
rect 31269 7046 31281 7098
rect 31333 7046 31345 7098
rect 31397 7046 31409 7098
rect 31461 7046 31473 7098
rect 31525 7046 31531 7098
rect 552 7024 31531 7046
rect 6914 6944 6920 6996
rect 6972 6944 6978 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7331 6987 7389 6993
rect 7331 6984 7343 6987
rect 7064 6956 7343 6984
rect 7064 6944 7070 6956
rect 7331 6953 7343 6956
rect 7377 6953 7389 6987
rect 7331 6947 7389 6953
rect 8018 6944 8024 6996
rect 8076 6984 8082 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 8076 6956 8217 6984
rect 8076 6944 8082 6956
rect 8205 6953 8217 6956
rect 8251 6953 8263 6987
rect 8205 6947 8263 6953
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 9217 6987 9275 6993
rect 9217 6984 9229 6987
rect 8536 6956 9229 6984
rect 8536 6944 8542 6956
rect 9217 6953 9229 6956
rect 9263 6953 9275 6987
rect 9217 6947 9275 6953
rect 9674 6944 9680 6996
rect 9732 6944 9738 6996
rect 9766 6944 9772 6996
rect 9824 6984 9830 6996
rect 10413 6987 10471 6993
rect 10413 6984 10425 6987
rect 9824 6956 10425 6984
rect 9824 6944 9830 6956
rect 10413 6953 10425 6956
rect 10459 6953 10471 6987
rect 10413 6947 10471 6953
rect 10502 6944 10508 6996
rect 10560 6944 10566 6996
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 12253 6987 12311 6993
rect 12253 6984 12265 6987
rect 11112 6956 12265 6984
rect 11112 6944 11118 6956
rect 12253 6953 12265 6956
rect 12299 6953 12311 6987
rect 12253 6947 12311 6953
rect 14550 6944 14556 6996
rect 14608 6944 14614 6996
rect 15378 6944 15384 6996
rect 15436 6984 15442 6996
rect 15841 6987 15899 6993
rect 15841 6984 15853 6987
rect 15436 6956 15853 6984
rect 15436 6944 15442 6956
rect 15841 6953 15853 6956
rect 15887 6953 15899 6987
rect 16577 6987 16635 6993
rect 16577 6984 16589 6987
rect 15841 6947 15899 6953
rect 15948 6956 16589 6984
rect 6546 6857 6552 6860
rect 6248 6851 6306 6857
rect 6248 6817 6260 6851
rect 6294 6848 6306 6851
rect 6524 6851 6552 6857
rect 6294 6820 6408 6848
rect 6294 6817 6306 6820
rect 6248 6811 6306 6817
rect 6380 6712 6408 6820
rect 6524 6817 6536 6851
rect 6524 6811 6552 6817
rect 6546 6808 6552 6811
rect 6604 6808 6610 6860
rect 6822 6857 6828 6860
rect 6800 6851 6828 6857
rect 6800 6817 6812 6851
rect 6800 6811 6828 6817
rect 6822 6808 6828 6811
rect 6880 6808 6886 6860
rect 6932 6848 6960 6944
rect 7190 6876 7196 6928
rect 7248 6916 7254 6928
rect 7248 6888 8156 6916
rect 7248 6876 7254 6888
rect 7466 6857 7472 6860
rect 7044 6851 7102 6857
rect 7044 6848 7056 6851
rect 6932 6820 7056 6848
rect 7044 6817 7056 6820
rect 7090 6817 7102 6851
rect 7044 6811 7102 6817
rect 7434 6851 7472 6857
rect 7434 6817 7446 6851
rect 7434 6811 7472 6817
rect 7466 6808 7472 6811
rect 7524 6808 7530 6860
rect 7852 6857 7880 6888
rect 7561 6851 7619 6857
rect 7561 6817 7573 6851
rect 7607 6817 7619 6851
rect 7561 6811 7619 6817
rect 7837 6851 7895 6857
rect 7837 6817 7849 6851
rect 7883 6817 7895 6851
rect 7837 6811 7895 6817
rect 7576 6780 7604 6811
rect 7926 6808 7932 6860
rect 7984 6808 7990 6860
rect 8128 6857 8156 6888
rect 8220 6888 8616 6916
rect 8220 6860 8248 6888
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6817 8171 6851
rect 8113 6811 8171 6817
rect 8202 6808 8208 6860
rect 8260 6808 8266 6860
rect 8478 6808 8484 6860
rect 8536 6808 8542 6860
rect 8588 6857 8616 6888
rect 8662 6876 8668 6928
rect 8720 6876 8726 6928
rect 8754 6876 8760 6928
rect 8812 6916 8818 6928
rect 9692 6916 9720 6944
rect 8812 6888 9536 6916
rect 8812 6876 8818 6888
rect 8573 6851 8631 6857
rect 8573 6817 8585 6851
rect 8619 6817 8631 6851
rect 8680 6847 8708 6876
rect 8573 6811 8631 6817
rect 8665 6841 8723 6847
rect 7944 6780 7972 6808
rect 8665 6807 8677 6841
rect 8711 6807 8723 6841
rect 8846 6808 8852 6860
rect 8904 6808 8910 6860
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 9508 6857 9536 6888
rect 9600 6888 9720 6916
rect 10520 6916 10548 6944
rect 11149 6919 11207 6925
rect 11149 6916 11161 6919
rect 10520 6888 11161 6916
rect 9600 6857 9628 6888
rect 11149 6885 11161 6888
rect 11195 6885 11207 6919
rect 11149 6879 11207 6885
rect 11330 6876 11336 6928
rect 11388 6876 11394 6928
rect 11698 6876 11704 6928
rect 11756 6916 11762 6928
rect 14568 6916 14596 6944
rect 15948 6916 15976 6956
rect 16577 6953 16589 6956
rect 16623 6953 16635 6987
rect 16577 6947 16635 6953
rect 16758 6944 16764 6996
rect 16816 6944 16822 6996
rect 18414 6944 18420 6996
rect 18472 6984 18478 6996
rect 18874 6984 18880 6996
rect 18472 6956 18880 6984
rect 18472 6944 18478 6956
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 19521 6987 19579 6993
rect 19521 6953 19533 6987
rect 19567 6984 19579 6987
rect 19886 6984 19892 6996
rect 19567 6956 19892 6984
rect 19567 6953 19579 6956
rect 19521 6947 19579 6953
rect 19886 6944 19892 6956
rect 19944 6944 19950 6996
rect 20162 6944 20168 6996
rect 20220 6944 20226 6996
rect 20990 6944 20996 6996
rect 21048 6944 21054 6996
rect 21082 6944 21088 6996
rect 21140 6984 21146 6996
rect 21140 6956 22048 6984
rect 21140 6944 21146 6956
rect 11756 6888 11928 6916
rect 14568 6888 15976 6916
rect 11756 6876 11762 6888
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 9272 6820 9321 6848
rect 9272 6808 9278 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 9585 6851 9643 6857
rect 9585 6817 9597 6851
rect 9631 6817 9643 6851
rect 9585 6811 9643 6817
rect 8665 6801 8723 6807
rect 8386 6780 8392 6792
rect 7576 6752 7880 6780
rect 7944 6752 8392 6780
rect 7374 6712 7380 6724
rect 6380 6684 7380 6712
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 6319 6647 6377 6653
rect 6319 6613 6331 6647
rect 6365 6644 6377 6647
rect 6454 6644 6460 6656
rect 6365 6616 6460 6644
rect 6365 6613 6377 6616
rect 6319 6607 6377 6613
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 6595 6647 6653 6653
rect 6595 6613 6607 6647
rect 6641 6644 6653 6647
rect 6730 6644 6736 6656
rect 6641 6616 6736 6644
rect 6641 6613 6653 6616
rect 6595 6607 6653 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 6871 6647 6929 6653
rect 6871 6613 6883 6647
rect 6917 6644 6929 6647
rect 7006 6644 7012 6656
rect 6917 6616 7012 6644
rect 6917 6613 6929 6616
rect 6871 6607 6929 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7190 6653 7196 6656
rect 7147 6647 7196 6653
rect 7147 6613 7159 6647
rect 7193 6613 7196 6647
rect 7147 6607 7196 6613
rect 7190 6604 7196 6607
rect 7248 6604 7254 6656
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7340 6616 7757 6644
rect 7340 6604 7346 6616
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 7852 6644 7880 6752
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 8754 6740 8760 6792
rect 8812 6740 8818 6792
rect 9324 6780 9352 6811
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 10505 6851 10563 6857
rect 10505 6848 10517 6851
rect 10468 6820 10517 6848
rect 10468 6808 10474 6820
rect 10505 6817 10517 6820
rect 10551 6817 10563 6851
rect 10505 6811 10563 6817
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 10689 6851 10747 6857
rect 10689 6817 10701 6851
rect 10735 6848 10747 6851
rect 11241 6851 11299 6857
rect 11241 6848 11253 6851
rect 10735 6820 11253 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 9324 6752 10097 6780
rect 7929 6715 7987 6721
rect 7929 6681 7941 6715
rect 7975 6712 7987 6715
rect 9582 6712 9588 6724
rect 7975 6684 9588 6712
rect 7975 6681 7987 6684
rect 7929 6675 7987 6681
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 9766 6672 9772 6724
rect 9824 6672 9830 6724
rect 10069 6712 10097 6752
rect 10134 6740 10140 6792
rect 10192 6740 10198 6792
rect 10612 6724 10640 6811
rect 11164 6792 11192 6820
rect 11241 6817 11253 6820
rect 11287 6817 11299 6851
rect 11348 6847 11376 6876
rect 11241 6811 11299 6817
rect 11333 6841 11391 6847
rect 11333 6807 11345 6841
rect 11379 6807 11391 6841
rect 11422 6808 11428 6860
rect 11480 6808 11486 6860
rect 11900 6857 11928 6888
rect 16206 6876 16212 6928
rect 16264 6876 16270 6928
rect 16776 6916 16804 6944
rect 16684 6888 16804 6916
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 11532 6820 11621 6848
rect 11333 6801 11391 6807
rect 11146 6740 11152 6792
rect 11204 6740 11210 6792
rect 11532 6724 11560 6820
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 11885 6851 11943 6857
rect 11885 6817 11897 6851
rect 11931 6848 11943 6851
rect 12250 6848 12256 6860
rect 11931 6820 12256 6848
rect 11931 6817 11943 6820
rect 11885 6811 11943 6817
rect 12250 6808 12256 6820
rect 12308 6848 12314 6860
rect 12345 6851 12403 6857
rect 12345 6848 12357 6851
rect 12308 6820 12357 6848
rect 12308 6808 12314 6820
rect 12345 6817 12357 6820
rect 12391 6817 12403 6851
rect 12345 6811 12403 6817
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 12693 6851 12751 6857
rect 12693 6848 12705 6851
rect 12584 6820 12705 6848
rect 12584 6808 12590 6820
rect 12693 6817 12705 6820
rect 12739 6817 12751 6851
rect 12693 6811 12751 6817
rect 14452 6851 14510 6857
rect 14452 6817 14464 6851
rect 14498 6848 14510 6851
rect 14826 6848 14832 6860
rect 14498 6820 14832 6848
rect 14498 6817 14510 6820
rect 14452 6811 14510 6817
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 14918 6808 14924 6860
rect 14976 6848 14982 6860
rect 14976 6820 15424 6848
rect 14976 6808 14982 6820
rect 12437 6783 12495 6789
rect 12437 6780 12449 6783
rect 11624 6752 12449 6780
rect 10594 6712 10600 6724
rect 10069 6684 10600 6712
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 10686 6672 10692 6724
rect 10744 6672 10750 6724
rect 11514 6672 11520 6724
rect 11572 6672 11578 6724
rect 9677 6647 9735 6653
rect 9677 6644 9689 6647
rect 7852 6616 9689 6644
rect 7745 6607 7803 6613
rect 9677 6613 9689 6616
rect 9723 6613 9735 6647
rect 10704 6644 10732 6672
rect 11624 6644 11652 6752
rect 12437 6749 12449 6752
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 13630 6740 13636 6792
rect 13688 6780 13694 6792
rect 14185 6783 14243 6789
rect 14185 6780 14197 6783
rect 13688 6752 14197 6780
rect 13688 6740 13694 6752
rect 14185 6749 14197 6752
rect 14231 6749 14243 6783
rect 14185 6743 14243 6749
rect 12342 6712 12348 6724
rect 11992 6684 12348 6712
rect 11992 6653 12020 6684
rect 12342 6672 12348 6684
rect 12400 6672 12406 6724
rect 15396 6712 15424 6820
rect 15470 6808 15476 6860
rect 15528 6808 15534 6860
rect 15933 6851 15991 6857
rect 15933 6817 15945 6851
rect 15979 6848 15991 6851
rect 16224 6848 16252 6876
rect 16684 6857 16712 6888
rect 17586 6876 17592 6928
rect 17644 6876 17650 6928
rect 19702 6916 19708 6928
rect 18984 6888 19708 6916
rect 15979 6820 16252 6848
rect 16393 6851 16451 6857
rect 15979 6817 15991 6820
rect 15933 6811 15991 6817
rect 16393 6817 16405 6851
rect 16439 6817 16451 6851
rect 16393 6811 16451 6817
rect 16669 6851 16727 6857
rect 16669 6817 16681 6851
rect 16715 6817 16727 6851
rect 16669 6811 16727 6817
rect 15488 6780 15516 6808
rect 16301 6783 16359 6789
rect 16301 6780 16313 6783
rect 15488 6752 16313 6780
rect 16301 6749 16313 6752
rect 16347 6749 16359 6783
rect 16301 6743 16359 6749
rect 16408 6780 16436 6811
rect 16758 6808 16764 6860
rect 16816 6848 16822 6860
rect 16945 6851 17003 6857
rect 16945 6848 16957 6851
rect 16816 6820 16957 6848
rect 16816 6808 16822 6820
rect 16945 6817 16957 6820
rect 16991 6848 17003 6851
rect 17604 6848 17632 6876
rect 18690 6848 18696 6860
rect 16991 6820 17632 6848
rect 17788 6820 18696 6848
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17788 6780 17816 6820
rect 18690 6808 18696 6820
rect 18748 6848 18754 6860
rect 18984 6857 19012 6888
rect 19702 6876 19708 6888
rect 19760 6876 19766 6928
rect 20180 6916 20208 6944
rect 21008 6916 21036 6944
rect 22020 6916 22048 6956
rect 23934 6944 23940 6996
rect 23992 6984 23998 6996
rect 24578 6984 24584 6996
rect 23992 6956 24584 6984
rect 23992 6944 23998 6956
rect 24578 6944 24584 6956
rect 24636 6944 24642 6996
rect 24857 6987 24915 6993
rect 24857 6953 24869 6987
rect 24903 6984 24915 6987
rect 25498 6984 25504 6996
rect 24903 6956 25504 6984
rect 24903 6953 24915 6956
rect 24857 6947 24915 6953
rect 25498 6944 25504 6956
rect 25556 6944 25562 6996
rect 24026 6916 24032 6928
rect 20088 6888 20208 6916
rect 20824 6888 21036 6916
rect 21284 6888 21956 6916
rect 22020 6888 23152 6916
rect 18969 6851 19027 6857
rect 18969 6848 18981 6851
rect 18748 6820 18981 6848
rect 18748 6808 18754 6820
rect 18969 6817 18981 6820
rect 19015 6817 19027 6851
rect 18969 6811 19027 6817
rect 19061 6851 19119 6857
rect 19061 6817 19073 6851
rect 19107 6817 19119 6851
rect 19061 6811 19119 6817
rect 16408 6752 17816 6780
rect 16408 6712 16436 6752
rect 17862 6740 17868 6792
rect 17920 6740 17926 6792
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 19076 6780 19104 6811
rect 19334 6808 19340 6860
rect 19392 6808 19398 6860
rect 20088 6857 20116 6888
rect 19521 6851 19579 6857
rect 19521 6817 19533 6851
rect 19567 6817 19579 6851
rect 19521 6811 19579 6817
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 20073 6851 20131 6857
rect 19843 6820 20024 6848
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 18840 6752 19104 6780
rect 19153 6783 19211 6789
rect 18840 6740 18846 6752
rect 19153 6749 19165 6783
rect 19199 6780 19211 6783
rect 19536 6780 19564 6811
rect 19199 6752 19564 6780
rect 19996 6780 20024 6820
rect 20073 6817 20085 6851
rect 20119 6817 20131 6851
rect 20073 6811 20131 6817
rect 20165 6851 20223 6857
rect 20165 6817 20177 6851
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 20180 6780 20208 6811
rect 20438 6808 20444 6860
rect 20496 6808 20502 6860
rect 20625 6851 20683 6857
rect 20625 6817 20637 6851
rect 20671 6848 20683 6851
rect 20824 6848 20852 6888
rect 21284 6860 21312 6888
rect 21928 6860 21956 6888
rect 20671 6820 20852 6848
rect 20901 6851 20959 6857
rect 20671 6817 20683 6820
rect 20625 6811 20683 6817
rect 20901 6817 20913 6851
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 19996 6752 20208 6780
rect 19199 6749 19211 6752
rect 19153 6743 19211 6749
rect 15396 6684 16436 6712
rect 17880 6712 17908 6740
rect 18233 6715 18291 6721
rect 18233 6712 18245 6715
rect 17880 6684 18245 6712
rect 18233 6681 18245 6684
rect 18279 6681 18291 6715
rect 19610 6712 19616 6724
rect 18233 6675 18291 6681
rect 18340 6684 19616 6712
rect 10704 6616 11652 6644
rect 11977 6647 12035 6653
rect 9677 6607 9735 6613
rect 11977 6613 11989 6647
rect 12023 6613 12035 6647
rect 11977 6607 12035 6613
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 13170 6644 13176 6656
rect 12308 6616 13176 6644
rect 12308 6604 12314 6616
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 13817 6647 13875 6653
rect 13817 6644 13829 6647
rect 13780 6616 13829 6644
rect 13780 6604 13786 6616
rect 13817 6613 13829 6616
rect 13863 6613 13875 6647
rect 13817 6607 13875 6613
rect 15562 6604 15568 6656
rect 15620 6604 15626 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18340 6644 18368 6684
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 19996 6721 20024 6752
rect 20530 6740 20536 6792
rect 20588 6780 20594 6792
rect 20916 6780 20944 6811
rect 21266 6808 21272 6860
rect 21324 6808 21330 6860
rect 21536 6851 21594 6857
rect 21536 6817 21548 6851
rect 21582 6848 21594 6851
rect 21818 6848 21824 6860
rect 21582 6820 21824 6848
rect 21582 6817 21594 6820
rect 21536 6811 21594 6817
rect 21818 6808 21824 6820
rect 21876 6808 21882 6860
rect 21910 6808 21916 6860
rect 21968 6808 21974 6860
rect 23124 6857 23152 6888
rect 23492 6888 24032 6916
rect 23017 6851 23075 6857
rect 23017 6848 23029 6851
rect 22388 6820 23029 6848
rect 22388 6792 22416 6820
rect 23017 6817 23029 6820
rect 23063 6817 23075 6851
rect 23017 6811 23075 6817
rect 23109 6851 23167 6857
rect 23109 6817 23121 6851
rect 23155 6817 23167 6851
rect 23492 6848 23520 6888
rect 24026 6876 24032 6888
rect 24084 6916 24090 6928
rect 25222 6916 25228 6928
rect 24084 6888 25228 6916
rect 24084 6876 24090 6888
rect 23109 6811 23167 6817
rect 23216 6820 23520 6848
rect 20588 6752 20944 6780
rect 20588 6740 20594 6752
rect 22370 6740 22376 6792
rect 22428 6740 22434 6792
rect 23032 6780 23060 6811
rect 23216 6780 23244 6820
rect 23566 6808 23572 6860
rect 23624 6808 23630 6860
rect 23658 6808 23664 6860
rect 23716 6808 23722 6860
rect 23937 6851 23995 6857
rect 23937 6817 23949 6851
rect 23983 6817 23995 6851
rect 23937 6811 23995 6817
rect 23032 6752 23244 6780
rect 23290 6740 23296 6792
rect 23348 6780 23354 6792
rect 23952 6780 23980 6811
rect 24210 6808 24216 6860
rect 24268 6808 24274 6860
rect 24305 6851 24363 6857
rect 24305 6817 24317 6851
rect 24351 6848 24363 6851
rect 24394 6848 24400 6860
rect 24351 6820 24400 6848
rect 24351 6817 24363 6820
rect 24305 6811 24363 6817
rect 24394 6808 24400 6820
rect 24452 6808 24458 6860
rect 24486 6808 24492 6860
rect 24544 6808 24550 6860
rect 24673 6851 24731 6857
rect 24673 6817 24685 6851
rect 24719 6817 24731 6851
rect 24673 6811 24731 6817
rect 24765 6851 24823 6857
rect 24765 6817 24777 6851
rect 24811 6848 24823 6851
rect 24872 6848 24900 6888
rect 25222 6876 25228 6888
rect 25280 6876 25286 6928
rect 24811 6820 24900 6848
rect 24811 6817 24823 6820
rect 24765 6811 24823 6817
rect 23348 6752 23980 6780
rect 23348 6740 23354 6752
rect 24118 6740 24124 6792
rect 24176 6780 24182 6792
rect 24688 6780 24716 6811
rect 24176 6752 24716 6780
rect 24176 6740 24182 6752
rect 19981 6715 20039 6721
rect 19981 6681 19993 6715
rect 20027 6712 20039 6715
rect 24029 6715 24087 6721
rect 20027 6684 20944 6712
rect 20027 6681 20039 6684
rect 19981 6675 20039 6681
rect 20916 6656 20944 6684
rect 24029 6681 24041 6715
rect 24075 6712 24087 6715
rect 24946 6712 24952 6724
rect 24075 6684 24952 6712
rect 24075 6681 24087 6684
rect 24029 6675 24087 6681
rect 24946 6672 24952 6684
rect 25004 6672 25010 6724
rect 18012 6616 18368 6644
rect 18012 6604 18018 6616
rect 18690 6604 18696 6656
rect 18748 6644 18754 6656
rect 18877 6647 18935 6653
rect 18877 6644 18889 6647
rect 18748 6616 18889 6644
rect 18748 6604 18754 6616
rect 18877 6613 18889 6616
rect 18923 6613 18935 6647
rect 18877 6607 18935 6613
rect 19518 6604 19524 6656
rect 19576 6644 19582 6656
rect 19705 6647 19763 6653
rect 19705 6644 19717 6647
rect 19576 6616 19717 6644
rect 19576 6604 19582 6616
rect 19705 6613 19717 6616
rect 19751 6613 19763 6647
rect 19705 6607 19763 6613
rect 20257 6647 20315 6653
rect 20257 6613 20269 6647
rect 20303 6644 20315 6647
rect 20533 6647 20591 6653
rect 20533 6644 20545 6647
rect 20303 6616 20545 6644
rect 20303 6613 20315 6616
rect 20257 6607 20315 6613
rect 20533 6613 20545 6616
rect 20579 6613 20591 6647
rect 20533 6607 20591 6613
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 20809 6647 20867 6653
rect 20809 6644 20821 6647
rect 20772 6616 20821 6644
rect 20772 6604 20778 6616
rect 20809 6613 20821 6616
rect 20855 6613 20867 6647
rect 20809 6607 20867 6613
rect 20898 6604 20904 6656
rect 20956 6604 20962 6656
rect 21174 6604 21180 6656
rect 21232 6644 21238 6656
rect 22186 6644 22192 6656
rect 21232 6616 22192 6644
rect 21232 6604 21238 6616
rect 22186 6604 22192 6616
rect 22244 6604 22250 6656
rect 22646 6604 22652 6656
rect 22704 6604 22710 6656
rect 22738 6604 22744 6656
rect 22796 6644 22802 6656
rect 22925 6647 22983 6653
rect 22925 6644 22937 6647
rect 22796 6616 22937 6644
rect 22796 6604 22802 6616
rect 22925 6613 22937 6616
rect 22971 6613 22983 6647
rect 22925 6607 22983 6613
rect 23106 6604 23112 6656
rect 23164 6644 23170 6656
rect 23201 6647 23259 6653
rect 23201 6644 23213 6647
rect 23164 6616 23213 6644
rect 23164 6604 23170 6616
rect 23201 6613 23213 6616
rect 23247 6613 23259 6647
rect 23201 6607 23259 6613
rect 23474 6604 23480 6656
rect 23532 6604 23538 6656
rect 23750 6604 23756 6656
rect 23808 6644 23814 6656
rect 24302 6644 24308 6656
rect 23808 6616 24308 6644
rect 23808 6604 23814 6616
rect 24302 6604 24308 6616
rect 24360 6604 24366 6656
rect 24578 6604 24584 6656
rect 24636 6604 24642 6656
rect 552 6554 31372 6576
rect 552 6502 4250 6554
rect 4302 6502 4314 6554
rect 4366 6502 4378 6554
rect 4430 6502 4442 6554
rect 4494 6502 4506 6554
rect 4558 6502 11955 6554
rect 12007 6502 12019 6554
rect 12071 6502 12083 6554
rect 12135 6502 12147 6554
rect 12199 6502 12211 6554
rect 12263 6502 19660 6554
rect 19712 6502 19724 6554
rect 19776 6502 19788 6554
rect 19840 6502 19852 6554
rect 19904 6502 19916 6554
rect 19968 6502 27365 6554
rect 27417 6502 27429 6554
rect 27481 6502 27493 6554
rect 27545 6502 27557 6554
rect 27609 6502 27621 6554
rect 27673 6502 31372 6554
rect 552 6480 31372 6502
rect 6454 6400 6460 6452
rect 6512 6400 6518 6452
rect 7282 6400 7288 6452
rect 7340 6400 7346 6452
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 8067 6443 8125 6449
rect 8067 6440 8079 6443
rect 7524 6412 8079 6440
rect 7524 6400 7530 6412
rect 8067 6409 8079 6412
rect 8113 6409 8125 6443
rect 8067 6403 8125 6409
rect 8202 6400 8208 6452
rect 8260 6400 8266 6452
rect 8527 6443 8585 6449
rect 8527 6409 8539 6443
rect 8573 6440 8585 6443
rect 10134 6440 10140 6452
rect 8573 6412 10140 6440
rect 8573 6409 8585 6412
rect 8527 6403 8585 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 10284 6412 10517 6440
rect 10284 6400 10290 6412
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 10594 6400 10600 6452
rect 10652 6400 10658 6452
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 11296 6412 12434 6440
rect 11296 6400 11302 6412
rect 6472 6304 6500 6400
rect 7300 6372 7328 6400
rect 8220 6372 8248 6400
rect 9490 6372 9496 6384
rect 7300 6344 8156 6372
rect 8220 6344 9496 6372
rect 8128 6304 8156 6344
rect 9490 6332 9496 6344
rect 9548 6332 9554 6384
rect 9674 6332 9680 6384
rect 9732 6332 9738 6384
rect 9858 6332 9864 6384
rect 9916 6372 9922 6384
rect 9916 6344 10272 6372
rect 9916 6332 9922 6344
rect 10134 6304 10140 6316
rect 6472 6276 7696 6304
rect 8128 6276 8708 6304
rect 7098 6196 7104 6248
rect 7156 6196 7162 6248
rect 7190 6196 7196 6248
rect 7248 6196 7254 6248
rect 7668 6245 7696 6276
rect 7342 6239 7400 6245
rect 7342 6205 7354 6239
rect 7388 6236 7400 6239
rect 7515 6239 7573 6245
rect 7515 6236 7527 6239
rect 7388 6208 7527 6236
rect 7388 6205 7400 6208
rect 7342 6199 7400 6205
rect 7515 6205 7527 6208
rect 7561 6205 7573 6239
rect 7515 6199 7573 6205
rect 7618 6239 7696 6245
rect 7618 6205 7630 6239
rect 7664 6208 7696 6239
rect 7664 6205 7676 6208
rect 7618 6199 7676 6205
rect 7834 6196 7840 6248
rect 7892 6245 7898 6248
rect 7892 6239 7920 6245
rect 7908 6205 7920 6239
rect 7892 6199 7920 6205
rect 7892 6196 7898 6199
rect 8018 6196 8024 6248
rect 8076 6236 8082 6248
rect 8680 6245 8708 6276
rect 8772 6276 9352 6304
rect 8138 6239 8196 6245
rect 8138 6236 8150 6239
rect 8076 6208 8150 6236
rect 8076 6196 8082 6208
rect 8138 6205 8150 6208
rect 8184 6205 8196 6239
rect 8424 6239 8482 6245
rect 8424 6236 8436 6239
rect 8138 6199 8196 6205
rect 8312 6208 8436 6236
rect 7116 6100 7144 6196
rect 7208 6168 7236 6196
rect 8312 6168 8340 6208
rect 8424 6205 8436 6208
rect 8470 6205 8482 6239
rect 8424 6199 8482 6205
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 8665 6199 8723 6205
rect 7208 6140 8340 6168
rect 8570 6128 8576 6180
rect 8628 6168 8634 6180
rect 8772 6168 8800 6276
rect 9324 6248 9352 6276
rect 9416 6276 10140 6304
rect 8849 6239 8907 6245
rect 8849 6205 8861 6239
rect 8895 6236 8907 6239
rect 8895 6208 9260 6236
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 8628 6140 8800 6168
rect 8628 6128 8634 6140
rect 8938 6128 8944 6180
rect 8996 6128 9002 6180
rect 9030 6128 9036 6180
rect 9088 6168 9094 6180
rect 9125 6171 9183 6177
rect 9125 6168 9137 6171
rect 9088 6140 9137 6168
rect 9088 6128 9094 6140
rect 9125 6137 9137 6140
rect 9171 6137 9183 6171
rect 9232 6168 9260 6208
rect 9306 6196 9312 6248
rect 9364 6196 9370 6248
rect 9416 6245 9444 6276
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 9401 6239 9459 6245
rect 9401 6205 9413 6239
rect 9447 6205 9459 6239
rect 9401 6199 9459 6205
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6236 9551 6239
rect 10042 6236 10048 6248
rect 9539 6208 10048 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 10244 6236 10272 6344
rect 10318 6264 10324 6316
rect 10376 6264 10382 6316
rect 10612 6245 10640 6400
rect 12406 6372 12434 6412
rect 12710 6400 12716 6452
rect 12768 6400 12774 6452
rect 16758 6440 16764 6452
rect 15672 6412 16764 6440
rect 12989 6375 13047 6381
rect 12989 6372 13001 6375
rect 12406 6344 13001 6372
rect 12989 6341 13001 6344
rect 13035 6341 13047 6375
rect 12989 6335 13047 6341
rect 13265 6375 13323 6381
rect 13265 6341 13277 6375
rect 13311 6372 13323 6375
rect 15286 6372 15292 6384
rect 13311 6344 15292 6372
rect 13311 6341 13323 6344
rect 13265 6335 13323 6341
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 11054 6304 11060 6316
rect 10744 6276 11060 6304
rect 10744 6264 10750 6276
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 13906 6304 13912 6316
rect 12820 6276 13912 6304
rect 10597 6239 10655 6245
rect 10244 6208 10456 6236
rect 9677 6171 9735 6177
rect 9232 6140 9628 6168
rect 9125 6131 9183 6137
rect 7239 6103 7297 6109
rect 7239 6100 7251 6103
rect 7116 6072 7251 6100
rect 7239 6069 7251 6072
rect 7285 6069 7297 6103
rect 7239 6063 7297 6069
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 7791 6103 7849 6109
rect 7791 6100 7803 6103
rect 7432 6072 7803 6100
rect 7432 6060 7438 6072
rect 7791 6069 7803 6072
rect 7837 6069 7849 6103
rect 7791 6063 7849 6069
rect 8754 6060 8760 6112
rect 8812 6060 8818 6112
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9309 6103 9367 6109
rect 9309 6100 9321 6103
rect 9272 6072 9321 6100
rect 9272 6060 9278 6072
rect 9309 6069 9321 6072
rect 9355 6069 9367 6103
rect 9600 6100 9628 6140
rect 9677 6137 9689 6171
rect 9723 6168 9735 6171
rect 10321 6171 10379 6177
rect 10321 6168 10333 6171
rect 9723 6140 10333 6168
rect 9723 6137 9735 6140
rect 9677 6131 9735 6137
rect 10321 6137 10333 6140
rect 10367 6137 10379 6171
rect 10428 6168 10456 6208
rect 10597 6205 10609 6239
rect 10643 6205 10655 6239
rect 10597 6199 10655 6205
rect 10778 6196 10784 6248
rect 10836 6196 10842 6248
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 12820 6245 12848 6276
rect 13906 6264 13912 6276
rect 13964 6264 13970 6316
rect 12805 6239 12863 6245
rect 11204 6208 12756 6236
rect 11204 6196 11210 6208
rect 10873 6171 10931 6177
rect 10873 6168 10885 6171
rect 10428 6140 10885 6168
rect 10321 6131 10379 6137
rect 10873 6137 10885 6140
rect 10919 6137 10931 6171
rect 10873 6131 10931 6137
rect 11324 6171 11382 6177
rect 11324 6137 11336 6171
rect 11370 6168 11382 6171
rect 11790 6168 11796 6180
rect 11370 6140 11796 6168
rect 11370 6137 11382 6140
rect 11324 6131 11382 6137
rect 11790 6128 11796 6140
rect 11848 6128 11854 6180
rect 12728 6168 12756 6208
rect 12805 6205 12817 6239
rect 12851 6205 12863 6239
rect 12805 6199 12863 6205
rect 13081 6239 13139 6245
rect 13081 6205 13093 6239
rect 13127 6205 13139 6239
rect 13081 6199 13139 6205
rect 13096 6168 13124 6199
rect 13170 6196 13176 6248
rect 13228 6196 13234 6248
rect 13814 6196 13820 6248
rect 13872 6196 13878 6248
rect 15194 6196 15200 6248
rect 15252 6196 15258 6248
rect 15672 6245 15700 6412
rect 16758 6400 16764 6412
rect 16816 6400 16822 6452
rect 17773 6443 17831 6449
rect 17773 6409 17785 6443
rect 17819 6440 17831 6443
rect 18598 6440 18604 6452
rect 17819 6412 18604 6440
rect 17819 6409 17831 6412
rect 17773 6403 17831 6409
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 19058 6400 19064 6452
rect 19116 6400 19122 6452
rect 19334 6400 19340 6452
rect 19392 6400 19398 6452
rect 19518 6400 19524 6452
rect 19576 6400 19582 6452
rect 20254 6400 20260 6452
rect 20312 6440 20318 6452
rect 21177 6443 21235 6449
rect 21177 6440 21189 6443
rect 20312 6412 21189 6440
rect 20312 6400 20318 6412
rect 21177 6409 21189 6412
rect 21223 6409 21235 6443
rect 21177 6403 21235 6409
rect 21726 6400 21732 6452
rect 21784 6400 21790 6452
rect 21818 6400 21824 6452
rect 21876 6400 21882 6452
rect 21910 6400 21916 6452
rect 21968 6440 21974 6452
rect 22557 6443 22615 6449
rect 22557 6440 22569 6443
rect 21968 6412 22569 6440
rect 21968 6400 21974 6412
rect 22557 6409 22569 6412
rect 22603 6409 22615 6443
rect 22557 6403 22615 6409
rect 22833 6443 22891 6449
rect 22833 6409 22845 6443
rect 22879 6440 22891 6443
rect 23658 6440 23664 6452
rect 22879 6412 23664 6440
rect 22879 6409 22891 6412
rect 22833 6403 22891 6409
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 23937 6443 23995 6449
rect 23937 6409 23949 6443
rect 23983 6440 23995 6443
rect 24486 6440 24492 6452
rect 23983 6412 24492 6440
rect 23983 6409 23995 6412
rect 23937 6403 23995 6409
rect 24486 6400 24492 6412
rect 24544 6400 24550 6452
rect 17497 6375 17555 6381
rect 17497 6341 17509 6375
rect 17543 6372 17555 6375
rect 18046 6372 18052 6384
rect 17543 6344 18052 6372
rect 17543 6341 17555 6344
rect 17497 6335 17555 6341
rect 18046 6332 18052 6344
rect 18104 6332 18110 6384
rect 18322 6332 18328 6384
rect 18380 6372 18386 6384
rect 19150 6372 19156 6384
rect 18380 6344 19156 6372
rect 18380 6332 18386 6344
rect 19150 6332 19156 6344
rect 19208 6332 19214 6384
rect 17954 6264 17960 6316
rect 18012 6264 18018 6316
rect 18690 6304 18696 6316
rect 18156 6276 18696 6304
rect 15657 6239 15715 6245
rect 15657 6205 15669 6239
rect 15703 6205 15715 6239
rect 15657 6199 15715 6205
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6205 15899 6239
rect 15841 6199 15899 6205
rect 16117 6239 16175 6245
rect 16117 6205 16129 6239
rect 16163 6236 16175 6239
rect 16850 6236 16856 6248
rect 16163 6208 16856 6236
rect 16163 6205 16175 6208
rect 16117 6199 16175 6205
rect 13725 6171 13783 6177
rect 13725 6168 13737 6171
rect 12728 6140 13124 6168
rect 13188 6140 13737 6168
rect 10594 6100 10600 6112
rect 9600 6072 10600 6100
rect 9309 6063 9367 6069
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 12437 6103 12495 6109
rect 12437 6100 12449 6103
rect 12308 6072 12449 6100
rect 12308 6060 12314 6072
rect 12437 6069 12449 6072
rect 12483 6069 12495 6103
rect 12437 6063 12495 6069
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 13188 6100 13216 6140
rect 13725 6137 13737 6140
rect 13771 6137 13783 6171
rect 13725 6131 13783 6137
rect 13909 6171 13967 6177
rect 13909 6137 13921 6171
rect 13955 6137 13967 6171
rect 15212 6168 15240 6196
rect 15856 6168 15884 6199
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6205 17923 6239
rect 17972 6236 18000 6264
rect 18156 6245 18184 6276
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17972 6208 18061 6236
rect 17865 6199 17923 6205
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 18141 6239 18199 6245
rect 18141 6205 18153 6239
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 15212 6140 15884 6168
rect 15933 6171 15991 6177
rect 13909 6131 13967 6137
rect 15933 6137 15945 6171
rect 15979 6168 15991 6171
rect 16362 6171 16420 6177
rect 16362 6168 16374 6171
rect 15979 6140 16374 6168
rect 15979 6137 15991 6140
rect 15933 6131 15991 6137
rect 16362 6137 16374 6140
rect 16408 6137 16420 6171
rect 17880 6168 17908 6199
rect 18322 6196 18328 6248
rect 18380 6196 18386 6248
rect 18417 6239 18475 6245
rect 18417 6205 18429 6239
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 18340 6168 18368 6196
rect 17880 6140 18368 6168
rect 16362 6131 16420 6137
rect 12676 6072 13216 6100
rect 12676 6060 12682 6072
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 13924 6100 13952 6131
rect 13688 6072 13952 6100
rect 13688 6060 13694 6072
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 15654 6100 15660 6112
rect 15252 6072 15660 6100
rect 15252 6060 15258 6072
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 18432 6100 18460 6199
rect 18874 6196 18880 6248
rect 18932 6196 18938 6248
rect 18969 6239 19027 6245
rect 18969 6205 18981 6239
rect 19015 6230 19027 6239
rect 19150 6236 19156 6248
rect 19076 6230 19156 6236
rect 19015 6208 19156 6230
rect 19015 6205 19104 6208
rect 18969 6202 19104 6205
rect 18969 6199 19027 6202
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 18785 6171 18843 6177
rect 18785 6137 18797 6171
rect 18831 6168 18843 6171
rect 19352 6168 19380 6400
rect 19536 6304 19564 6400
rect 20806 6332 20812 6384
rect 20864 6372 20870 6384
rect 21836 6372 21864 6400
rect 24213 6375 24271 6381
rect 24213 6372 24225 6375
rect 20864 6344 21680 6372
rect 21836 6344 24225 6372
rect 20864 6332 20870 6344
rect 21266 6304 21272 6316
rect 19444 6276 19564 6304
rect 20824 6276 21272 6304
rect 19444 6245 19472 6276
rect 19429 6239 19487 6245
rect 19429 6205 19441 6239
rect 19475 6205 19487 6239
rect 19429 6199 19487 6205
rect 19521 6239 19579 6245
rect 19521 6205 19533 6239
rect 19567 6236 19579 6239
rect 20824 6236 20852 6276
rect 21266 6264 21272 6276
rect 21324 6264 21330 6316
rect 21652 6304 21680 6344
rect 24213 6341 24225 6344
rect 24259 6341 24271 6375
rect 24213 6335 24271 6341
rect 23750 6304 23756 6316
rect 21652 6276 23756 6304
rect 19567 6208 20852 6236
rect 19567 6205 19579 6208
rect 19521 6199 19579 6205
rect 20898 6196 20904 6248
rect 20956 6236 20962 6248
rect 21652 6245 21680 6276
rect 21085 6239 21143 6245
rect 21085 6236 21097 6239
rect 20956 6208 21097 6236
rect 20956 6196 20962 6208
rect 21085 6205 21097 6208
rect 21131 6205 21143 6239
rect 21085 6199 21143 6205
rect 21545 6239 21603 6245
rect 21545 6205 21557 6239
rect 21591 6205 21603 6239
rect 21545 6199 21603 6205
rect 21637 6239 21695 6245
rect 21637 6205 21649 6239
rect 21683 6205 21695 6239
rect 21637 6199 21695 6205
rect 18831 6140 19380 6168
rect 19788 6171 19846 6177
rect 18831 6137 18843 6140
rect 18785 6131 18843 6137
rect 19788 6137 19800 6171
rect 19834 6168 19846 6171
rect 20070 6168 20076 6180
rect 19834 6140 20076 6168
rect 19834 6137 19846 6140
rect 19788 6131 19846 6137
rect 20070 6128 20076 6140
rect 20128 6128 20134 6180
rect 20346 6128 20352 6180
rect 20404 6128 20410 6180
rect 21266 6168 21272 6180
rect 20916 6140 21272 6168
rect 19242 6100 19248 6112
rect 18432 6072 19248 6100
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 19337 6103 19395 6109
rect 19337 6069 19349 6103
rect 19383 6100 19395 6103
rect 20364 6100 20392 6128
rect 20916 6109 20944 6140
rect 21266 6128 21272 6140
rect 21324 6128 21330 6180
rect 21560 6168 21588 6199
rect 21726 6196 21732 6248
rect 21784 6196 21790 6248
rect 22002 6196 22008 6248
rect 22060 6196 22066 6248
rect 22094 6196 22100 6248
rect 22152 6196 22158 6248
rect 22186 6196 22192 6248
rect 22244 6196 22250 6248
rect 22278 6196 22284 6248
rect 22336 6236 22342 6248
rect 22664 6245 22692 6276
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 23845 6249 23903 6255
rect 22649 6239 22707 6245
rect 22336 6208 22600 6236
rect 22336 6196 22342 6208
rect 21744 6168 21772 6196
rect 21560 6140 21772 6168
rect 19383 6072 20392 6100
rect 20901 6103 20959 6109
rect 19383 6069 19395 6072
rect 19337 6063 19395 6069
rect 20901 6069 20913 6103
rect 20947 6069 20959 6103
rect 20901 6063 20959 6069
rect 21450 6060 21456 6112
rect 21508 6060 21514 6112
rect 22020 6109 22048 6196
rect 22572 6168 22600 6208
rect 22649 6205 22661 6239
rect 22695 6205 22707 6239
rect 22649 6199 22707 6205
rect 22741 6239 22799 6245
rect 22741 6205 22753 6239
rect 22787 6236 22799 6239
rect 22787 6208 22968 6236
rect 22787 6205 22799 6208
rect 22741 6199 22799 6205
rect 22940 6180 22968 6208
rect 23198 6196 23204 6248
rect 23256 6196 23262 6248
rect 23293 6239 23351 6245
rect 23293 6205 23305 6239
rect 23339 6205 23351 6239
rect 23293 6199 23351 6205
rect 22922 6168 22928 6180
rect 22572 6140 22928 6168
rect 22922 6128 22928 6140
rect 22980 6128 22986 6180
rect 23014 6128 23020 6180
rect 23072 6168 23078 6180
rect 23308 6168 23336 6199
rect 23382 6196 23388 6248
rect 23440 6236 23446 6248
rect 23477 6239 23535 6245
rect 23477 6236 23489 6239
rect 23440 6208 23489 6236
rect 23440 6196 23446 6208
rect 23477 6205 23489 6208
rect 23523 6205 23535 6239
rect 23845 6215 23857 6249
rect 23891 6215 23903 6249
rect 23845 6209 23903 6215
rect 24305 6239 24363 6245
rect 23477 6199 23535 6205
rect 23860 6180 23888 6209
rect 24305 6205 24317 6239
rect 24351 6236 24363 6239
rect 25314 6236 25320 6248
rect 24351 6208 25320 6236
rect 24351 6205 24363 6208
rect 24305 6199 24363 6205
rect 25314 6196 25320 6208
rect 25372 6196 25378 6248
rect 23072 6140 23336 6168
rect 23072 6128 23078 6140
rect 23842 6128 23848 6180
rect 23900 6128 23906 6180
rect 22005 6103 22063 6109
rect 22005 6069 22017 6103
rect 22051 6069 22063 6103
rect 22005 6063 22063 6069
rect 22278 6060 22284 6112
rect 22336 6060 22342 6112
rect 22830 6060 22836 6112
rect 22888 6100 22894 6112
rect 23109 6103 23167 6109
rect 23109 6100 23121 6103
rect 22888 6072 23121 6100
rect 22888 6060 22894 6072
rect 23109 6069 23121 6072
rect 23155 6069 23167 6103
rect 23109 6063 23167 6069
rect 23290 6060 23296 6112
rect 23348 6060 23354 6112
rect 552 6010 31531 6032
rect 552 5958 8102 6010
rect 8154 5958 8166 6010
rect 8218 5958 8230 6010
rect 8282 5958 8294 6010
rect 8346 5958 8358 6010
rect 8410 5958 15807 6010
rect 15859 5958 15871 6010
rect 15923 5958 15935 6010
rect 15987 5958 15999 6010
rect 16051 5958 16063 6010
rect 16115 5958 23512 6010
rect 23564 5958 23576 6010
rect 23628 5958 23640 6010
rect 23692 5958 23704 6010
rect 23756 5958 23768 6010
rect 23820 5958 31217 6010
rect 31269 5958 31281 6010
rect 31333 5958 31345 6010
rect 31397 5958 31409 6010
rect 31461 5958 31473 6010
rect 31525 5958 31531 6010
rect 552 5936 31531 5958
rect 6730 5856 6736 5908
rect 6788 5856 6794 5908
rect 7006 5856 7012 5908
rect 7064 5856 7070 5908
rect 7834 5905 7840 5908
rect 7791 5899 7840 5905
rect 7791 5865 7803 5899
rect 7837 5865 7840 5899
rect 7791 5859 7840 5865
rect 7834 5856 7840 5859
rect 7892 5856 7898 5908
rect 8478 5856 8484 5908
rect 8536 5856 8542 5908
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 8938 5896 8944 5908
rect 8619 5868 8944 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 6748 5760 6776 5856
rect 7024 5828 7052 5856
rect 8496 5828 8524 5856
rect 9140 5828 9168 5859
rect 9214 5856 9220 5908
rect 9272 5856 9278 5908
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 9548 5868 9674 5896
rect 9548 5856 9554 5868
rect 7024 5800 7855 5828
rect 8496 5800 9168 5828
rect 7688 5763 7746 5769
rect 7688 5760 7700 5763
rect 6748 5732 7700 5760
rect 7688 5729 7700 5732
rect 7734 5729 7746 5763
rect 7827 5760 7855 5800
rect 8046 5763 8104 5769
rect 8046 5760 8058 5763
rect 7827 5732 8058 5760
rect 7688 5723 7746 5729
rect 8046 5729 8058 5732
rect 8092 5729 8104 5763
rect 8046 5723 8104 5729
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5760 8447 5763
rect 8481 5763 8539 5769
rect 8481 5760 8493 5763
rect 8435 5732 8493 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 8481 5729 8493 5732
rect 8527 5760 8539 5763
rect 8570 5760 8576 5772
rect 8527 5732 8576 5760
rect 8527 5729 8539 5732
rect 8481 5723 8539 5729
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 8874 5763 8932 5769
rect 8874 5760 8886 5763
rect 8680 5732 8886 5760
rect 8680 5704 8708 5732
rect 8874 5729 8886 5732
rect 8920 5760 8932 5763
rect 9030 5760 9036 5772
rect 8920 5732 9036 5760
rect 8920 5729 8932 5732
rect 8874 5723 8932 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 6546 5652 6552 5704
rect 6604 5652 6610 5704
rect 6822 5652 6828 5704
rect 6880 5692 6886 5704
rect 6880 5664 8156 5692
rect 6880 5652 6886 5664
rect 6564 5624 6592 5652
rect 7975 5627 8033 5633
rect 7975 5624 7987 5627
rect 6564 5596 7987 5624
rect 7975 5593 7987 5596
rect 8021 5593 8033 5627
rect 7975 5587 8033 5593
rect 8128 5556 8156 5664
rect 8662 5652 8668 5704
rect 8720 5652 8726 5704
rect 9140 5692 9168 5800
rect 9232 5769 9260 5856
rect 9646 5828 9674 5868
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 10781 5899 10839 5905
rect 10781 5896 10793 5899
rect 10100 5868 10793 5896
rect 10100 5856 10106 5868
rect 10781 5865 10793 5868
rect 10827 5865 10839 5899
rect 10781 5859 10839 5865
rect 10796 5828 10824 5859
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 13814 5896 13820 5908
rect 12400 5868 13820 5896
rect 12400 5856 12406 5868
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 14458 5896 14464 5908
rect 14415 5868 14464 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 14458 5856 14464 5868
rect 14516 5896 14522 5908
rect 14516 5868 14596 5896
rect 14516 5856 14522 5868
rect 12538 5831 12596 5837
rect 12538 5828 12550 5831
rect 9646 5800 10732 5828
rect 10796 5800 12550 5828
rect 9674 5769 9680 5772
rect 9217 5763 9275 5769
rect 9217 5729 9229 5763
rect 9263 5729 9275 5763
rect 9668 5760 9680 5769
rect 9635 5732 9680 5760
rect 9217 5723 9275 5729
rect 9668 5723 9680 5732
rect 9674 5720 9680 5723
rect 9732 5720 9738 5772
rect 10704 5760 10732 5800
rect 12538 5797 12550 5800
rect 12584 5797 12596 5831
rect 13630 5828 13636 5840
rect 12538 5791 12596 5797
rect 12820 5800 13636 5828
rect 11057 5763 11115 5769
rect 11057 5760 11069 5763
rect 10704 5732 11069 5760
rect 11057 5729 11069 5732
rect 11103 5760 11115 5763
rect 11330 5760 11336 5772
rect 11103 5732 11336 5760
rect 11103 5729 11115 5732
rect 11057 5723 11115 5729
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 12820 5704 12848 5800
rect 13630 5788 13636 5800
rect 13688 5828 13694 5840
rect 14568 5828 14596 5868
rect 17862 5856 17868 5908
rect 17920 5856 17926 5908
rect 18782 5856 18788 5908
rect 18840 5856 18846 5908
rect 19337 5899 19395 5905
rect 19337 5865 19349 5899
rect 19383 5896 19395 5899
rect 20438 5896 20444 5908
rect 19383 5868 20444 5896
rect 19383 5865 19395 5868
rect 19337 5859 19395 5865
rect 20438 5856 20444 5868
rect 20496 5856 20502 5908
rect 20530 5856 20536 5908
rect 20588 5896 20594 5908
rect 21910 5896 21916 5908
rect 20588 5868 21916 5896
rect 20588 5856 20594 5868
rect 21910 5856 21916 5868
rect 21968 5856 21974 5908
rect 22554 5856 22560 5908
rect 22612 5856 22618 5908
rect 22741 5899 22799 5905
rect 22741 5865 22753 5899
rect 22787 5896 22799 5899
rect 23290 5896 23296 5908
rect 22787 5868 23296 5896
rect 22787 5865 22799 5868
rect 22741 5859 22799 5865
rect 23290 5856 23296 5868
rect 23348 5856 23354 5908
rect 24118 5856 24124 5908
rect 24176 5856 24182 5908
rect 14706 5831 14764 5837
rect 14706 5828 14718 5831
rect 13688 5800 14504 5828
rect 14568 5800 14718 5828
rect 13688 5788 13694 5800
rect 13256 5763 13314 5769
rect 13256 5729 13268 5763
rect 13302 5760 13314 5763
rect 13538 5760 13544 5772
rect 13302 5732 13544 5760
rect 13302 5729 13314 5732
rect 13256 5723 13314 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 14476 5769 14504 5800
rect 14706 5797 14718 5800
rect 14752 5797 14764 5831
rect 14706 5791 14764 5797
rect 14461 5763 14519 5769
rect 14461 5729 14473 5763
rect 14507 5729 14519 5763
rect 15010 5760 15016 5772
rect 14461 5723 14519 5729
rect 14568 5732 15016 5760
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 9140 5664 9413 5692
rect 9401 5661 9413 5664
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 11149 5695 11207 5701
rect 11149 5692 11161 5695
rect 10928 5664 11161 5692
rect 10928 5652 10934 5664
rect 11149 5661 11161 5664
rect 11195 5692 11207 5695
rect 11422 5692 11428 5704
rect 11195 5664 11428 5692
rect 11195 5661 11207 5664
rect 11149 5655 11207 5661
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 12802 5652 12808 5704
rect 12860 5652 12866 5704
rect 12989 5695 13047 5701
rect 12989 5661 13001 5695
rect 13035 5661 13047 5695
rect 14568 5692 14596 5732
rect 15010 5720 15016 5732
rect 15068 5760 15074 5772
rect 15068 5732 15608 5760
rect 15068 5720 15074 5732
rect 12989 5655 13047 5661
rect 14016 5664 14596 5692
rect 15580 5692 15608 5732
rect 15654 5720 15660 5772
rect 15712 5760 15718 5772
rect 16373 5763 16431 5769
rect 16373 5760 16385 5763
rect 15712 5732 16385 5760
rect 15712 5720 15718 5732
rect 16373 5729 16385 5732
rect 16419 5729 16431 5763
rect 16373 5723 16431 5729
rect 17681 5763 17739 5769
rect 17681 5729 17693 5763
rect 17727 5760 17739 5763
rect 17880 5760 17908 5856
rect 17727 5732 17908 5760
rect 17948 5763 18006 5769
rect 17727 5729 17739 5732
rect 17681 5723 17739 5729
rect 17948 5729 17960 5763
rect 17994 5760 18006 5763
rect 18800 5760 18828 5856
rect 20714 5828 20720 5840
rect 20548 5800 20720 5828
rect 19150 5760 19156 5772
rect 17994 5732 18736 5760
rect 18800 5732 19156 5760
rect 17994 5729 18006 5732
rect 17948 5723 18006 5729
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 15580 5664 16129 5692
rect 8297 5627 8355 5633
rect 8297 5593 8309 5627
rect 8343 5624 8355 5627
rect 8343 5596 9444 5624
rect 8343 5593 8355 5596
rect 8297 5587 8355 5593
rect 8803 5559 8861 5565
rect 8803 5556 8815 5559
rect 8128 5528 8815 5556
rect 8803 5525 8815 5528
rect 8849 5525 8861 5559
rect 9416 5556 9444 5596
rect 10962 5584 10968 5636
rect 11020 5624 11026 5636
rect 11020 5596 11468 5624
rect 11020 5584 11026 5596
rect 9674 5556 9680 5568
rect 9416 5528 9680 5556
rect 8803 5519 8861 5525
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 11440 5565 11468 5596
rect 11425 5559 11483 5565
rect 11425 5525 11437 5559
rect 11471 5525 11483 5559
rect 13004 5556 13032 5655
rect 14016 5556 14044 5664
rect 16117 5661 16129 5664
rect 16163 5661 16175 5695
rect 18708 5692 18736 5732
rect 19150 5720 19156 5732
rect 19208 5760 19214 5772
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 19208 5732 19257 5760
rect 19208 5720 19214 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 19521 5763 19579 5769
rect 19521 5760 19533 5763
rect 19392 5732 19533 5760
rect 19392 5720 19398 5732
rect 19521 5729 19533 5732
rect 19567 5729 19579 5763
rect 19521 5723 19579 5729
rect 19981 5763 20039 5769
rect 19981 5729 19993 5763
rect 20027 5760 20039 5763
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 20027 5732 20177 5760
rect 20027 5729 20039 5732
rect 19981 5723 20039 5729
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 20257 5763 20315 5769
rect 20257 5729 20269 5763
rect 20303 5760 20315 5763
rect 20346 5760 20352 5772
rect 20303 5732 20352 5760
rect 20303 5729 20315 5732
rect 20257 5723 20315 5729
rect 19613 5695 19671 5701
rect 19613 5692 19625 5695
rect 18708 5664 19625 5692
rect 16117 5655 16175 5661
rect 19613 5661 19625 5664
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 20070 5652 20076 5704
rect 20128 5692 20134 5704
rect 20272 5692 20300 5723
rect 20346 5720 20352 5732
rect 20404 5720 20410 5772
rect 20548 5769 20576 5800
rect 20714 5788 20720 5800
rect 20772 5788 20778 5840
rect 21358 5788 21364 5840
rect 21416 5788 21422 5840
rect 22572 5828 22600 5856
rect 22296 5800 22600 5828
rect 23017 5831 23075 5837
rect 20533 5763 20591 5769
rect 20533 5729 20545 5763
rect 20579 5729 20591 5763
rect 20533 5723 20591 5729
rect 20625 5763 20683 5769
rect 20625 5729 20637 5763
rect 20671 5729 20683 5763
rect 20625 5723 20683 5729
rect 20128 5664 20300 5692
rect 20128 5652 20134 5664
rect 19058 5584 19064 5636
rect 19116 5584 19122 5636
rect 19242 5584 19248 5636
rect 19300 5624 19306 5636
rect 20640 5624 20668 5723
rect 20806 5720 20812 5772
rect 20864 5720 20870 5772
rect 20898 5720 20904 5772
rect 20956 5760 20962 5772
rect 21085 5763 21143 5769
rect 21085 5760 21097 5763
rect 20956 5732 21097 5760
rect 20956 5720 20962 5732
rect 21085 5729 21097 5732
rect 21131 5729 21143 5763
rect 21085 5723 21143 5729
rect 21450 5720 21456 5772
rect 21508 5720 21514 5772
rect 21634 5720 21640 5772
rect 21692 5720 21698 5772
rect 21729 5763 21787 5769
rect 21729 5729 21741 5763
rect 21775 5760 21787 5763
rect 21818 5760 21824 5772
rect 21775 5732 21824 5760
rect 21775 5729 21787 5732
rect 21729 5723 21787 5729
rect 21818 5720 21824 5732
rect 21876 5720 21882 5772
rect 21910 5720 21916 5772
rect 21968 5760 21974 5772
rect 22296 5769 22324 5800
rect 23017 5797 23029 5831
rect 23063 5828 23075 5831
rect 24136 5828 24164 5856
rect 23063 5800 24164 5828
rect 23063 5797 23075 5800
rect 23017 5791 23075 5797
rect 22005 5763 22063 5769
rect 22005 5760 22017 5763
rect 21968 5732 22017 5760
rect 21968 5720 21974 5732
rect 22005 5729 22017 5732
rect 22051 5729 22063 5763
rect 22005 5723 22063 5729
rect 22281 5763 22339 5769
rect 22281 5729 22293 5763
rect 22327 5729 22339 5763
rect 22281 5723 22339 5729
rect 22373 5763 22431 5769
rect 22373 5729 22385 5763
rect 22419 5729 22431 5763
rect 22373 5723 22431 5729
rect 20714 5652 20720 5704
rect 20772 5692 20778 5704
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 20772 5664 21005 5692
rect 20772 5652 20778 5664
rect 20993 5661 21005 5664
rect 21039 5661 21051 5695
rect 20993 5655 21051 5661
rect 21358 5652 21364 5704
rect 21416 5692 21422 5704
rect 22388 5692 22416 5723
rect 22462 5720 22468 5772
rect 22520 5720 22526 5772
rect 22649 5763 22707 5769
rect 22649 5729 22661 5763
rect 22695 5729 22707 5763
rect 22649 5723 22707 5729
rect 23109 5763 23167 5769
rect 23109 5729 23121 5763
rect 23155 5760 23167 5763
rect 23385 5763 23443 5769
rect 23155 5732 23336 5760
rect 23155 5729 23167 5732
rect 23109 5723 23167 5729
rect 21416 5664 22416 5692
rect 21416 5652 21422 5664
rect 19300 5596 20668 5624
rect 19300 5584 19306 5596
rect 21542 5584 21548 5636
rect 21600 5624 21606 5636
rect 22370 5624 22376 5636
rect 21600 5596 22376 5624
rect 21600 5584 21606 5596
rect 22370 5584 22376 5596
rect 22428 5624 22434 5636
rect 22664 5624 22692 5723
rect 23308 5692 23336 5732
rect 23385 5729 23397 5763
rect 23431 5760 23443 5763
rect 26142 5760 26148 5772
rect 23431 5732 26148 5760
rect 23431 5729 23443 5732
rect 23385 5723 23443 5729
rect 26142 5720 26148 5732
rect 26200 5720 26206 5772
rect 25866 5692 25872 5704
rect 23308 5664 25872 5692
rect 25866 5652 25872 5664
rect 25924 5652 25930 5704
rect 22428 5596 22692 5624
rect 22428 5584 22434 5596
rect 22922 5584 22928 5636
rect 22980 5624 22986 5636
rect 23293 5627 23351 5633
rect 23293 5624 23305 5627
rect 22980 5596 23305 5624
rect 22980 5584 22986 5596
rect 23293 5593 23305 5596
rect 23339 5624 23351 5627
rect 24210 5624 24216 5636
rect 23339 5596 24216 5624
rect 23339 5593 23351 5596
rect 23293 5587 23351 5593
rect 24210 5584 24216 5596
rect 24268 5584 24274 5636
rect 13004 5528 14044 5556
rect 15841 5559 15899 5565
rect 11425 5519 11483 5525
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 16298 5556 16304 5568
rect 15887 5528 16304 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 17310 5516 17316 5568
rect 17368 5556 17374 5568
rect 17497 5559 17555 5565
rect 17497 5556 17509 5559
rect 17368 5528 17509 5556
rect 17368 5516 17374 5528
rect 17497 5525 17509 5528
rect 17543 5525 17555 5559
rect 17497 5519 17555 5525
rect 19889 5559 19947 5565
rect 19889 5525 19901 5559
rect 19935 5556 19947 5559
rect 20441 5559 20499 5565
rect 20441 5556 20453 5559
rect 19935 5528 20453 5556
rect 19935 5525 19947 5528
rect 19889 5519 19947 5525
rect 20441 5525 20453 5528
rect 20487 5525 20499 5559
rect 20441 5519 20499 5525
rect 20530 5516 20536 5568
rect 20588 5556 20594 5568
rect 20717 5559 20775 5565
rect 20717 5556 20729 5559
rect 20588 5528 20729 5556
rect 20588 5516 20594 5528
rect 20717 5525 20729 5528
rect 20763 5525 20775 5559
rect 20717 5519 20775 5525
rect 21910 5516 21916 5568
rect 21968 5516 21974 5568
rect 22189 5559 22247 5565
rect 22189 5525 22201 5559
rect 22235 5556 22247 5559
rect 24854 5556 24860 5568
rect 22235 5528 24860 5556
rect 22235 5525 22247 5528
rect 22189 5519 22247 5525
rect 24854 5516 24860 5528
rect 24912 5516 24918 5568
rect 552 5466 31372 5488
rect 552 5414 4250 5466
rect 4302 5414 4314 5466
rect 4366 5414 4378 5466
rect 4430 5414 4442 5466
rect 4494 5414 4506 5466
rect 4558 5414 11955 5466
rect 12007 5414 12019 5466
rect 12071 5414 12083 5466
rect 12135 5414 12147 5466
rect 12199 5414 12211 5466
rect 12263 5414 19660 5466
rect 19712 5414 19724 5466
rect 19776 5414 19788 5466
rect 19840 5414 19852 5466
rect 19904 5414 19916 5466
rect 19968 5414 27365 5466
rect 27417 5414 27429 5466
rect 27481 5414 27493 5466
rect 27545 5414 27557 5466
rect 27609 5414 27621 5466
rect 27673 5414 31372 5466
rect 552 5392 31372 5414
rect 9582 5312 9588 5364
rect 9640 5312 9646 5364
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 10137 5355 10195 5361
rect 10137 5352 10149 5355
rect 9732 5324 10149 5352
rect 9732 5312 9738 5324
rect 10137 5321 10149 5324
rect 10183 5321 10195 5355
rect 11054 5352 11060 5364
rect 10137 5315 10195 5321
rect 10888 5324 11060 5352
rect 9600 5284 9628 5312
rect 10689 5287 10747 5293
rect 10689 5284 10701 5287
rect 9600 5256 10701 5284
rect 10689 5253 10701 5256
rect 10735 5253 10747 5287
rect 10689 5247 10747 5253
rect 8036 5188 8524 5216
rect 8036 5157 8064 5188
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5117 8079 5151
rect 8021 5111 8079 5117
rect 8386 5108 8392 5160
rect 8444 5108 8450 5160
rect 8496 5148 8524 5188
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 10888 5225 10916 5324
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 12526 5312 12532 5364
rect 12584 5312 12590 5364
rect 13078 5312 13084 5364
rect 13136 5312 13142 5364
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 15289 5355 15347 5361
rect 14608 5324 15240 5352
rect 14608 5312 14614 5324
rect 15212 5284 15240 5324
rect 15289 5321 15301 5355
rect 15335 5352 15347 5355
rect 15470 5352 15476 5364
rect 15335 5324 15476 5352
rect 15335 5321 15347 5324
rect 15289 5315 15347 5321
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 16301 5355 16359 5361
rect 16301 5321 16313 5355
rect 16347 5352 16359 5355
rect 16669 5355 16727 5361
rect 16669 5352 16681 5355
rect 16347 5324 16681 5352
rect 16347 5321 16359 5324
rect 16301 5315 16359 5321
rect 16669 5321 16681 5324
rect 16715 5321 16727 5355
rect 16669 5315 16727 5321
rect 19242 5312 19248 5364
rect 19300 5312 19306 5364
rect 19334 5312 19340 5364
rect 19392 5312 19398 5364
rect 19521 5355 19579 5361
rect 19521 5321 19533 5355
rect 19567 5352 19579 5355
rect 20530 5352 20536 5364
rect 19567 5324 20536 5352
rect 19567 5321 19579 5324
rect 19521 5315 19579 5321
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 20806 5352 20812 5364
rect 20640 5324 20812 5352
rect 16022 5284 16028 5296
rect 15212 5256 16028 5284
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 18785 5287 18843 5293
rect 18785 5253 18797 5287
rect 18831 5284 18843 5287
rect 19352 5284 19380 5312
rect 18831 5256 19380 5284
rect 19797 5287 19855 5293
rect 18831 5253 18843 5256
rect 18785 5247 18843 5253
rect 19797 5253 19809 5287
rect 19843 5284 19855 5287
rect 20640 5284 20668 5324
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 21450 5312 21456 5364
rect 21508 5312 21514 5364
rect 21729 5355 21787 5361
rect 21729 5321 21741 5355
rect 21775 5352 21787 5355
rect 22002 5352 22008 5364
rect 21775 5324 22008 5352
rect 21775 5321 21787 5324
rect 21729 5315 21787 5321
rect 22002 5312 22008 5324
rect 22060 5312 22066 5364
rect 22281 5355 22339 5361
rect 22281 5321 22293 5355
rect 22327 5352 22339 5355
rect 24578 5352 24584 5364
rect 22327 5324 24584 5352
rect 22327 5321 22339 5324
rect 22281 5315 22339 5321
rect 24578 5312 24584 5324
rect 24636 5312 24642 5364
rect 20898 5284 20904 5296
rect 19843 5256 20668 5284
rect 20824 5256 20904 5284
rect 19843 5253 19855 5256
rect 19797 5247 19855 5253
rect 10873 5219 10931 5225
rect 9456 5188 10640 5216
rect 9456 5176 9462 5188
rect 8496 5120 9996 5148
rect 8634 5083 8692 5089
rect 8634 5080 8646 5083
rect 8220 5052 8646 5080
rect 8220 5021 8248 5052
rect 8634 5049 8646 5052
rect 8680 5049 8692 5083
rect 8634 5043 8692 5049
rect 8205 5015 8263 5021
rect 8205 4981 8217 5015
rect 8251 4981 8263 5015
rect 8205 4975 8263 4981
rect 9766 4972 9772 5024
rect 9824 4972 9830 5024
rect 9968 5021 9996 5120
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10612 5157 10640 5188
rect 10873 5185 10885 5219
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5216 13783 5219
rect 15470 5216 15476 5228
rect 13771 5188 15476 5216
rect 13771 5185 13783 5188
rect 13725 5179 13783 5185
rect 10505 5151 10563 5157
rect 10505 5148 10517 5151
rect 10100 5120 10517 5148
rect 10100 5108 10106 5120
rect 10505 5117 10517 5120
rect 10551 5117 10563 5151
rect 10505 5111 10563 5117
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 10781 5151 10839 5157
rect 10781 5117 10793 5151
rect 10827 5117 10839 5151
rect 10781 5111 10839 5117
rect 10410 5040 10416 5092
rect 10468 5080 10474 5092
rect 10796 5080 10824 5111
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 11572 5120 12449 5148
rect 11572 5108 11578 5120
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 13817 5151 13875 5157
rect 12768 5120 13676 5148
rect 12768 5108 12774 5120
rect 10468 5052 10824 5080
rect 10468 5040 10474 5052
rect 10870 5040 10876 5092
rect 10928 5080 10934 5092
rect 11118 5083 11176 5089
rect 11118 5080 11130 5083
rect 10928 5052 11130 5080
rect 10928 5040 10934 5052
rect 11118 5049 11130 5052
rect 11164 5049 11176 5083
rect 11118 5043 11176 5049
rect 13081 5083 13139 5089
rect 13081 5049 13093 5083
rect 13127 5080 13139 5083
rect 13127 5052 13584 5080
rect 13127 5049 13139 5052
rect 13081 5043 13139 5049
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 4981 10011 5015
rect 9953 4975 10011 4981
rect 10134 4972 10140 5024
rect 10192 4972 10198 5024
rect 11606 4972 11612 5024
rect 11664 5012 11670 5024
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 11664 4984 12265 5012
rect 11664 4972 11670 4984
rect 12253 4981 12265 4984
rect 12299 4981 12311 5015
rect 12253 4975 12311 4981
rect 13262 4972 13268 5024
rect 13320 4972 13326 5024
rect 13556 5021 13584 5052
rect 13541 5015 13599 5021
rect 13541 4981 13553 5015
rect 13587 4981 13599 5015
rect 13648 5012 13676 5120
rect 13817 5117 13829 5151
rect 13863 5117 13875 5151
rect 13817 5111 13875 5117
rect 13832 5080 13860 5111
rect 13906 5108 13912 5160
rect 13964 5108 13970 5160
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14458 5148 14464 5160
rect 14047 5120 14464 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 14568 5157 14596 5188
rect 15470 5176 15476 5188
rect 15528 5216 15534 5228
rect 15528 5188 16160 5216
rect 15528 5176 15534 5188
rect 14553 5151 14611 5157
rect 14553 5117 14565 5151
rect 14599 5117 14611 5151
rect 14553 5111 14611 5117
rect 14918 5108 14924 5160
rect 14976 5108 14982 5160
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5148 15255 5151
rect 15286 5148 15292 5160
rect 15243 5120 15292 5148
rect 15243 5117 15255 5120
rect 15197 5111 15255 5117
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 15436 5120 15577 5148
rect 15436 5108 15442 5120
rect 15565 5117 15577 5120
rect 15611 5117 15623 5151
rect 15565 5111 15623 5117
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 16022 5148 16028 5160
rect 15887 5120 16028 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 16132 5157 16160 5188
rect 16850 5176 16856 5228
rect 16908 5216 16914 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16908 5188 17049 5216
rect 16908 5176 16914 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 20254 5216 20260 5228
rect 17037 5179 17095 5185
rect 19904 5188 20260 5216
rect 17310 5157 17316 5160
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5148 16175 5151
rect 17304 5148 17316 5157
rect 16163 5120 17316 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 17304 5111 17316 5120
rect 17310 5108 17316 5111
rect 17368 5108 17374 5160
rect 19150 5157 19156 5160
rect 18877 5151 18935 5157
rect 18877 5117 18889 5151
rect 18923 5117 18935 5151
rect 19145 5148 19156 5157
rect 19111 5120 19156 5148
rect 18877 5111 18935 5117
rect 19145 5111 19156 5120
rect 14090 5080 14096 5092
rect 13832 5052 14096 5080
rect 14090 5040 14096 5052
rect 14148 5080 14154 5092
rect 14829 5083 14887 5089
rect 14148 5052 14596 5080
rect 14148 5040 14154 5052
rect 14568 5024 14596 5052
rect 14829 5049 14841 5083
rect 14875 5080 14887 5083
rect 15102 5080 15108 5092
rect 14875 5052 15108 5080
rect 14875 5049 14887 5052
rect 14829 5043 14887 5049
rect 15102 5040 15108 5052
rect 15160 5040 15166 5092
rect 15657 5083 15715 5089
rect 15657 5049 15669 5083
rect 15703 5080 15715 5083
rect 16206 5080 16212 5092
rect 15703 5052 16212 5080
rect 15703 5049 15715 5052
rect 15657 5043 15715 5049
rect 16206 5040 16212 5052
rect 16264 5040 16270 5092
rect 16853 5083 16911 5089
rect 16853 5080 16865 5083
rect 16776 5052 16865 5080
rect 16776 5024 16804 5052
rect 16853 5049 16865 5052
rect 16899 5049 16911 5083
rect 18892 5080 18920 5111
rect 19150 5108 19156 5111
rect 19208 5108 19214 5160
rect 19613 5151 19671 5157
rect 19613 5117 19625 5151
rect 19659 5148 19671 5151
rect 19702 5148 19708 5160
rect 19659 5120 19708 5148
rect 19659 5117 19671 5120
rect 19613 5111 19671 5117
rect 19702 5108 19708 5120
rect 19760 5108 19766 5160
rect 19904 5157 19932 5188
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 20824 5216 20852 5256
rect 20898 5244 20904 5256
rect 20956 5244 20962 5296
rect 21910 5284 21916 5296
rect 21192 5256 21916 5284
rect 20364 5188 20852 5216
rect 19889 5151 19947 5157
rect 19889 5117 19901 5151
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 19978 5108 19984 5160
rect 20036 5108 20042 5160
rect 20364 5148 20392 5188
rect 20548 5157 20576 5188
rect 20272 5120 20392 5148
rect 20441 5151 20499 5157
rect 20272 5080 20300 5120
rect 20441 5117 20453 5151
rect 20487 5117 20499 5151
rect 20441 5111 20499 5117
rect 20533 5151 20591 5157
rect 20533 5117 20545 5151
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 18892 5052 20300 5080
rect 20349 5083 20407 5089
rect 16853 5043 16911 5049
rect 20349 5049 20361 5083
rect 20395 5049 20407 5083
rect 20456 5080 20484 5111
rect 20622 5108 20628 5160
rect 20680 5108 20686 5160
rect 20993 5151 21051 5157
rect 20993 5117 21005 5151
rect 21039 5148 21051 5151
rect 21192 5148 21220 5256
rect 21910 5244 21916 5256
rect 21968 5244 21974 5296
rect 22094 5244 22100 5296
rect 22152 5284 22158 5296
rect 25682 5284 25688 5296
rect 22152 5256 25688 5284
rect 22152 5244 22158 5256
rect 25682 5244 25688 5256
rect 25740 5244 25746 5296
rect 22922 5216 22928 5228
rect 22204 5188 22928 5216
rect 21039 5120 21220 5148
rect 21269 5151 21327 5157
rect 21039 5117 21051 5120
rect 20993 5111 21051 5117
rect 21269 5117 21281 5151
rect 21315 5117 21327 5151
rect 21269 5111 21327 5117
rect 20640 5080 20668 5108
rect 21082 5080 21088 5092
rect 20456 5052 20668 5080
rect 20824 5052 21088 5080
rect 20349 5043 20407 5049
rect 14277 5015 14335 5021
rect 14277 5012 14289 5015
rect 13648 4984 14289 5012
rect 13541 4975 13599 4981
rect 14277 4981 14289 4984
rect 14323 4981 14335 5015
rect 14277 4975 14335 4981
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 14645 5015 14703 5021
rect 14645 5012 14657 5015
rect 14608 4984 14657 5012
rect 14608 4972 14614 4984
rect 14645 4981 14657 4984
rect 14691 4981 14703 5015
rect 14645 4975 14703 4981
rect 15013 5015 15071 5021
rect 15013 4981 15025 5015
rect 15059 5012 15071 5015
rect 15194 5012 15200 5024
rect 15059 4984 15200 5012
rect 15059 4981 15071 4984
rect 15013 4975 15071 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 15933 5015 15991 5021
rect 15933 5012 15945 5015
rect 15436 4984 15945 5012
rect 15436 4972 15442 4984
rect 15933 4981 15945 4984
rect 15979 4981 15991 5015
rect 15933 4975 15991 4981
rect 16022 4972 16028 5024
rect 16080 5012 16086 5024
rect 16390 5012 16396 5024
rect 16080 4984 16396 5012
rect 16080 4972 16086 4984
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 16482 4972 16488 5024
rect 16540 4972 16546 5024
rect 16666 5021 16672 5024
rect 16653 5015 16672 5021
rect 16653 4981 16665 5015
rect 16653 4975 16672 4981
rect 16666 4972 16672 4975
rect 16724 4972 16730 5024
rect 16758 4972 16764 5024
rect 16816 4972 16822 5024
rect 18417 5015 18475 5021
rect 18417 4981 18429 5015
rect 18463 5012 18475 5015
rect 19518 5012 19524 5024
rect 18463 4984 19524 5012
rect 18463 4981 18475 4984
rect 18417 4975 18475 4981
rect 19518 4972 19524 4984
rect 19576 4972 19582 5024
rect 20070 4972 20076 5024
rect 20128 4972 20134 5024
rect 20364 5012 20392 5043
rect 20530 5012 20536 5024
rect 20364 4984 20536 5012
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 20625 5015 20683 5021
rect 20625 4981 20637 5015
rect 20671 5012 20683 5015
rect 20824 5012 20852 5052
rect 21082 5040 21088 5052
rect 21140 5040 21146 5092
rect 21284 5080 21312 5111
rect 21542 5108 21548 5160
rect 21600 5108 21606 5160
rect 21637 5151 21695 5157
rect 21637 5117 21649 5151
rect 21683 5148 21695 5151
rect 21910 5148 21916 5160
rect 21683 5120 21916 5148
rect 21683 5117 21695 5120
rect 21637 5111 21695 5117
rect 21910 5108 21916 5120
rect 21968 5108 21974 5160
rect 22094 5108 22100 5160
rect 22152 5108 22158 5160
rect 22204 5157 22232 5188
rect 22922 5176 22928 5188
rect 22980 5176 22986 5228
rect 23382 5176 23388 5228
rect 23440 5176 23446 5228
rect 22189 5151 22247 5157
rect 22189 5117 22201 5151
rect 22235 5117 22247 5151
rect 22189 5111 22247 5117
rect 22005 5083 22063 5089
rect 21284 5052 21680 5080
rect 20671 4984 20852 5012
rect 20901 5015 20959 5021
rect 20671 4981 20683 4984
rect 20625 4975 20683 4981
rect 20901 4981 20913 5015
rect 20947 5012 20959 5015
rect 21177 5015 21235 5021
rect 21177 5012 21189 5015
rect 20947 4984 21189 5012
rect 20947 4981 20959 4984
rect 20901 4975 20959 4981
rect 21177 4981 21189 4984
rect 21223 4981 21235 5015
rect 21652 5012 21680 5052
rect 22005 5049 22017 5083
rect 22051 5080 22063 5083
rect 23400 5080 23428 5176
rect 22051 5052 23428 5080
rect 22051 5049 22063 5052
rect 22005 5043 22063 5049
rect 22738 5012 22744 5024
rect 21652 4984 22744 5012
rect 21177 4975 21235 4981
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 552 4922 31531 4944
rect 552 4870 8102 4922
rect 8154 4870 8166 4922
rect 8218 4870 8230 4922
rect 8282 4870 8294 4922
rect 8346 4870 8358 4922
rect 8410 4870 15807 4922
rect 15859 4870 15871 4922
rect 15923 4870 15935 4922
rect 15987 4870 15999 4922
rect 16051 4870 16063 4922
rect 16115 4870 23512 4922
rect 23564 4870 23576 4922
rect 23628 4870 23640 4922
rect 23692 4870 23704 4922
rect 23756 4870 23768 4922
rect 23820 4870 31217 4922
rect 31269 4870 31281 4922
rect 31333 4870 31345 4922
rect 31397 4870 31409 4922
rect 31461 4870 31473 4922
rect 31525 4870 31531 4922
rect 552 4848 31531 4870
rect 9306 4768 9312 4820
rect 9364 4768 9370 4820
rect 9861 4811 9919 4817
rect 9861 4777 9873 4811
rect 9907 4808 9919 4811
rect 10134 4808 10140 4820
rect 9907 4780 10140 4808
rect 9907 4777 9919 4780
rect 9861 4771 9919 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10318 4768 10324 4820
rect 10376 4808 10382 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10376 4780 10701 4808
rect 10376 4768 10382 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 10689 4771 10747 4777
rect 10870 4768 10876 4820
rect 10928 4768 10934 4820
rect 11330 4768 11336 4820
rect 11388 4808 11394 4820
rect 11388 4780 11744 4808
rect 11388 4768 11394 4780
rect 9217 4675 9275 4681
rect 9217 4641 9229 4675
rect 9263 4672 9275 4675
rect 9324 4672 9352 4768
rect 9677 4743 9735 4749
rect 9677 4709 9689 4743
rect 9723 4740 9735 4743
rect 9766 4740 9772 4752
rect 9723 4712 9772 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 9766 4700 9772 4712
rect 9824 4740 9830 4752
rect 10229 4743 10287 4749
rect 10229 4740 10241 4743
rect 9824 4712 10241 4740
rect 9824 4700 9830 4712
rect 10229 4709 10241 4712
rect 10275 4740 10287 4743
rect 10888 4740 10916 4768
rect 11514 4740 11520 4752
rect 10275 4712 10916 4740
rect 11348 4712 11520 4740
rect 10275 4709 10287 4712
rect 10229 4703 10287 4709
rect 9263 4644 9352 4672
rect 9263 4641 9275 4644
rect 9217 4635 9275 4641
rect 9490 4632 9496 4684
rect 9548 4632 9554 4684
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 10042 4672 10048 4684
rect 9999 4644 10048 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10134 4632 10140 4684
rect 10192 4632 10198 4684
rect 10321 4675 10379 4681
rect 10321 4641 10333 4675
rect 10367 4672 10379 4675
rect 10502 4672 10508 4684
rect 10367 4644 10508 4672
rect 10367 4641 10379 4644
rect 10321 4635 10379 4641
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 10594 4632 10600 4684
rect 10652 4632 10658 4684
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 11348 4681 11376 4712
rect 11514 4700 11520 4712
rect 11572 4700 11578 4752
rect 10781 4675 10839 4681
rect 10781 4672 10793 4675
rect 10744 4644 10793 4672
rect 10744 4632 10750 4644
rect 10781 4641 10793 4644
rect 10827 4672 10839 4675
rect 11333 4675 11391 4681
rect 11333 4672 11345 4675
rect 10827 4644 11345 4672
rect 10827 4641 10839 4644
rect 10781 4635 10839 4641
rect 11333 4641 11345 4644
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 10612 4604 10640 4632
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 8812 4576 10456 4604
rect 10612 4576 11253 4604
rect 8812 4564 8818 4576
rect 9306 4428 9312 4480
rect 9364 4428 9370 4480
rect 10428 4468 10456 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11348 4604 11376 4635
rect 11422 4632 11428 4684
rect 11480 4632 11486 4684
rect 11716 4681 11744 4780
rect 11790 4768 11796 4820
rect 11848 4768 11854 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 13173 4811 13231 4817
rect 13173 4808 13185 4811
rect 13136 4780 13185 4808
rect 13136 4768 13142 4780
rect 13173 4777 13185 4780
rect 13219 4777 13231 4811
rect 13173 4771 13231 4777
rect 13262 4768 13268 4820
rect 13320 4768 13326 4820
rect 13449 4811 13507 4817
rect 13449 4777 13461 4811
rect 13495 4808 13507 4811
rect 13538 4808 13544 4820
rect 13495 4780 13544 4808
rect 13495 4777 13507 4780
rect 13449 4771 13507 4777
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 14090 4768 14096 4820
rect 14148 4768 14154 4820
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 16117 4811 16175 4817
rect 16117 4808 16129 4811
rect 14700 4780 16129 4808
rect 14700 4768 14706 4780
rect 16117 4777 16129 4780
rect 16163 4777 16175 4811
rect 16117 4771 16175 4777
rect 16206 4768 16212 4820
rect 16264 4768 16270 4820
rect 16482 4768 16488 4820
rect 16540 4768 16546 4820
rect 16577 4811 16635 4817
rect 16577 4777 16589 4811
rect 16623 4808 16635 4811
rect 16758 4808 16764 4820
rect 16623 4780 16764 4808
rect 16623 4777 16635 4780
rect 16577 4771 16635 4777
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 19886 4768 19892 4820
rect 19944 4768 19950 4820
rect 20070 4768 20076 4820
rect 20128 4808 20134 4820
rect 21174 4808 21180 4820
rect 20128 4780 21180 4808
rect 20128 4768 20134 4780
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 21910 4768 21916 4820
rect 21968 4808 21974 4820
rect 23842 4808 23848 4820
rect 21968 4780 23848 4808
rect 21968 4768 21974 4780
rect 23842 4768 23848 4780
rect 23900 4768 23906 4820
rect 12084 4712 13032 4740
rect 12084 4681 12112 4712
rect 13004 4684 13032 4712
rect 11701 4675 11759 4681
rect 11701 4641 11713 4675
rect 11747 4641 11759 4675
rect 11701 4635 11759 4641
rect 12069 4675 12127 4681
rect 12069 4641 12081 4675
rect 12115 4641 12127 4675
rect 12897 4675 12955 4681
rect 12897 4672 12909 4675
rect 12069 4635 12127 4641
rect 12176 4644 12909 4672
rect 12176 4604 12204 4644
rect 12897 4641 12909 4644
rect 12943 4641 12955 4675
rect 12897 4635 12955 4641
rect 11348 4576 12204 4604
rect 12345 4607 12403 4613
rect 11241 4567 11299 4573
rect 12345 4573 12357 4607
rect 12391 4604 12403 4607
rect 12805 4607 12863 4613
rect 12805 4604 12817 4607
rect 12391 4576 12817 4604
rect 12391 4573 12403 4576
rect 12345 4567 12403 4573
rect 12805 4573 12817 4576
rect 12851 4573 12863 4607
rect 12912 4604 12940 4635
rect 12986 4632 12992 4684
rect 13044 4632 13050 4684
rect 13081 4675 13139 4681
rect 13081 4641 13093 4675
rect 13127 4641 13139 4675
rect 13280 4672 13308 4768
rect 14108 4740 14136 4768
rect 14016 4712 14136 4740
rect 14016 4681 14044 4712
rect 14182 4700 14188 4752
rect 14240 4740 14246 4752
rect 14240 4712 16160 4740
rect 14240 4700 14246 4712
rect 13633 4675 13691 4681
rect 13633 4672 13645 4675
rect 13280 4644 13645 4672
rect 13081 4635 13139 4641
rect 13633 4641 13645 4644
rect 13679 4641 13691 4675
rect 13633 4635 13691 4641
rect 14001 4675 14059 4681
rect 14001 4641 14013 4675
rect 14047 4641 14059 4675
rect 14001 4635 14059 4641
rect 13096 4604 13124 4635
rect 14090 4632 14096 4684
rect 14148 4632 14154 4684
rect 14274 4632 14280 4684
rect 14332 4632 14338 4684
rect 14645 4675 14703 4681
rect 14645 4641 14657 4675
rect 14691 4641 14703 4675
rect 14645 4635 14703 4641
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 14826 4672 14832 4684
rect 14783 4644 14832 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 12912 4576 13124 4604
rect 12805 4567 12863 4573
rect 13814 4564 13820 4616
rect 13872 4604 13878 4616
rect 14660 4604 14688 4635
rect 14826 4632 14832 4644
rect 14884 4632 14890 4684
rect 15381 4675 15439 4681
rect 15381 4641 15393 4675
rect 15427 4641 15439 4675
rect 15381 4635 15439 4641
rect 13872 4576 14688 4604
rect 15396 4604 15424 4635
rect 15470 4632 15476 4684
rect 15528 4672 15534 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 15528 4644 15669 4672
rect 15528 4632 15534 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 15838 4632 15844 4684
rect 15896 4632 15902 4684
rect 15930 4632 15936 4684
rect 15988 4632 15994 4684
rect 16132 4681 16160 4712
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4641 16175 4675
rect 16224 4672 16252 4768
rect 16500 4740 16528 4768
rect 16408 4712 16528 4740
rect 16301 4675 16359 4681
rect 16301 4672 16313 4675
rect 16224 4644 16313 4672
rect 16117 4635 16175 4641
rect 16301 4641 16313 4644
rect 16347 4641 16359 4675
rect 16301 4635 16359 4641
rect 16408 4604 16436 4712
rect 16666 4700 16672 4752
rect 16724 4700 16730 4752
rect 16482 4632 16488 4684
rect 16540 4632 16546 4684
rect 15396 4576 16436 4604
rect 13872 4564 13878 4576
rect 10505 4539 10563 4545
rect 10505 4505 10517 4539
rect 10551 4536 10563 4539
rect 10594 4536 10600 4548
rect 10551 4508 10600 4536
rect 10551 4505 10563 4508
rect 10505 4499 10563 4505
rect 10594 4496 10600 4508
rect 10652 4496 10658 4548
rect 11422 4496 11428 4548
rect 11480 4536 11486 4548
rect 12253 4539 12311 4545
rect 12253 4536 12265 4539
rect 11480 4508 12265 4536
rect 11480 4496 11486 4508
rect 12253 4505 12265 4508
rect 12299 4505 12311 4539
rect 12253 4499 12311 4505
rect 12710 4496 12716 4548
rect 12768 4496 12774 4548
rect 15565 4539 15623 4545
rect 15565 4505 15577 4539
rect 15611 4536 15623 4539
rect 15654 4536 15660 4548
rect 15611 4508 15660 4536
rect 15611 4505 15623 4508
rect 15565 4499 15623 4505
rect 15654 4496 15660 4508
rect 15712 4496 15718 4548
rect 15933 4539 15991 4545
rect 15933 4505 15945 4539
rect 15979 4536 15991 4539
rect 16684 4536 16712 4700
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 19904 4681 19932 4768
rect 20732 4712 20944 4740
rect 16945 4675 17003 4681
rect 16945 4672 16957 4675
rect 16908 4644 16957 4672
rect 16908 4632 16914 4644
rect 16945 4641 16957 4644
rect 16991 4641 17003 4675
rect 17201 4675 17259 4681
rect 17201 4672 17213 4675
rect 16945 4635 17003 4641
rect 17052 4644 17213 4672
rect 17052 4604 17080 4644
rect 17201 4641 17213 4644
rect 17247 4641 17259 4675
rect 17201 4635 17259 4641
rect 19889 4675 19947 4681
rect 19889 4641 19901 4675
rect 19935 4641 19947 4675
rect 19889 4635 19947 4641
rect 20438 4632 20444 4684
rect 20496 4632 20502 4684
rect 20732 4681 20760 4712
rect 20717 4675 20775 4681
rect 20717 4641 20729 4675
rect 20763 4641 20775 4675
rect 20717 4635 20775 4641
rect 20809 4675 20867 4681
rect 20809 4641 20821 4675
rect 20855 4641 20867 4675
rect 20809 4635 20867 4641
rect 15979 4508 16712 4536
rect 16776 4576 17080 4604
rect 15979 4505 15991 4508
rect 15933 4499 15991 4505
rect 11517 4471 11575 4477
rect 11517 4468 11529 4471
rect 10428 4440 11529 4468
rect 11517 4437 11529 4440
rect 11563 4437 11575 4471
rect 11517 4431 11575 4437
rect 11790 4428 11796 4480
rect 11848 4468 11854 4480
rect 12161 4471 12219 4477
rect 12161 4468 12173 4471
rect 11848 4440 12173 4468
rect 11848 4428 11854 4440
rect 12161 4437 12173 4440
rect 12207 4468 12219 4471
rect 12728 4468 12756 4496
rect 12207 4440 12756 4468
rect 12207 4437 12219 4440
rect 12161 4431 12219 4437
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 14277 4471 14335 4477
rect 14277 4468 14289 4471
rect 14240 4440 14289 4468
rect 14240 4428 14246 4440
rect 14277 4437 14289 4440
rect 14323 4437 14335 4471
rect 14277 4431 14335 4437
rect 15838 4428 15844 4480
rect 15896 4468 15902 4480
rect 16390 4468 16396 4480
rect 15896 4440 16396 4468
rect 15896 4428 15902 4440
rect 16390 4428 16396 4440
rect 16448 4468 16454 4480
rect 16776 4468 16804 4576
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 20162 4604 20168 4616
rect 19392 4576 20168 4604
rect 19392 4564 19398 4576
rect 20162 4564 20168 4576
rect 20220 4564 20226 4616
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4604 20683 4607
rect 20824 4604 20852 4635
rect 20671 4576 20852 4604
rect 20916 4604 20944 4712
rect 20990 4632 20996 4684
rect 21048 4632 21054 4684
rect 22830 4604 22836 4616
rect 20916 4576 22836 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 20349 4539 20407 4545
rect 20349 4505 20361 4539
rect 20395 4536 20407 4539
rect 20901 4539 20959 4545
rect 20901 4536 20913 4539
rect 20395 4508 20913 4536
rect 20395 4505 20407 4508
rect 20349 4499 20407 4505
rect 20901 4505 20913 4508
rect 20947 4505 20959 4539
rect 20901 4499 20959 4505
rect 21358 4496 21364 4548
rect 21416 4496 21422 4548
rect 16448 4440 16804 4468
rect 16448 4428 16454 4440
rect 18322 4428 18328 4480
rect 18380 4428 18386 4480
rect 19981 4471 20039 4477
rect 19981 4437 19993 4471
rect 20027 4468 20039 4471
rect 21376 4468 21404 4496
rect 20027 4440 21404 4468
rect 20027 4437 20039 4440
rect 19981 4431 20039 4437
rect 552 4378 31372 4400
rect 552 4326 4250 4378
rect 4302 4326 4314 4378
rect 4366 4326 4378 4378
rect 4430 4326 4442 4378
rect 4494 4326 4506 4378
rect 4558 4326 11955 4378
rect 12007 4326 12019 4378
rect 12071 4326 12083 4378
rect 12135 4326 12147 4378
rect 12199 4326 12211 4378
rect 12263 4326 19660 4378
rect 19712 4326 19724 4378
rect 19776 4326 19788 4378
rect 19840 4326 19852 4378
rect 19904 4326 19916 4378
rect 19968 4326 27365 4378
rect 27417 4326 27429 4378
rect 27481 4326 27493 4378
rect 27545 4326 27557 4378
rect 27609 4326 27621 4378
rect 27673 4326 31372 4378
rect 552 4304 31372 4326
rect 9306 4224 9312 4276
rect 9364 4264 9370 4276
rect 9677 4267 9735 4273
rect 9677 4264 9689 4267
rect 9364 4236 9689 4264
rect 9364 4224 9370 4236
rect 9677 4233 9689 4236
rect 9723 4233 9735 4267
rect 11790 4264 11796 4276
rect 9677 4227 9735 4233
rect 10980 4236 11796 4264
rect 9490 4156 9496 4208
rect 9548 4196 9554 4208
rect 9858 4196 9864 4208
rect 9548 4168 9864 4196
rect 9548 4156 9554 4168
rect 9858 4156 9864 4168
rect 9916 4196 9922 4208
rect 10045 4199 10103 4205
rect 10045 4196 10057 4199
rect 9916 4168 10057 4196
rect 9916 4156 9922 4168
rect 10045 4165 10057 4168
rect 10091 4165 10103 4199
rect 10045 4159 10103 4165
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 10980 4128 11008 4236
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 15286 4224 15292 4276
rect 15344 4264 15350 4276
rect 15838 4264 15844 4276
rect 15344 4236 15844 4264
rect 15344 4224 15350 4236
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 18322 4224 18328 4276
rect 18380 4264 18386 4276
rect 21910 4264 21916 4276
rect 18380 4236 21916 4264
rect 18380 4224 18386 4236
rect 21910 4224 21916 4236
rect 21968 4224 21974 4276
rect 11241 4199 11299 4205
rect 11241 4165 11253 4199
rect 11287 4165 11299 4199
rect 11241 4159 11299 4165
rect 8536 4100 9076 4128
rect 8536 4088 8542 4100
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 8754 3884 8760 3936
rect 8812 3884 8818 3936
rect 8956 3924 8984 4023
rect 9048 3992 9076 4100
rect 10152 4100 11008 4128
rect 11256 4128 11284 4159
rect 19518 4156 19524 4208
rect 19576 4196 19582 4208
rect 20622 4196 20628 4208
rect 19576 4168 20628 4196
rect 19576 4156 19582 4168
rect 20622 4156 20628 4168
rect 20680 4156 20686 4208
rect 11256 4100 11744 4128
rect 10152 4072 10180 4100
rect 10134 4020 10140 4072
rect 10192 4020 10198 4072
rect 10321 4063 10379 4069
rect 10321 4029 10333 4063
rect 10367 4060 10379 4063
rect 10502 4060 10508 4072
rect 10367 4032 10508 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 10612 4069 10640 4100
rect 10980 4069 11008 4100
rect 10597 4063 10655 4069
rect 10597 4029 10609 4063
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 11422 4060 11428 4072
rect 11287 4032 11428 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 11609 4063 11667 4069
rect 11609 4029 11621 4063
rect 11655 4029 11667 4063
rect 11716 4060 11744 4100
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 15657 4131 15715 4137
rect 15657 4128 15669 4131
rect 14976 4100 15669 4128
rect 14976 4088 14982 4100
rect 15657 4097 15669 4100
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 14182 4069 14188 4072
rect 11865 4063 11923 4069
rect 11865 4060 11877 4063
rect 11716 4032 11877 4060
rect 11609 4023 11667 4029
rect 11865 4029 11877 4032
rect 11911 4029 11923 4063
rect 11865 4023 11923 4029
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4029 13967 4063
rect 14176 4060 14188 4069
rect 14143 4032 14188 4060
rect 13909 4023 13967 4029
rect 14176 4023 14188 4032
rect 11624 3992 11652 4023
rect 13924 3992 13952 4023
rect 14182 4020 14188 4023
rect 14240 4020 14246 4072
rect 14936 3992 14964 4088
rect 9048 3964 14964 3992
rect 15924 3995 15982 4001
rect 15924 3961 15936 3995
rect 15970 3992 15982 3995
rect 16390 3992 16396 4004
rect 15970 3964 16396 3992
rect 15970 3961 15982 3964
rect 15924 3955 15982 3961
rect 16390 3952 16396 3964
rect 16448 3952 16454 4004
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 8956 3896 9505 3924
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 10137 3927 10195 3933
rect 10137 3924 10149 3927
rect 9723 3896 10149 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 10137 3893 10149 3896
rect 10183 3893 10195 3927
rect 10137 3887 10195 3893
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10284 3896 10517 3924
rect 10284 3884 10290 3896
rect 10505 3893 10517 3896
rect 10551 3924 10563 3927
rect 10594 3924 10600 3936
rect 10551 3896 10600 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10594 3884 10600 3896
rect 10652 3924 10658 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10652 3896 11069 3924
rect 10652 3884 10658 3896
rect 11057 3893 11069 3896
rect 11103 3924 11115 3927
rect 12986 3924 12992 3936
rect 11103 3896 12992 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 17034 3884 17040 3936
rect 17092 3884 17098 3936
rect 552 3834 31531 3856
rect 552 3782 8102 3834
rect 8154 3782 8166 3834
rect 8218 3782 8230 3834
rect 8282 3782 8294 3834
rect 8346 3782 8358 3834
rect 8410 3782 15807 3834
rect 15859 3782 15871 3834
rect 15923 3782 15935 3834
rect 15987 3782 15999 3834
rect 16051 3782 16063 3834
rect 16115 3782 23512 3834
rect 23564 3782 23576 3834
rect 23628 3782 23640 3834
rect 23692 3782 23704 3834
rect 23756 3782 23768 3834
rect 23820 3782 31217 3834
rect 31269 3782 31281 3834
rect 31333 3782 31345 3834
rect 31397 3782 31409 3834
rect 31461 3782 31473 3834
rect 31525 3782 31531 3834
rect 552 3760 31531 3782
rect 9858 3680 9864 3732
rect 9916 3680 9922 3732
rect 10029 3723 10087 3729
rect 10029 3689 10041 3723
rect 10075 3720 10087 3723
rect 10134 3720 10140 3732
rect 10075 3692 10140 3720
rect 10075 3689 10087 3692
rect 10029 3683 10087 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 12621 3723 12679 3729
rect 12621 3720 12633 3723
rect 10336 3692 12633 3720
rect 8656 3655 8714 3661
rect 8656 3621 8668 3655
rect 8702 3652 8714 3655
rect 8754 3652 8760 3664
rect 8702 3624 8760 3652
rect 8702 3621 8714 3624
rect 8656 3615 8714 3621
rect 8754 3612 8760 3624
rect 8812 3612 8818 3664
rect 10226 3612 10232 3664
rect 10284 3612 10290 3664
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 8478 3584 8484 3596
rect 8435 3556 8484 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 9030 3544 9036 3596
rect 9088 3584 9094 3596
rect 10336 3584 10364 3692
rect 12621 3689 12633 3692
rect 12667 3689 12679 3723
rect 12621 3683 12679 3689
rect 14274 3680 14280 3732
rect 14332 3720 14338 3732
rect 14461 3723 14519 3729
rect 14461 3720 14473 3723
rect 14332 3692 14473 3720
rect 14332 3680 14338 3692
rect 14461 3689 14473 3692
rect 14507 3689 14519 3723
rect 14461 3683 14519 3689
rect 16117 3723 16175 3729
rect 16117 3689 16129 3723
rect 16163 3720 16175 3723
rect 16390 3720 16396 3732
rect 16163 3692 16396 3720
rect 16163 3689 16175 3692
rect 16117 3683 16175 3689
rect 16390 3680 16396 3692
rect 16448 3680 16454 3732
rect 12170 3655 12228 3661
rect 12170 3652 12182 3655
rect 9088 3556 10364 3584
rect 11026 3624 12182 3652
rect 9088 3544 9094 3556
rect 10502 3448 10508 3460
rect 10060 3420 10508 3448
rect 10060 3389 10088 3420
rect 10502 3408 10508 3420
rect 10560 3448 10566 3460
rect 11026 3448 11054 3624
rect 12170 3621 12182 3624
rect 12216 3621 12228 3655
rect 12170 3615 12228 3621
rect 12820 3624 14044 3652
rect 12820 3596 12848 3624
rect 12437 3587 12495 3593
rect 12437 3553 12449 3587
rect 12483 3584 12495 3587
rect 12802 3584 12808 3596
rect 12483 3556 12808 3584
rect 12483 3553 12495 3556
rect 12437 3547 12495 3553
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 12986 3544 12992 3596
rect 13044 3584 13050 3596
rect 14016 3593 14044 3624
rect 14090 3612 14096 3664
rect 14148 3652 14154 3664
rect 15378 3652 15384 3664
rect 14148 3624 15384 3652
rect 14148 3612 14154 3624
rect 14200 3593 14228 3624
rect 15378 3612 15384 3624
rect 15436 3652 15442 3664
rect 16206 3652 16212 3664
rect 15436 3624 16212 3652
rect 15436 3612 15442 3624
rect 16206 3612 16212 3624
rect 16264 3652 16270 3664
rect 17034 3652 17040 3664
rect 16264 3624 17040 3652
rect 16264 3612 16270 3624
rect 17034 3612 17040 3624
rect 17092 3652 17098 3664
rect 17190 3655 17248 3661
rect 17190 3652 17202 3655
rect 17092 3624 17202 3652
rect 17092 3612 17098 3624
rect 17190 3621 17202 3624
rect 17236 3621 17248 3655
rect 17190 3615 17248 3621
rect 13734 3587 13792 3593
rect 13734 3584 13746 3587
rect 13044 3556 13746 3584
rect 13044 3544 13050 3556
rect 13734 3553 13746 3556
rect 13780 3553 13792 3587
rect 13734 3547 13792 3553
rect 14001 3587 14059 3593
rect 14001 3553 14013 3587
rect 14047 3553 14059 3587
rect 14001 3547 14059 3553
rect 14185 3587 14243 3593
rect 14185 3553 14197 3587
rect 14231 3553 14243 3587
rect 14185 3547 14243 3553
rect 15010 3544 15016 3596
rect 15068 3593 15074 3596
rect 15068 3584 15079 3593
rect 15068 3556 15194 3584
rect 15068 3547 15079 3556
rect 15068 3544 15074 3547
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 14507 3488 14933 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 15166 3516 15194 3556
rect 16114 3544 16120 3596
rect 16172 3584 16178 3596
rect 16301 3587 16359 3593
rect 16301 3584 16313 3587
rect 16172 3556 16313 3584
rect 16172 3544 16178 3556
rect 16301 3553 16313 3556
rect 16347 3553 16359 3587
rect 16301 3547 16359 3553
rect 16393 3587 16451 3593
rect 16393 3553 16405 3587
rect 16439 3584 16451 3587
rect 16482 3584 16488 3596
rect 16439 3556 16488 3584
rect 16439 3553 16451 3556
rect 16393 3547 16451 3553
rect 16408 3516 16436 3547
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 16850 3544 16856 3596
rect 16908 3584 16914 3596
rect 16945 3587 17003 3593
rect 16945 3584 16957 3587
rect 16908 3556 16957 3584
rect 16908 3544 16914 3556
rect 16945 3553 16957 3556
rect 16991 3553 17003 3587
rect 16945 3547 17003 3553
rect 15166 3488 16436 3516
rect 14921 3479 14979 3485
rect 10560 3420 11054 3448
rect 14277 3451 14335 3457
rect 10560 3408 10566 3420
rect 14277 3417 14289 3451
rect 14323 3448 14335 3451
rect 15286 3448 15292 3460
rect 14323 3420 15292 3448
rect 14323 3417 14335 3420
rect 14277 3411 14335 3417
rect 15286 3408 15292 3420
rect 15344 3408 15350 3460
rect 15749 3451 15807 3457
rect 15749 3417 15761 3451
rect 15795 3448 15807 3451
rect 16485 3451 16543 3457
rect 16485 3448 16497 3451
rect 15795 3420 16497 3448
rect 15795 3417 15807 3420
rect 15749 3411 15807 3417
rect 16485 3417 16497 3420
rect 16531 3417 16543 3451
rect 16485 3411 16543 3417
rect 9769 3383 9827 3389
rect 9769 3349 9781 3383
rect 9815 3380 9827 3383
rect 10045 3383 10103 3389
rect 10045 3380 10057 3383
rect 9815 3352 10057 3380
rect 9815 3349 9827 3352
rect 9769 3343 9827 3349
rect 10045 3349 10057 3352
rect 10091 3349 10103 3383
rect 10045 3343 10103 3349
rect 10318 3340 10324 3392
rect 10376 3380 10382 3392
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 10376 3352 11069 3380
rect 10376 3340 10382 3352
rect 11057 3349 11069 3352
rect 11103 3349 11115 3383
rect 11057 3343 11115 3349
rect 15841 3383 15899 3389
rect 15841 3349 15853 3383
rect 15887 3380 15899 3383
rect 16114 3380 16120 3392
rect 15887 3352 16120 3380
rect 15887 3349 15899 3352
rect 15841 3343 15899 3349
rect 16114 3340 16120 3352
rect 16172 3340 16178 3392
rect 18325 3383 18383 3389
rect 18325 3349 18337 3383
rect 18371 3380 18383 3383
rect 23198 3380 23204 3392
rect 18371 3352 23204 3380
rect 18371 3349 18383 3352
rect 18325 3343 18383 3349
rect 23198 3340 23204 3352
rect 23256 3340 23262 3392
rect 552 3290 31372 3312
rect 552 3238 4250 3290
rect 4302 3238 4314 3290
rect 4366 3238 4378 3290
rect 4430 3238 4442 3290
rect 4494 3238 4506 3290
rect 4558 3238 11955 3290
rect 12007 3238 12019 3290
rect 12071 3238 12083 3290
rect 12135 3238 12147 3290
rect 12199 3238 12211 3290
rect 12263 3238 19660 3290
rect 19712 3238 19724 3290
rect 19776 3238 19788 3290
rect 19840 3238 19852 3290
rect 19904 3238 19916 3290
rect 19968 3238 27365 3290
rect 27417 3238 27429 3290
rect 27481 3238 27493 3290
rect 27545 3238 27557 3290
rect 27609 3238 27621 3290
rect 27673 3238 31372 3290
rect 552 3216 31372 3238
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 11698 2836 11704 2848
rect 9732 2808 11704 2836
rect 9732 2796 9738 2808
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 552 2746 31531 2768
rect 552 2694 8102 2746
rect 8154 2694 8166 2746
rect 8218 2694 8230 2746
rect 8282 2694 8294 2746
rect 8346 2694 8358 2746
rect 8410 2694 15807 2746
rect 15859 2694 15871 2746
rect 15923 2694 15935 2746
rect 15987 2694 15999 2746
rect 16051 2694 16063 2746
rect 16115 2694 23512 2746
rect 23564 2694 23576 2746
rect 23628 2694 23640 2746
rect 23692 2694 23704 2746
rect 23756 2694 23768 2746
rect 23820 2694 31217 2746
rect 31269 2694 31281 2746
rect 31333 2694 31345 2746
rect 31397 2694 31409 2746
rect 31461 2694 31473 2746
rect 31525 2694 31531 2746
rect 552 2672 31531 2694
rect 552 2202 31372 2224
rect 552 2150 4250 2202
rect 4302 2150 4314 2202
rect 4366 2150 4378 2202
rect 4430 2150 4442 2202
rect 4494 2150 4506 2202
rect 4558 2150 11955 2202
rect 12007 2150 12019 2202
rect 12071 2150 12083 2202
rect 12135 2150 12147 2202
rect 12199 2150 12211 2202
rect 12263 2150 19660 2202
rect 19712 2150 19724 2202
rect 19776 2150 19788 2202
rect 19840 2150 19852 2202
rect 19904 2150 19916 2202
rect 19968 2150 27365 2202
rect 27417 2150 27429 2202
rect 27481 2150 27493 2202
rect 27545 2150 27557 2202
rect 27609 2150 27621 2202
rect 27673 2150 31372 2202
rect 552 2128 31372 2150
rect 552 1658 31531 1680
rect 552 1606 8102 1658
rect 8154 1606 8166 1658
rect 8218 1606 8230 1658
rect 8282 1606 8294 1658
rect 8346 1606 8358 1658
rect 8410 1606 15807 1658
rect 15859 1606 15871 1658
rect 15923 1606 15935 1658
rect 15987 1606 15999 1658
rect 16051 1606 16063 1658
rect 16115 1606 23512 1658
rect 23564 1606 23576 1658
rect 23628 1606 23640 1658
rect 23692 1606 23704 1658
rect 23756 1606 23768 1658
rect 23820 1606 31217 1658
rect 31269 1606 31281 1658
rect 31333 1606 31345 1658
rect 31397 1606 31409 1658
rect 31461 1606 31473 1658
rect 31525 1606 31531 1658
rect 552 1584 31531 1606
rect 552 1114 31372 1136
rect 552 1062 4250 1114
rect 4302 1062 4314 1114
rect 4366 1062 4378 1114
rect 4430 1062 4442 1114
rect 4494 1062 4506 1114
rect 4558 1062 11955 1114
rect 12007 1062 12019 1114
rect 12071 1062 12083 1114
rect 12135 1062 12147 1114
rect 12199 1062 12211 1114
rect 12263 1062 19660 1114
rect 19712 1062 19724 1114
rect 19776 1062 19788 1114
rect 19840 1062 19852 1114
rect 19904 1062 19916 1114
rect 19968 1062 27365 1114
rect 27417 1062 27429 1114
rect 27481 1062 27493 1114
rect 27545 1062 27557 1114
rect 27609 1062 27621 1114
rect 27673 1062 31372 1114
rect 552 1040 31372 1062
rect 8021 1003 8079 1009
rect 8021 969 8033 1003
rect 8067 1000 8079 1003
rect 8662 1000 8668 1012
rect 8067 972 8668 1000
rect 8067 969 8079 972
rect 8021 963 8079 969
rect 8662 960 8668 972
rect 8720 960 8726 1012
rect 7834 756 7840 808
rect 7892 756 7898 808
rect 552 570 31531 592
rect 552 518 8102 570
rect 8154 518 8166 570
rect 8218 518 8230 570
rect 8282 518 8294 570
rect 8346 518 8358 570
rect 8410 518 15807 570
rect 15859 518 15871 570
rect 15923 518 15935 570
rect 15987 518 15999 570
rect 16051 518 16063 570
rect 16115 518 23512 570
rect 23564 518 23576 570
rect 23628 518 23640 570
rect 23692 518 23704 570
rect 23756 518 23768 570
rect 23820 518 31217 570
rect 31269 518 31281 570
rect 31333 518 31345 570
rect 31397 518 31409 570
rect 31461 518 31473 570
rect 31525 518 31531 570
rect 552 496 31531 518
rect 16022 416 16028 468
rect 16080 456 16086 468
rect 16298 456 16304 468
rect 16080 428 16304 456
rect 16080 416 16086 428
rect 16298 416 16304 428
rect 16356 416 16362 468
<< via1 >>
rect 8102 19014 8154 19066
rect 8166 19014 8218 19066
rect 8230 19014 8282 19066
rect 8294 19014 8346 19066
rect 8358 19014 8410 19066
rect 15807 19014 15859 19066
rect 15871 19014 15923 19066
rect 15935 19014 15987 19066
rect 15999 19014 16051 19066
rect 16063 19014 16115 19066
rect 23512 19014 23564 19066
rect 23576 19014 23628 19066
rect 23640 19014 23692 19066
rect 23704 19014 23756 19066
rect 23768 19014 23820 19066
rect 31217 19014 31269 19066
rect 31281 19014 31333 19066
rect 31345 19014 31397 19066
rect 31409 19014 31461 19066
rect 31473 19014 31525 19066
rect 4250 18470 4302 18522
rect 4314 18470 4366 18522
rect 4378 18470 4430 18522
rect 4442 18470 4494 18522
rect 4506 18470 4558 18522
rect 11955 18470 12007 18522
rect 12019 18470 12071 18522
rect 12083 18470 12135 18522
rect 12147 18470 12199 18522
rect 12211 18470 12263 18522
rect 19660 18470 19712 18522
rect 19724 18470 19776 18522
rect 19788 18470 19840 18522
rect 19852 18470 19904 18522
rect 19916 18470 19968 18522
rect 27365 18470 27417 18522
rect 27429 18470 27481 18522
rect 27493 18470 27545 18522
rect 27557 18470 27609 18522
rect 27621 18470 27673 18522
rect 8102 17926 8154 17978
rect 8166 17926 8218 17978
rect 8230 17926 8282 17978
rect 8294 17926 8346 17978
rect 8358 17926 8410 17978
rect 15807 17926 15859 17978
rect 15871 17926 15923 17978
rect 15935 17926 15987 17978
rect 15999 17926 16051 17978
rect 16063 17926 16115 17978
rect 23512 17926 23564 17978
rect 23576 17926 23628 17978
rect 23640 17926 23692 17978
rect 23704 17926 23756 17978
rect 23768 17926 23820 17978
rect 31217 17926 31269 17978
rect 31281 17926 31333 17978
rect 31345 17926 31397 17978
rect 31409 17926 31461 17978
rect 31473 17926 31525 17978
rect 20996 17552 21048 17604
rect 21180 17484 21232 17536
rect 4250 17382 4302 17434
rect 4314 17382 4366 17434
rect 4378 17382 4430 17434
rect 4442 17382 4494 17434
rect 4506 17382 4558 17434
rect 11955 17382 12007 17434
rect 12019 17382 12071 17434
rect 12083 17382 12135 17434
rect 12147 17382 12199 17434
rect 12211 17382 12263 17434
rect 19660 17382 19712 17434
rect 19724 17382 19776 17434
rect 19788 17382 19840 17434
rect 19852 17382 19904 17434
rect 19916 17382 19968 17434
rect 27365 17382 27417 17434
rect 27429 17382 27481 17434
rect 27493 17382 27545 17434
rect 27557 17382 27609 17434
rect 27621 17382 27673 17434
rect 11336 17280 11388 17332
rect 21272 17280 21324 17332
rect 21824 17280 21876 17332
rect 23296 17280 23348 17332
rect 9772 17076 9824 17128
rect 12348 17212 12400 17264
rect 11520 17076 11572 17128
rect 8668 17008 8720 17060
rect 11152 17008 11204 17060
rect 11244 17008 11296 17060
rect 11888 17076 11940 17128
rect 12072 17119 12124 17128
rect 12072 17085 12081 17119
rect 12081 17085 12115 17119
rect 12115 17085 12124 17119
rect 12072 17076 12124 17085
rect 12624 17119 12676 17128
rect 12624 17085 12633 17119
rect 12633 17085 12667 17119
rect 12667 17085 12676 17119
rect 12624 17076 12676 17085
rect 12992 17119 13044 17128
rect 12992 17085 13001 17119
rect 13001 17085 13035 17119
rect 13035 17085 13044 17119
rect 12992 17076 13044 17085
rect 13820 17119 13872 17128
rect 13820 17085 13829 17119
rect 13829 17085 13863 17119
rect 13863 17085 13872 17119
rect 13820 17076 13872 17085
rect 14004 17076 14056 17128
rect 19524 17144 19576 17196
rect 20352 17119 20404 17128
rect 20352 17085 20361 17119
rect 20361 17085 20395 17119
rect 20395 17085 20404 17119
rect 20352 17076 20404 17085
rect 22100 17212 22152 17264
rect 22284 17212 22336 17264
rect 23940 17212 23992 17264
rect 20996 17119 21048 17128
rect 20444 17008 20496 17060
rect 20996 17085 21005 17119
rect 21005 17085 21039 17119
rect 21039 17085 21048 17119
rect 20996 17076 21048 17085
rect 21456 17119 21508 17128
rect 21456 17085 21465 17119
rect 21465 17085 21499 17119
rect 21499 17085 21508 17119
rect 21456 17076 21508 17085
rect 21640 17076 21692 17128
rect 22744 17144 22796 17196
rect 22008 17119 22060 17128
rect 22008 17085 22017 17119
rect 22017 17085 22051 17119
rect 22051 17085 22060 17119
rect 22008 17076 22060 17085
rect 21088 17008 21140 17060
rect 22376 17119 22428 17128
rect 22376 17085 22385 17119
rect 22385 17085 22419 17119
rect 22419 17085 22428 17119
rect 22376 17076 22428 17085
rect 24952 17076 25004 17128
rect 11520 16940 11572 16992
rect 12532 16983 12584 16992
rect 12532 16949 12541 16983
rect 12541 16949 12575 16983
rect 12575 16949 12584 16983
rect 12532 16940 12584 16949
rect 13728 16940 13780 16992
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 13912 16940 13964 16949
rect 14924 16983 14976 16992
rect 14924 16949 14933 16983
rect 14933 16949 14967 16983
rect 14967 16949 14976 16983
rect 14924 16940 14976 16949
rect 19248 16940 19300 16992
rect 20812 16983 20864 16992
rect 20812 16949 20821 16983
rect 20821 16949 20855 16983
rect 20855 16949 20864 16983
rect 20812 16940 20864 16949
rect 21640 16983 21692 16992
rect 21640 16949 21649 16983
rect 21649 16949 21683 16983
rect 21683 16949 21692 16983
rect 21640 16940 21692 16949
rect 21916 16940 21968 16992
rect 22652 16940 22704 16992
rect 25136 17008 25188 17060
rect 23020 16983 23072 16992
rect 23020 16949 23029 16983
rect 23029 16949 23063 16983
rect 23063 16949 23072 16983
rect 23020 16940 23072 16949
rect 8102 16838 8154 16890
rect 8166 16838 8218 16890
rect 8230 16838 8282 16890
rect 8294 16838 8346 16890
rect 8358 16838 8410 16890
rect 15807 16838 15859 16890
rect 15871 16838 15923 16890
rect 15935 16838 15987 16890
rect 15999 16838 16051 16890
rect 16063 16838 16115 16890
rect 23512 16838 23564 16890
rect 23576 16838 23628 16890
rect 23640 16838 23692 16890
rect 23704 16838 23756 16890
rect 23768 16838 23820 16890
rect 31217 16838 31269 16890
rect 31281 16838 31333 16890
rect 31345 16838 31397 16890
rect 31409 16838 31461 16890
rect 31473 16838 31525 16890
rect 7932 16736 7984 16788
rect 8760 16668 8812 16720
rect 10876 16668 10928 16720
rect 12624 16736 12676 16788
rect 13820 16779 13872 16788
rect 13820 16745 13829 16779
rect 13829 16745 13863 16779
rect 13863 16745 13872 16779
rect 13820 16736 13872 16745
rect 14004 16736 14056 16788
rect 14924 16736 14976 16788
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 10692 16600 10744 16652
rect 10968 16643 11020 16652
rect 10968 16609 10977 16643
rect 10977 16609 11011 16643
rect 11011 16609 11020 16643
rect 10968 16600 11020 16609
rect 11060 16643 11112 16652
rect 11060 16609 11069 16643
rect 11069 16609 11103 16643
rect 11103 16609 11112 16643
rect 11060 16600 11112 16609
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11244 16600 11296 16609
rect 11336 16643 11388 16652
rect 11336 16609 11345 16643
rect 11345 16609 11379 16643
rect 11379 16609 11388 16643
rect 11336 16600 11388 16609
rect 12072 16600 12124 16652
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 12440 16600 12492 16652
rect 10508 16464 10560 16516
rect 10600 16464 10652 16516
rect 11704 16532 11756 16584
rect 13728 16643 13780 16652
rect 13728 16609 13737 16643
rect 13737 16609 13771 16643
rect 13771 16609 13780 16643
rect 13728 16600 13780 16609
rect 14648 16600 14700 16652
rect 14924 16643 14976 16652
rect 14924 16609 14933 16643
rect 14933 16609 14967 16643
rect 14967 16609 14976 16643
rect 14924 16600 14976 16609
rect 15568 16668 15620 16720
rect 20260 16668 20312 16720
rect 15752 16600 15804 16652
rect 10968 16464 11020 16516
rect 16120 16532 16172 16584
rect 16856 16532 16908 16584
rect 19248 16643 19300 16652
rect 19248 16609 19257 16643
rect 19257 16609 19291 16643
rect 19291 16609 19300 16643
rect 19248 16600 19300 16609
rect 19340 16643 19392 16652
rect 19340 16609 19349 16643
rect 19349 16609 19383 16643
rect 19383 16609 19392 16643
rect 19340 16600 19392 16609
rect 19524 16600 19576 16652
rect 21364 16736 21416 16788
rect 21456 16736 21508 16788
rect 22652 16736 22704 16788
rect 22744 16779 22796 16788
rect 22744 16745 22753 16779
rect 22753 16745 22787 16779
rect 22787 16745 22796 16779
rect 22744 16736 22796 16745
rect 22836 16736 22888 16788
rect 23112 16736 23164 16788
rect 20904 16668 20956 16720
rect 21088 16668 21140 16720
rect 21272 16668 21324 16720
rect 13728 16464 13780 16516
rect 14464 16464 14516 16516
rect 15016 16464 15068 16516
rect 11428 16396 11480 16448
rect 12440 16439 12492 16448
rect 12440 16405 12449 16439
rect 12449 16405 12483 16439
rect 12483 16405 12492 16439
rect 12440 16396 12492 16405
rect 12808 16439 12860 16448
rect 12808 16405 12817 16439
rect 12817 16405 12851 16439
rect 12851 16405 12860 16439
rect 12808 16396 12860 16405
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 13176 16396 13228 16448
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 13452 16396 13504 16448
rect 14924 16396 14976 16448
rect 15200 16396 15252 16448
rect 19432 16439 19484 16448
rect 19432 16405 19441 16439
rect 19441 16405 19475 16439
rect 19475 16405 19484 16439
rect 19432 16396 19484 16405
rect 19524 16396 19576 16448
rect 19984 16439 20036 16448
rect 19984 16405 19993 16439
rect 19993 16405 20027 16439
rect 20027 16405 20036 16439
rect 19984 16396 20036 16405
rect 20076 16396 20128 16448
rect 20352 16575 20404 16584
rect 20352 16541 20361 16575
rect 20361 16541 20395 16575
rect 20395 16541 20404 16575
rect 20352 16532 20404 16541
rect 21456 16643 21508 16652
rect 21456 16609 21465 16643
rect 21465 16609 21499 16643
rect 21499 16609 21508 16643
rect 21456 16600 21508 16609
rect 21272 16532 21324 16584
rect 21732 16600 21784 16652
rect 22008 16643 22060 16652
rect 22008 16609 22017 16643
rect 22017 16609 22051 16643
rect 22051 16609 22060 16643
rect 22008 16600 22060 16609
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 23296 16711 23348 16720
rect 23296 16677 23305 16711
rect 23305 16677 23339 16711
rect 23339 16677 23348 16711
rect 23296 16668 23348 16677
rect 22744 16532 22796 16584
rect 23664 16643 23716 16652
rect 23664 16609 23673 16643
rect 23673 16609 23707 16643
rect 23707 16609 23716 16643
rect 23664 16600 23716 16609
rect 23756 16532 23808 16584
rect 20536 16396 20588 16448
rect 24308 16464 24360 16516
rect 21180 16396 21232 16448
rect 22468 16396 22520 16448
rect 23572 16396 23624 16448
rect 24584 16396 24636 16448
rect 4250 16294 4302 16346
rect 4314 16294 4366 16346
rect 4378 16294 4430 16346
rect 4442 16294 4494 16346
rect 4506 16294 4558 16346
rect 11955 16294 12007 16346
rect 12019 16294 12071 16346
rect 12083 16294 12135 16346
rect 12147 16294 12199 16346
rect 12211 16294 12263 16346
rect 19660 16294 19712 16346
rect 19724 16294 19776 16346
rect 19788 16294 19840 16346
rect 19852 16294 19904 16346
rect 19916 16294 19968 16346
rect 27365 16294 27417 16346
rect 27429 16294 27481 16346
rect 27493 16294 27545 16346
rect 27557 16294 27609 16346
rect 27621 16294 27673 16346
rect 7472 16192 7524 16244
rect 9772 16124 9824 16176
rect 9864 16124 9916 16176
rect 10968 16235 11020 16244
rect 10968 16201 10977 16235
rect 10977 16201 11011 16235
rect 11011 16201 11020 16235
rect 10968 16192 11020 16201
rect 11060 16192 11112 16244
rect 12348 16192 12400 16244
rect 12624 16192 12676 16244
rect 13912 16192 13964 16244
rect 14004 16235 14056 16244
rect 14004 16201 14013 16235
rect 14013 16201 14047 16235
rect 14047 16201 14056 16235
rect 14004 16192 14056 16201
rect 14556 16192 14608 16244
rect 15752 16192 15804 16244
rect 9772 16031 9824 16040
rect 9772 15997 9781 16031
rect 9781 15997 9815 16031
rect 9815 15997 9824 16031
rect 9772 15988 9824 15997
rect 10140 15988 10192 16040
rect 10508 15988 10560 16040
rect 10692 15988 10744 16040
rect 10968 15988 11020 16040
rect 11520 16056 11572 16108
rect 11888 16124 11940 16176
rect 14832 16124 14884 16176
rect 16304 16124 16356 16176
rect 11244 15988 11296 16040
rect 12440 16056 12492 16108
rect 12624 16031 12676 16040
rect 12624 15997 12633 16031
rect 12633 15997 12667 16031
rect 12667 15997 12676 16031
rect 12624 15988 12676 15997
rect 12808 16031 12860 16040
rect 12808 15997 12817 16031
rect 12817 15997 12851 16031
rect 12851 15997 12860 16031
rect 12808 15988 12860 15997
rect 13084 16031 13136 16040
rect 13084 15997 13093 16031
rect 13093 15997 13127 16031
rect 13127 15997 13136 16031
rect 13084 15988 13136 15997
rect 13360 16031 13412 16040
rect 13360 15997 13369 16031
rect 13369 15997 13403 16031
rect 13403 15997 13412 16031
rect 13360 15988 13412 15997
rect 8024 15852 8076 15904
rect 10140 15895 10192 15904
rect 10140 15861 10149 15895
rect 10149 15861 10183 15895
rect 10183 15861 10192 15895
rect 10140 15852 10192 15861
rect 10324 15852 10376 15904
rect 10508 15852 10560 15904
rect 10968 15852 11020 15904
rect 11152 15852 11204 15904
rect 11520 15895 11572 15904
rect 11520 15861 11529 15895
rect 11529 15861 11563 15895
rect 11563 15861 11572 15895
rect 11520 15852 11572 15861
rect 12348 15895 12400 15904
rect 12348 15861 12357 15895
rect 12357 15861 12391 15895
rect 12391 15861 12400 15895
rect 12348 15852 12400 15861
rect 12716 15895 12768 15904
rect 12716 15861 12725 15895
rect 12725 15861 12759 15895
rect 12759 15861 12768 15895
rect 12716 15852 12768 15861
rect 12808 15852 12860 15904
rect 13820 15920 13872 15972
rect 14464 16031 14516 16040
rect 14464 15997 14473 16031
rect 14473 15997 14507 16031
rect 14507 15997 14516 16031
rect 14464 15988 14516 15997
rect 15292 15988 15344 16040
rect 15660 15988 15712 16040
rect 16120 15988 16172 16040
rect 18236 16192 18288 16244
rect 19524 16192 19576 16244
rect 20260 16192 20312 16244
rect 20812 16192 20864 16244
rect 20904 16192 20956 16244
rect 21364 16192 21416 16244
rect 22100 16235 22152 16244
rect 22100 16201 22109 16235
rect 22109 16201 22143 16235
rect 22143 16201 22152 16235
rect 22100 16192 22152 16201
rect 22468 16192 22520 16244
rect 19800 16124 19852 16176
rect 18788 16056 18840 16108
rect 19616 16056 19668 16108
rect 23296 16192 23348 16244
rect 23664 16192 23716 16244
rect 23388 16124 23440 16176
rect 17960 15988 18012 16040
rect 18328 16031 18380 16040
rect 18328 15997 18337 16031
rect 18337 15997 18371 16031
rect 18371 15997 18380 16031
rect 18328 15988 18380 15997
rect 19432 16031 19484 16040
rect 19432 15997 19441 16031
rect 19441 15997 19475 16031
rect 19475 15997 19484 16031
rect 19432 15988 19484 15997
rect 14740 15852 14792 15904
rect 14832 15895 14884 15904
rect 14832 15861 14841 15895
rect 14841 15861 14875 15895
rect 14875 15861 14884 15895
rect 14832 15852 14884 15861
rect 15476 15895 15528 15904
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 18420 15895 18472 15904
rect 18420 15861 18429 15895
rect 18429 15861 18463 15895
rect 18463 15861 18472 15895
rect 18420 15852 18472 15861
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 19156 15852 19208 15904
rect 19432 15852 19484 15904
rect 19984 16031 20036 16040
rect 19984 15997 19993 16031
rect 19993 15997 20027 16031
rect 20027 15997 20036 16031
rect 19984 15988 20036 15997
rect 20352 15988 20404 16040
rect 20904 16031 20956 16040
rect 20904 15997 20913 16031
rect 20913 15997 20947 16031
rect 20947 15997 20956 16031
rect 20904 15988 20956 15997
rect 21180 15988 21232 16040
rect 21364 16031 21416 16040
rect 21364 15997 21373 16031
rect 21373 15997 21407 16031
rect 21407 15997 21416 16031
rect 21364 15988 21416 15997
rect 22376 16056 22428 16108
rect 22744 16056 22796 16108
rect 22192 16031 22244 16040
rect 22192 15997 22201 16031
rect 22201 15997 22235 16031
rect 22235 15997 22244 16031
rect 22192 15988 22244 15997
rect 22468 15988 22520 16040
rect 22836 15988 22888 16040
rect 23296 16031 23348 16040
rect 23296 15997 23305 16031
rect 23305 15997 23339 16031
rect 23339 15997 23348 16031
rect 23296 15988 23348 15997
rect 23572 16031 23624 16040
rect 23572 15997 23581 16031
rect 23581 15997 23615 16031
rect 23615 15997 23624 16031
rect 23572 15988 23624 15997
rect 24308 16124 24360 16176
rect 24032 16056 24084 16108
rect 20260 15852 20312 15904
rect 21088 15852 21140 15904
rect 21272 15852 21324 15904
rect 21548 15895 21600 15904
rect 21548 15861 21557 15895
rect 21557 15861 21591 15895
rect 21591 15861 21600 15895
rect 21548 15852 21600 15861
rect 21824 15895 21876 15904
rect 21824 15861 21833 15895
rect 21833 15861 21867 15895
rect 21867 15861 21876 15895
rect 21824 15852 21876 15861
rect 21916 15852 21968 15904
rect 22560 15852 22612 15904
rect 22836 15852 22888 15904
rect 25228 16056 25280 16108
rect 24308 15988 24360 16040
rect 26424 15988 26476 16040
rect 24124 15852 24176 15904
rect 26608 15852 26660 15904
rect 8102 15750 8154 15802
rect 8166 15750 8218 15802
rect 8230 15750 8282 15802
rect 8294 15750 8346 15802
rect 8358 15750 8410 15802
rect 15807 15750 15859 15802
rect 15871 15750 15923 15802
rect 15935 15750 15987 15802
rect 15999 15750 16051 15802
rect 16063 15750 16115 15802
rect 23512 15750 23564 15802
rect 23576 15750 23628 15802
rect 23640 15750 23692 15802
rect 23704 15750 23756 15802
rect 23768 15750 23820 15802
rect 31217 15750 31269 15802
rect 31281 15750 31333 15802
rect 31345 15750 31397 15802
rect 31409 15750 31461 15802
rect 31473 15750 31525 15802
rect 9772 15648 9824 15700
rect 9956 15648 10008 15700
rect 10324 15648 10376 15700
rect 10600 15648 10652 15700
rect 10876 15648 10928 15700
rect 8484 15444 8536 15496
rect 8944 15555 8996 15564
rect 8944 15521 8953 15555
rect 8953 15521 8987 15555
rect 8987 15521 8996 15555
rect 8944 15512 8996 15521
rect 9496 15555 9548 15564
rect 9496 15521 9505 15555
rect 9505 15521 9539 15555
rect 9539 15521 9548 15555
rect 9496 15512 9548 15521
rect 9680 15512 9732 15564
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 10324 15555 10376 15564
rect 10324 15521 10333 15555
rect 10333 15521 10367 15555
rect 10367 15521 10376 15555
rect 10324 15512 10376 15521
rect 11060 15580 11112 15632
rect 10692 15512 10744 15564
rect 11428 15648 11480 15700
rect 12624 15648 12676 15700
rect 14832 15648 14884 15700
rect 15476 15648 15528 15700
rect 15660 15648 15712 15700
rect 11888 15580 11940 15632
rect 11428 15555 11480 15564
rect 11428 15521 11437 15555
rect 11437 15521 11471 15555
rect 11471 15521 11480 15555
rect 11428 15512 11480 15521
rect 8576 15376 8628 15428
rect 9588 15376 9640 15428
rect 11060 15444 11112 15496
rect 11704 15512 11756 15564
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 8300 15308 8352 15360
rect 9128 15308 9180 15360
rect 10784 15376 10836 15428
rect 12164 15555 12216 15564
rect 12164 15521 12173 15555
rect 12173 15521 12207 15555
rect 12207 15521 12216 15555
rect 12164 15512 12216 15521
rect 12440 15555 12492 15564
rect 12440 15521 12449 15555
rect 12449 15521 12483 15555
rect 12483 15521 12492 15555
rect 12440 15512 12492 15521
rect 12900 15512 12952 15564
rect 12992 15512 13044 15564
rect 13268 15512 13320 15564
rect 13728 15555 13780 15564
rect 13728 15521 13737 15555
rect 13737 15521 13771 15555
rect 13771 15521 13780 15555
rect 13728 15512 13780 15521
rect 13912 15555 13964 15564
rect 13912 15521 13921 15555
rect 13921 15521 13955 15555
rect 13955 15521 13964 15555
rect 13912 15512 13964 15521
rect 14740 15580 14792 15632
rect 14280 15376 14332 15428
rect 11428 15308 11480 15360
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 14188 15308 14240 15360
rect 15476 15376 15528 15428
rect 16672 15553 16724 15564
rect 16672 15519 16681 15553
rect 16681 15519 16715 15553
rect 16715 15519 16724 15553
rect 16672 15512 16724 15519
rect 16856 15512 16908 15564
rect 17960 15512 18012 15564
rect 18328 15648 18380 15700
rect 18972 15648 19024 15700
rect 19064 15648 19116 15700
rect 19524 15648 19576 15700
rect 18420 15580 18472 15632
rect 18328 15555 18380 15564
rect 18328 15521 18337 15555
rect 18337 15521 18371 15555
rect 18371 15521 18380 15555
rect 18328 15512 18380 15521
rect 19064 15555 19116 15564
rect 19064 15521 19073 15555
rect 19073 15521 19107 15555
rect 19107 15521 19116 15555
rect 19064 15512 19116 15521
rect 18880 15444 18932 15496
rect 19432 15512 19484 15564
rect 19800 15623 19852 15632
rect 19800 15589 19809 15623
rect 19809 15589 19843 15623
rect 19843 15589 19852 15623
rect 19800 15580 19852 15589
rect 17500 15376 17552 15428
rect 16672 15308 16724 15360
rect 17316 15351 17368 15360
rect 17316 15317 17325 15351
rect 17325 15317 17359 15351
rect 17359 15317 17368 15351
rect 17316 15308 17368 15317
rect 18144 15351 18196 15360
rect 18144 15317 18153 15351
rect 18153 15317 18187 15351
rect 18187 15317 18196 15351
rect 18144 15308 18196 15317
rect 19064 15308 19116 15360
rect 19340 15376 19392 15428
rect 20076 15580 20128 15632
rect 20536 15648 20588 15700
rect 22100 15648 22152 15700
rect 22284 15648 22336 15700
rect 20720 15512 20772 15564
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 22468 15580 22520 15632
rect 21916 15555 21968 15564
rect 21916 15521 21925 15555
rect 21925 15521 21959 15555
rect 21959 15521 21968 15555
rect 21916 15512 21968 15521
rect 22008 15555 22060 15564
rect 22008 15521 22017 15555
rect 22017 15521 22051 15555
rect 22051 15521 22060 15555
rect 22008 15512 22060 15521
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 22376 15555 22428 15564
rect 22376 15521 22385 15555
rect 22385 15521 22419 15555
rect 22419 15521 22428 15555
rect 22376 15512 22428 15521
rect 22928 15648 22980 15700
rect 23296 15648 23348 15700
rect 24952 15691 25004 15700
rect 24952 15657 24961 15691
rect 24961 15657 24995 15691
rect 24995 15657 25004 15691
rect 24952 15648 25004 15657
rect 24032 15580 24084 15632
rect 24124 15623 24176 15632
rect 24124 15589 24133 15623
rect 24133 15589 24167 15623
rect 24167 15589 24176 15623
rect 24124 15580 24176 15589
rect 23296 15444 23348 15496
rect 23848 15444 23900 15496
rect 24216 15555 24268 15564
rect 24216 15521 24225 15555
rect 24225 15521 24259 15555
rect 24259 15521 24268 15555
rect 24216 15512 24268 15521
rect 25688 15580 25740 15632
rect 24584 15555 24636 15564
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 24860 15555 24912 15564
rect 24860 15521 24869 15555
rect 24869 15521 24903 15555
rect 24903 15521 24912 15555
rect 24860 15512 24912 15521
rect 26332 15444 26384 15496
rect 20996 15376 21048 15428
rect 22192 15419 22244 15428
rect 22192 15385 22201 15419
rect 22201 15385 22235 15419
rect 22235 15385 22244 15419
rect 22192 15376 22244 15385
rect 25320 15376 25372 15428
rect 19432 15308 19484 15360
rect 19524 15308 19576 15360
rect 20352 15308 20404 15360
rect 21180 15308 21232 15360
rect 21364 15351 21416 15360
rect 21364 15317 21373 15351
rect 21373 15317 21407 15351
rect 21407 15317 21416 15351
rect 21364 15308 21416 15317
rect 21640 15351 21692 15360
rect 21640 15317 21649 15351
rect 21649 15317 21683 15351
rect 21683 15317 21692 15351
rect 21640 15308 21692 15317
rect 22100 15308 22152 15360
rect 23480 15308 23532 15360
rect 24216 15308 24268 15360
rect 4250 15206 4302 15258
rect 4314 15206 4366 15258
rect 4378 15206 4430 15258
rect 4442 15206 4494 15258
rect 4506 15206 4558 15258
rect 11955 15206 12007 15258
rect 12019 15206 12071 15258
rect 12083 15206 12135 15258
rect 12147 15206 12199 15258
rect 12211 15206 12263 15258
rect 19660 15206 19712 15258
rect 19724 15206 19776 15258
rect 19788 15206 19840 15258
rect 19852 15206 19904 15258
rect 19916 15206 19968 15258
rect 27365 15206 27417 15258
rect 27429 15206 27481 15258
rect 27493 15206 27545 15258
rect 27557 15206 27609 15258
rect 27621 15206 27673 15258
rect 8668 15104 8720 15156
rect 9772 15104 9824 15156
rect 10232 15104 10284 15156
rect 10508 15104 10560 15156
rect 12716 15104 12768 15156
rect 13636 15147 13688 15156
rect 13636 15113 13645 15147
rect 13645 15113 13679 15147
rect 13679 15113 13688 15147
rect 13636 15104 13688 15113
rect 13728 15104 13780 15156
rect 13912 15104 13964 15156
rect 17408 15104 17460 15156
rect 18328 15104 18380 15156
rect 19340 15104 19392 15156
rect 8484 14900 8536 14952
rect 8760 14900 8812 14952
rect 9588 15011 9640 15020
rect 9588 14977 9597 15011
rect 9597 14977 9631 15011
rect 9631 14977 9640 15011
rect 9588 14968 9640 14977
rect 9312 14900 9364 14952
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 7196 14764 7248 14816
rect 8300 14764 8352 14816
rect 9312 14807 9364 14816
rect 9312 14773 9321 14807
rect 9321 14773 9355 14807
rect 9355 14773 9364 14807
rect 9312 14764 9364 14773
rect 9496 14832 9548 14884
rect 9956 14943 10008 14952
rect 9956 14909 9965 14943
rect 9965 14909 9999 14943
rect 9999 14909 10008 14943
rect 9956 14900 10008 14909
rect 18604 15036 18656 15088
rect 20812 15104 20864 15156
rect 20352 15036 20404 15088
rect 22192 15104 22244 15156
rect 22560 15104 22612 15156
rect 23940 15147 23992 15156
rect 23940 15113 23949 15147
rect 23949 15113 23983 15147
rect 23983 15113 23992 15147
rect 23940 15104 23992 15113
rect 24216 15104 24268 15156
rect 28264 15104 28316 15156
rect 23204 15079 23256 15088
rect 23204 15045 23213 15079
rect 23213 15045 23247 15079
rect 23247 15045 23256 15079
rect 23204 15036 23256 15045
rect 10140 14900 10192 14952
rect 10324 14900 10376 14952
rect 10692 14900 10744 14952
rect 11520 14900 11572 14952
rect 11612 14900 11664 14952
rect 9772 14764 9824 14816
rect 10968 14832 11020 14884
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 10600 14764 10652 14816
rect 11336 14764 11388 14816
rect 11796 14832 11848 14884
rect 13084 14943 13136 14952
rect 13084 14909 13093 14943
rect 13093 14909 13127 14943
rect 13127 14909 13136 14943
rect 13084 14900 13136 14909
rect 13820 14900 13872 14952
rect 17776 14900 17828 14952
rect 18144 14900 18196 14952
rect 20260 14900 20312 14952
rect 25044 15079 25096 15088
rect 25044 15045 25053 15079
rect 25053 15045 25087 15079
rect 25087 15045 25096 15079
rect 25044 15036 25096 15045
rect 25136 15036 25188 15088
rect 23480 14968 23532 15020
rect 23388 14943 23440 14952
rect 23388 14909 23397 14943
rect 23397 14909 23431 14943
rect 23431 14909 23440 14943
rect 23388 14900 23440 14909
rect 23756 14900 23808 14952
rect 14004 14832 14056 14884
rect 15568 14832 15620 14884
rect 17132 14832 17184 14884
rect 12992 14764 13044 14816
rect 13176 14807 13228 14816
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 13544 14764 13596 14816
rect 14280 14764 14332 14816
rect 15200 14764 15252 14816
rect 21732 14832 21784 14884
rect 23020 14832 23072 14884
rect 21180 14764 21232 14816
rect 22652 14764 22704 14816
rect 23388 14764 23440 14816
rect 24124 14900 24176 14952
rect 24492 14943 24544 14952
rect 24492 14909 24501 14943
rect 24501 14909 24535 14943
rect 24535 14909 24544 14943
rect 24492 14900 24544 14909
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 24768 14900 24820 14952
rect 25228 14943 25280 14952
rect 25228 14909 25237 14943
rect 25237 14909 25271 14943
rect 25271 14909 25280 14943
rect 25228 14900 25280 14909
rect 25872 14832 25924 14884
rect 24400 14764 24452 14816
rect 24952 14764 25004 14816
rect 25504 14764 25556 14816
rect 25780 14764 25832 14816
rect 28264 14764 28316 14816
rect 29644 14764 29696 14816
rect 31668 14764 31720 14816
rect 8102 14662 8154 14714
rect 8166 14662 8218 14714
rect 8230 14662 8282 14714
rect 8294 14662 8346 14714
rect 8358 14662 8410 14714
rect 15807 14662 15859 14714
rect 15871 14662 15923 14714
rect 15935 14662 15987 14714
rect 15999 14662 16051 14714
rect 16063 14662 16115 14714
rect 23512 14662 23564 14714
rect 23576 14662 23628 14714
rect 23640 14662 23692 14714
rect 23704 14662 23756 14714
rect 23768 14662 23820 14714
rect 31217 14662 31269 14714
rect 31281 14662 31333 14714
rect 31345 14662 31397 14714
rect 31409 14662 31461 14714
rect 31473 14662 31525 14714
rect 7840 14560 7892 14612
rect 7932 14603 7984 14612
rect 7932 14569 7941 14603
rect 7941 14569 7975 14603
rect 7975 14569 7984 14603
rect 7932 14560 7984 14569
rect 7564 14492 7616 14544
rect 8944 14560 8996 14612
rect 10232 14560 10284 14612
rect 10692 14560 10744 14612
rect 11336 14560 11388 14612
rect 13084 14560 13136 14612
rect 15476 14560 15528 14612
rect 16212 14560 16264 14612
rect 16672 14560 16724 14612
rect 16856 14560 16908 14612
rect 17316 14560 17368 14612
rect 19064 14560 19116 14612
rect 19156 14560 19208 14612
rect 7840 14467 7892 14476
rect 7840 14433 7849 14467
rect 7849 14433 7883 14467
rect 7883 14433 7892 14467
rect 7840 14424 7892 14433
rect 8024 14467 8076 14476
rect 8024 14433 8033 14467
rect 8033 14433 8067 14467
rect 8067 14433 8076 14467
rect 8024 14424 8076 14433
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 8668 14467 8720 14476
rect 8668 14433 8677 14467
rect 8677 14433 8711 14467
rect 8711 14433 8720 14467
rect 8668 14424 8720 14433
rect 8300 14288 8352 14340
rect 11060 14492 11112 14544
rect 9128 14467 9180 14476
rect 9128 14433 9137 14467
rect 9137 14433 9171 14467
rect 9171 14433 9180 14467
rect 9128 14424 9180 14433
rect 9772 14424 9824 14476
rect 15200 14492 15252 14544
rect 8852 14356 8904 14408
rect 8944 14356 8996 14408
rect 10876 14356 10928 14408
rect 13268 14424 13320 14476
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 12808 14356 12860 14408
rect 13820 14467 13872 14476
rect 13820 14433 13829 14467
rect 13829 14433 13863 14467
rect 13863 14433 13872 14467
rect 13820 14424 13872 14433
rect 14188 14424 14240 14476
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 14648 14467 14700 14476
rect 14648 14433 14682 14467
rect 14682 14433 14700 14467
rect 14648 14424 14700 14433
rect 14004 14356 14056 14408
rect 16396 14467 16448 14476
rect 16396 14433 16405 14467
rect 16405 14433 16439 14467
rect 16439 14433 16448 14467
rect 16396 14424 16448 14433
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 16948 14424 17000 14433
rect 18420 14492 18472 14544
rect 17960 14467 18012 14476
rect 17960 14433 17969 14467
rect 17969 14433 18003 14467
rect 18003 14433 18012 14467
rect 17960 14424 18012 14433
rect 18052 14467 18104 14476
rect 18052 14433 18061 14467
rect 18061 14433 18095 14467
rect 18095 14433 18104 14467
rect 18052 14424 18104 14433
rect 18328 14424 18380 14476
rect 7104 14220 7156 14272
rect 8024 14220 8076 14272
rect 11612 14288 11664 14340
rect 13544 14288 13596 14340
rect 13820 14288 13872 14340
rect 18328 14288 18380 14340
rect 18604 14356 18656 14408
rect 19432 14467 19484 14476
rect 19432 14433 19441 14467
rect 19441 14433 19475 14467
rect 19475 14433 19484 14467
rect 19432 14424 19484 14433
rect 19524 14424 19576 14476
rect 21088 14560 21140 14612
rect 21732 14560 21784 14612
rect 22100 14560 22152 14612
rect 20720 14492 20772 14544
rect 18788 14288 18840 14340
rect 21548 14467 21600 14476
rect 21548 14433 21557 14467
rect 21557 14433 21591 14467
rect 21591 14433 21600 14467
rect 21548 14424 21600 14433
rect 21824 14424 21876 14476
rect 22100 14356 22152 14408
rect 20720 14288 20772 14340
rect 21732 14288 21784 14340
rect 22560 14560 22612 14612
rect 22836 14560 22888 14612
rect 23112 14492 23164 14544
rect 24032 14603 24084 14612
rect 24032 14569 24041 14603
rect 24041 14569 24075 14603
rect 24075 14569 24084 14603
rect 24032 14560 24084 14569
rect 24124 14560 24176 14612
rect 24308 14560 24360 14612
rect 24584 14560 24636 14612
rect 25688 14603 25740 14612
rect 25688 14569 25697 14603
rect 25697 14569 25731 14603
rect 25731 14569 25740 14603
rect 25688 14560 25740 14569
rect 25780 14560 25832 14612
rect 23940 14424 23992 14476
rect 24124 14467 24176 14476
rect 24124 14433 24133 14467
rect 24133 14433 24167 14467
rect 24167 14433 24176 14467
rect 24124 14424 24176 14433
rect 24400 14424 24452 14476
rect 24952 14465 25004 14476
rect 24952 14431 24961 14465
rect 24961 14431 24995 14465
rect 24995 14431 25004 14465
rect 24952 14424 25004 14431
rect 25504 14467 25556 14476
rect 25504 14433 25513 14467
rect 25513 14433 25547 14467
rect 25547 14433 25556 14467
rect 25504 14424 25556 14433
rect 25780 14467 25832 14476
rect 25780 14433 25789 14467
rect 25789 14433 25823 14467
rect 25823 14433 25832 14467
rect 25780 14424 25832 14433
rect 8484 14263 8536 14272
rect 8484 14229 8493 14263
rect 8493 14229 8527 14263
rect 8527 14229 8536 14263
rect 8484 14220 8536 14229
rect 9496 14220 9548 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 13728 14220 13780 14272
rect 16212 14263 16264 14272
rect 16212 14229 16221 14263
rect 16221 14229 16255 14263
rect 16255 14229 16264 14263
rect 16212 14220 16264 14229
rect 17316 14263 17368 14272
rect 17316 14229 17325 14263
rect 17325 14229 17359 14263
rect 17359 14229 17368 14263
rect 17316 14220 17368 14229
rect 17500 14220 17552 14272
rect 18420 14263 18472 14272
rect 18420 14229 18429 14263
rect 18429 14229 18463 14263
rect 18463 14229 18472 14263
rect 18420 14220 18472 14229
rect 18512 14220 18564 14272
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 20352 14263 20404 14272
rect 20352 14229 20361 14263
rect 20361 14229 20395 14263
rect 20395 14229 20404 14263
rect 20352 14220 20404 14229
rect 20444 14220 20496 14272
rect 21180 14220 21232 14272
rect 21456 14220 21508 14272
rect 24814 14356 24866 14408
rect 25688 14356 25740 14408
rect 22376 14220 22428 14272
rect 24216 14220 24268 14272
rect 24584 14263 24636 14272
rect 24584 14229 24593 14263
rect 24593 14229 24627 14263
rect 24627 14229 24636 14263
rect 24584 14220 24636 14229
rect 24952 14288 25004 14340
rect 25136 14263 25188 14272
rect 25136 14229 25145 14263
rect 25145 14229 25179 14263
rect 25179 14229 25188 14263
rect 25136 14220 25188 14229
rect 4250 14118 4302 14170
rect 4314 14118 4366 14170
rect 4378 14118 4430 14170
rect 4442 14118 4494 14170
rect 4506 14118 4558 14170
rect 11955 14118 12007 14170
rect 12019 14118 12071 14170
rect 12083 14118 12135 14170
rect 12147 14118 12199 14170
rect 12211 14118 12263 14170
rect 19660 14118 19712 14170
rect 19724 14118 19776 14170
rect 19788 14118 19840 14170
rect 19852 14118 19904 14170
rect 19916 14118 19968 14170
rect 27365 14118 27417 14170
rect 27429 14118 27481 14170
rect 27493 14118 27545 14170
rect 27557 14118 27609 14170
rect 27621 14118 27673 14170
rect 7840 14016 7892 14068
rect 7932 14016 7984 14068
rect 8576 14016 8628 14068
rect 7196 13948 7248 14000
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 7472 13880 7524 13932
rect 8116 13880 8168 13932
rect 8300 13880 8352 13932
rect 8944 14016 8996 14068
rect 9772 14016 9824 14068
rect 9864 14016 9916 14068
rect 10232 14016 10284 14068
rect 10140 13948 10192 14000
rect 10508 13991 10560 14000
rect 10508 13957 10517 13991
rect 10517 13957 10551 13991
rect 10551 13957 10560 13991
rect 10508 13948 10560 13957
rect 10784 13948 10836 14000
rect 11704 14016 11756 14068
rect 11796 13948 11848 14000
rect 13452 13948 13504 14000
rect 13912 13948 13964 14000
rect 7380 13849 7432 13864
rect 7380 13815 7397 13849
rect 7397 13815 7431 13849
rect 7431 13815 7432 13849
rect 7380 13812 7432 13815
rect 7656 13855 7708 13864
rect 7656 13821 7665 13855
rect 7665 13821 7699 13855
rect 7699 13821 7708 13855
rect 7656 13812 7708 13821
rect 7932 13855 7984 13864
rect 7932 13821 7941 13855
rect 7941 13821 7975 13855
rect 7975 13821 7984 13855
rect 7932 13812 7984 13821
rect 8208 13812 8260 13864
rect 7564 13744 7616 13796
rect 8576 13812 8628 13864
rect 8760 13812 8812 13864
rect 9312 13812 9364 13864
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 10876 13812 10928 13864
rect 10140 13744 10192 13796
rect 11888 13880 11940 13932
rect 12348 13880 12400 13932
rect 11612 13812 11664 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 13544 13880 13596 13932
rect 14188 14016 14240 14068
rect 17316 14016 17368 14068
rect 17960 14016 18012 14068
rect 18052 14016 18104 14068
rect 19248 14016 19300 14068
rect 20720 14016 20772 14068
rect 12164 13744 12216 13796
rect 12992 13812 13044 13864
rect 13728 13812 13780 13864
rect 9220 13676 9272 13728
rect 10048 13676 10100 13728
rect 11520 13676 11572 13728
rect 12624 13676 12676 13728
rect 13636 13744 13688 13796
rect 14464 13744 14516 13796
rect 14648 13812 14700 13864
rect 15292 13812 15344 13864
rect 16396 13948 16448 14000
rect 19524 13948 19576 14000
rect 15936 13855 15988 13864
rect 15936 13821 15945 13855
rect 15945 13821 15979 13855
rect 15979 13821 15988 13855
rect 15936 13812 15988 13821
rect 18788 13880 18840 13932
rect 23756 14016 23808 14068
rect 23848 14016 23900 14068
rect 25136 14016 25188 14068
rect 25320 14059 25372 14068
rect 25320 14025 25329 14059
rect 25329 14025 25363 14059
rect 25363 14025 25372 14059
rect 25320 14016 25372 14025
rect 25596 14059 25648 14068
rect 25596 14025 25605 14059
rect 25605 14025 25639 14059
rect 25639 14025 25648 14059
rect 25596 14016 25648 14025
rect 26148 14059 26200 14068
rect 26148 14025 26157 14059
rect 26157 14025 26191 14059
rect 26191 14025 26200 14059
rect 26148 14016 26200 14025
rect 26424 14059 26476 14068
rect 26424 14025 26433 14059
rect 26433 14025 26467 14059
rect 26467 14025 26476 14059
rect 26424 14016 26476 14025
rect 23480 13948 23532 14000
rect 24768 13948 24820 14000
rect 17224 13855 17276 13864
rect 17224 13821 17233 13855
rect 17233 13821 17267 13855
rect 17267 13821 17276 13855
rect 17224 13812 17276 13821
rect 17684 13855 17736 13864
rect 17684 13821 17693 13855
rect 17693 13821 17727 13855
rect 17727 13821 17736 13855
rect 17684 13812 17736 13821
rect 18052 13812 18104 13864
rect 18236 13855 18288 13864
rect 18236 13821 18245 13855
rect 18245 13821 18279 13855
rect 18279 13821 18288 13855
rect 18236 13812 18288 13821
rect 18328 13855 18380 13864
rect 18328 13821 18337 13855
rect 18337 13821 18371 13855
rect 18371 13821 18380 13855
rect 18328 13812 18380 13821
rect 13912 13676 13964 13728
rect 14740 13676 14792 13728
rect 16396 13744 16448 13796
rect 16948 13744 17000 13796
rect 20260 13744 20312 13796
rect 20996 13812 21048 13864
rect 21456 13880 21508 13932
rect 25228 13948 25280 14000
rect 21732 13812 21784 13864
rect 21456 13744 21508 13796
rect 22192 13855 22244 13864
rect 22192 13821 22201 13855
rect 22201 13821 22235 13855
rect 22235 13821 22244 13855
rect 22192 13812 22244 13821
rect 22284 13812 22336 13864
rect 23296 13812 23348 13864
rect 24216 13744 24268 13796
rect 15476 13676 15528 13728
rect 17132 13676 17184 13728
rect 19340 13676 19392 13728
rect 21732 13719 21784 13728
rect 21732 13685 21741 13719
rect 21741 13685 21775 13719
rect 21775 13685 21784 13719
rect 21732 13676 21784 13685
rect 22008 13719 22060 13728
rect 22008 13685 22017 13719
rect 22017 13685 22051 13719
rect 22051 13685 22060 13719
rect 22008 13676 22060 13685
rect 22100 13676 22152 13728
rect 24400 13812 24452 13864
rect 24492 13812 24544 13864
rect 24860 13855 24912 13864
rect 24860 13821 24869 13855
rect 24869 13821 24903 13855
rect 24903 13821 24912 13855
rect 24860 13812 24912 13821
rect 25596 13812 25648 13864
rect 25872 13812 25924 13864
rect 26332 13855 26384 13864
rect 26332 13821 26341 13855
rect 26341 13821 26375 13855
rect 26375 13821 26384 13855
rect 26332 13812 26384 13821
rect 26608 13855 26660 13864
rect 26608 13821 26617 13855
rect 26617 13821 26651 13855
rect 26651 13821 26660 13855
rect 26608 13812 26660 13821
rect 25412 13676 25464 13728
rect 25688 13676 25740 13728
rect 26700 13719 26752 13728
rect 26700 13685 26709 13719
rect 26709 13685 26743 13719
rect 26743 13685 26752 13719
rect 26700 13676 26752 13685
rect 8102 13574 8154 13626
rect 8166 13574 8218 13626
rect 8230 13574 8282 13626
rect 8294 13574 8346 13626
rect 8358 13574 8410 13626
rect 15807 13574 15859 13626
rect 15871 13574 15923 13626
rect 15935 13574 15987 13626
rect 15999 13574 16051 13626
rect 16063 13574 16115 13626
rect 23512 13574 23564 13626
rect 23576 13574 23628 13626
rect 23640 13574 23692 13626
rect 23704 13574 23756 13626
rect 23768 13574 23820 13626
rect 31217 13574 31269 13626
rect 31281 13574 31333 13626
rect 31345 13574 31397 13626
rect 31409 13574 31461 13626
rect 31473 13574 31525 13626
rect 7932 13472 7984 13524
rect 8392 13472 8444 13524
rect 8484 13472 8536 13524
rect 8668 13472 8720 13524
rect 7656 13404 7708 13456
rect 7932 13336 7984 13388
rect 8116 13379 8168 13388
rect 8116 13345 8125 13379
rect 8125 13345 8159 13379
rect 8159 13345 8168 13379
rect 8116 13336 8168 13345
rect 8024 13200 8076 13252
rect 9128 13404 9180 13456
rect 9220 13379 9272 13388
rect 9220 13345 9229 13379
rect 9229 13345 9263 13379
rect 9263 13345 9272 13379
rect 9220 13336 9272 13345
rect 9588 13515 9640 13524
rect 9588 13481 9597 13515
rect 9597 13481 9631 13515
rect 9631 13481 9640 13515
rect 9588 13472 9640 13481
rect 10140 13515 10192 13524
rect 10140 13481 10149 13515
rect 10149 13481 10183 13515
rect 10183 13481 10192 13515
rect 10140 13472 10192 13481
rect 10692 13472 10744 13524
rect 11060 13472 11112 13524
rect 12532 13472 12584 13524
rect 13360 13515 13412 13524
rect 13360 13481 13369 13515
rect 13369 13481 13403 13515
rect 13403 13481 13412 13515
rect 13360 13472 13412 13481
rect 13912 13472 13964 13524
rect 15660 13472 15712 13524
rect 16764 13472 16816 13524
rect 18052 13472 18104 13524
rect 18420 13472 18472 13524
rect 19064 13515 19116 13524
rect 19064 13481 19073 13515
rect 19073 13481 19107 13515
rect 19107 13481 19116 13515
rect 19064 13472 19116 13481
rect 20536 13472 20588 13524
rect 21548 13472 21600 13524
rect 22008 13472 22060 13524
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 10508 13336 10560 13388
rect 12256 13447 12308 13456
rect 11612 13379 11664 13388
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 11612 13336 11664 13345
rect 12256 13413 12290 13447
rect 12290 13413 12308 13447
rect 12256 13404 12308 13413
rect 17592 13404 17644 13456
rect 12716 13336 12768 13388
rect 13820 13379 13872 13388
rect 13820 13345 13829 13379
rect 13829 13345 13863 13379
rect 13863 13345 13872 13379
rect 13820 13336 13872 13345
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 7748 13132 7800 13184
rect 8116 13132 8168 13184
rect 9864 13175 9916 13184
rect 9864 13141 9873 13175
rect 9873 13141 9907 13175
rect 9907 13141 9916 13175
rect 9864 13132 9916 13141
rect 11244 13200 11296 13252
rect 16212 13336 16264 13388
rect 17776 13336 17828 13388
rect 17960 13379 18012 13388
rect 17960 13345 17994 13379
rect 17994 13345 18012 13379
rect 17960 13336 18012 13345
rect 20352 13404 20404 13456
rect 14004 13268 14056 13320
rect 14648 13268 14700 13320
rect 21456 13336 21508 13388
rect 21088 13268 21140 13320
rect 21272 13268 21324 13320
rect 21732 13336 21784 13388
rect 23204 13472 23256 13524
rect 22560 13404 22612 13456
rect 23664 13336 23716 13388
rect 21824 13268 21876 13320
rect 22192 13311 22244 13320
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 24216 13404 24268 13456
rect 24584 13404 24636 13456
rect 25320 13515 25372 13524
rect 25320 13481 25329 13515
rect 25329 13481 25363 13515
rect 25363 13481 25372 13515
rect 25320 13472 25372 13481
rect 25412 13472 25464 13524
rect 25964 13515 26016 13524
rect 25964 13481 25973 13515
rect 25973 13481 26007 13515
rect 26007 13481 26016 13515
rect 25964 13472 26016 13481
rect 26424 13472 26476 13524
rect 31668 13472 31720 13524
rect 24492 13336 24544 13388
rect 24860 13336 24912 13388
rect 25780 13404 25832 13456
rect 25504 13379 25556 13388
rect 25504 13345 25513 13379
rect 25513 13345 25547 13379
rect 25547 13345 25556 13379
rect 25504 13336 25556 13345
rect 25688 13336 25740 13388
rect 13912 13200 13964 13252
rect 11336 13132 11388 13184
rect 11520 13175 11572 13184
rect 11520 13141 11529 13175
rect 11529 13141 11563 13175
rect 11563 13141 11572 13175
rect 11520 13132 11572 13141
rect 11612 13132 11664 13184
rect 12992 13132 13044 13184
rect 14280 13132 14332 13184
rect 15476 13132 15528 13184
rect 21916 13200 21968 13252
rect 16856 13132 16908 13184
rect 20720 13132 20772 13184
rect 20904 13175 20956 13184
rect 20904 13141 20913 13175
rect 20913 13141 20947 13175
rect 20947 13141 20956 13175
rect 20904 13132 20956 13141
rect 21456 13175 21508 13184
rect 21456 13141 21465 13175
rect 21465 13141 21499 13175
rect 21499 13141 21508 13175
rect 21456 13132 21508 13141
rect 25964 13268 26016 13320
rect 26424 13132 26476 13184
rect 26516 13175 26568 13184
rect 26516 13141 26525 13175
rect 26525 13141 26559 13175
rect 26559 13141 26568 13175
rect 26516 13132 26568 13141
rect 28264 13132 28316 13184
rect 4250 13030 4302 13082
rect 4314 13030 4366 13082
rect 4378 13030 4430 13082
rect 4442 13030 4494 13082
rect 4506 13030 4558 13082
rect 11955 13030 12007 13082
rect 12019 13030 12071 13082
rect 12083 13030 12135 13082
rect 12147 13030 12199 13082
rect 12211 13030 12263 13082
rect 19660 13030 19712 13082
rect 19724 13030 19776 13082
rect 19788 13030 19840 13082
rect 19852 13030 19904 13082
rect 19916 13030 19968 13082
rect 27365 13030 27417 13082
rect 27429 13030 27481 13082
rect 27493 13030 27545 13082
rect 27557 13030 27609 13082
rect 27621 13030 27673 13082
rect 7564 12971 7616 12980
rect 7564 12937 7573 12971
rect 7573 12937 7607 12971
rect 7607 12937 7616 12971
rect 7564 12928 7616 12937
rect 7748 12928 7800 12980
rect 8944 12971 8996 12980
rect 8944 12937 8953 12971
rect 8953 12937 8987 12971
rect 8987 12937 8996 12971
rect 8944 12928 8996 12937
rect 9404 12928 9456 12980
rect 10968 12928 11020 12980
rect 13452 12928 13504 12980
rect 15384 12928 15436 12980
rect 16856 12928 16908 12980
rect 17684 12928 17736 12980
rect 18144 12928 18196 12980
rect 20168 12928 20220 12980
rect 24492 12971 24544 12980
rect 24492 12937 24501 12971
rect 24501 12937 24535 12971
rect 24535 12937 24544 12971
rect 24492 12928 24544 12937
rect 24676 12928 24728 12980
rect 25872 12928 25924 12980
rect 9036 12860 9088 12912
rect 8852 12792 8904 12844
rect 8116 12724 8168 12776
rect 8392 12724 8444 12776
rect 11060 12860 11112 12912
rect 12624 12860 12676 12912
rect 13636 12860 13688 12912
rect 15292 12860 15344 12912
rect 21364 12860 21416 12912
rect 10600 12792 10652 12844
rect 21088 12792 21140 12844
rect 9772 12724 9824 12776
rect 8760 12656 8812 12708
rect 9128 12656 9180 12708
rect 10416 12767 10468 12776
rect 10416 12733 10425 12767
rect 10425 12733 10459 12767
rect 10459 12733 10468 12767
rect 10416 12724 10468 12733
rect 11244 12724 11296 12776
rect 11152 12656 11204 12708
rect 11612 12656 11664 12708
rect 8484 12588 8536 12640
rect 9404 12588 9456 12640
rect 10140 12588 10192 12640
rect 12716 12767 12768 12776
rect 12716 12733 12725 12767
rect 12725 12733 12759 12767
rect 12759 12733 12768 12767
rect 12716 12724 12768 12733
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 13176 12767 13228 12776
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 15200 12767 15252 12776
rect 15200 12733 15209 12767
rect 15209 12733 15243 12767
rect 15243 12733 15252 12767
rect 15200 12724 15252 12733
rect 16948 12724 17000 12776
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 17776 12724 17828 12776
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 20996 12767 21048 12776
rect 20996 12733 21005 12767
rect 21005 12733 21039 12767
rect 21039 12733 21048 12767
rect 20996 12724 21048 12733
rect 12992 12656 13044 12708
rect 14004 12656 14056 12708
rect 17132 12656 17184 12708
rect 20812 12656 20864 12708
rect 21364 12724 21416 12776
rect 21548 12767 21600 12776
rect 21548 12733 21557 12767
rect 21557 12733 21591 12767
rect 21591 12733 21600 12767
rect 21548 12724 21600 12733
rect 21824 12767 21876 12776
rect 21824 12733 21833 12767
rect 21833 12733 21867 12767
rect 21867 12733 21876 12767
rect 21824 12724 21876 12733
rect 22652 12792 22704 12844
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 23848 12724 23900 12733
rect 23940 12767 23992 12776
rect 23940 12733 23949 12767
rect 23949 12733 23983 12767
rect 23983 12733 23992 12767
rect 23940 12724 23992 12733
rect 24032 12724 24084 12776
rect 24308 12767 24360 12776
rect 24308 12733 24317 12767
rect 24317 12733 24351 12767
rect 24351 12733 24360 12767
rect 24308 12724 24360 12733
rect 12624 12588 12676 12640
rect 13268 12631 13320 12640
rect 13268 12597 13277 12631
rect 13277 12597 13311 12631
rect 13311 12597 13320 12631
rect 13268 12588 13320 12597
rect 21088 12588 21140 12640
rect 24860 12860 24912 12912
rect 24952 12767 25004 12776
rect 24952 12733 24961 12767
rect 24961 12733 24995 12767
rect 24995 12733 25004 12767
rect 24952 12724 25004 12733
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 25780 12792 25832 12844
rect 26332 12767 26384 12776
rect 26332 12733 26341 12767
rect 26341 12733 26375 12767
rect 26375 12733 26384 12767
rect 26332 12724 26384 12733
rect 21640 12588 21692 12640
rect 22376 12588 22428 12640
rect 26056 12656 26108 12708
rect 24308 12588 24360 12640
rect 24400 12588 24452 12640
rect 8102 12486 8154 12538
rect 8166 12486 8218 12538
rect 8230 12486 8282 12538
rect 8294 12486 8346 12538
rect 8358 12486 8410 12538
rect 15807 12486 15859 12538
rect 15871 12486 15923 12538
rect 15935 12486 15987 12538
rect 15999 12486 16051 12538
rect 16063 12486 16115 12538
rect 23512 12486 23564 12538
rect 23576 12486 23628 12538
rect 23640 12486 23692 12538
rect 23704 12486 23756 12538
rect 23768 12486 23820 12538
rect 31217 12486 31269 12538
rect 31281 12486 31333 12538
rect 31345 12486 31397 12538
rect 31409 12486 31461 12538
rect 31473 12486 31525 12538
rect 8484 12427 8536 12436
rect 8484 12393 8493 12427
rect 8493 12393 8527 12427
rect 8527 12393 8536 12427
rect 8484 12384 8536 12393
rect 8576 12384 8628 12436
rect 8760 12427 8812 12436
rect 8760 12393 8769 12427
rect 8769 12393 8803 12427
rect 8803 12393 8812 12427
rect 8760 12384 8812 12393
rect 8852 12384 8904 12436
rect 9404 12384 9456 12436
rect 9864 12384 9916 12436
rect 10048 12384 10100 12436
rect 10232 12427 10284 12436
rect 10232 12393 10241 12427
rect 10241 12393 10275 12427
rect 10275 12393 10284 12427
rect 10232 12384 10284 12393
rect 11244 12384 11296 12436
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 11980 12427 12032 12436
rect 11980 12393 11989 12427
rect 11989 12393 12023 12427
rect 12023 12393 12032 12427
rect 11980 12384 12032 12393
rect 12716 12384 12768 12436
rect 7380 12248 7432 12300
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 8668 12180 8720 12232
rect 9220 12248 9272 12300
rect 9404 12291 9456 12300
rect 9404 12257 9412 12291
rect 9412 12257 9456 12291
rect 9404 12248 9456 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 10784 12316 10836 12368
rect 12992 12384 13044 12436
rect 13176 12384 13228 12436
rect 13360 12384 13412 12436
rect 10324 12291 10376 12300
rect 10324 12257 10333 12291
rect 10333 12257 10367 12291
rect 10367 12257 10376 12291
rect 10324 12248 10376 12257
rect 11060 12291 11112 12300
rect 11060 12257 11069 12291
rect 11069 12257 11103 12291
rect 11103 12257 11112 12291
rect 11060 12248 11112 12257
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 11612 12291 11664 12300
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 13176 12248 13228 12300
rect 13268 12291 13320 12300
rect 13268 12257 13277 12291
rect 13277 12257 13311 12291
rect 13311 12257 13320 12291
rect 13268 12248 13320 12257
rect 12808 12180 12860 12232
rect 14188 12316 14240 12368
rect 14280 12316 14332 12368
rect 13912 12248 13964 12300
rect 14096 12248 14148 12300
rect 17776 12384 17828 12436
rect 21640 12384 21692 12436
rect 21732 12384 21784 12436
rect 24400 12384 24452 12436
rect 28264 12384 28316 12436
rect 15476 12316 15528 12368
rect 14740 12248 14792 12300
rect 12900 12112 12952 12164
rect 8944 12044 8996 12096
rect 9220 12044 9272 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 13820 12112 13872 12164
rect 13452 12044 13504 12096
rect 13912 12087 13964 12096
rect 13912 12053 13921 12087
rect 13921 12053 13955 12087
rect 13955 12053 13964 12087
rect 13912 12044 13964 12053
rect 15200 12291 15252 12300
rect 15200 12257 15209 12291
rect 15209 12257 15243 12291
rect 15243 12257 15252 12291
rect 15200 12248 15252 12257
rect 15016 12180 15068 12232
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 15752 12291 15804 12300
rect 15752 12257 15761 12291
rect 15761 12257 15795 12291
rect 15795 12257 15804 12291
rect 15752 12248 15804 12257
rect 15844 12291 15896 12300
rect 15844 12257 15853 12291
rect 15853 12257 15887 12291
rect 15887 12257 15896 12291
rect 15844 12248 15896 12257
rect 15108 12112 15160 12164
rect 18604 12316 18656 12368
rect 17592 12291 17644 12300
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 26056 12316 26108 12368
rect 26148 12359 26200 12368
rect 26148 12325 26157 12359
rect 26157 12325 26191 12359
rect 26191 12325 26200 12359
rect 26148 12316 26200 12325
rect 17592 12248 17644 12257
rect 16304 12112 16356 12164
rect 17132 12112 17184 12164
rect 19524 12248 19576 12300
rect 20628 12291 20680 12300
rect 20628 12257 20637 12291
rect 20637 12257 20671 12291
rect 20671 12257 20680 12291
rect 20628 12248 20680 12257
rect 20720 12291 20772 12300
rect 20720 12257 20729 12291
rect 20729 12257 20763 12291
rect 20763 12257 20772 12291
rect 20720 12248 20772 12257
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 21548 12248 21600 12300
rect 24492 12248 24544 12300
rect 24584 12248 24636 12300
rect 24768 12291 24820 12300
rect 24768 12257 24777 12291
rect 24777 12257 24811 12291
rect 24811 12257 24820 12291
rect 24768 12248 24820 12257
rect 26516 12316 26568 12368
rect 15016 12044 15068 12096
rect 15568 12044 15620 12096
rect 16488 12087 16540 12096
rect 16488 12053 16497 12087
rect 16497 12053 16531 12087
rect 16531 12053 16540 12087
rect 16488 12044 16540 12053
rect 16856 12044 16908 12096
rect 18880 12112 18932 12164
rect 20904 12112 20956 12164
rect 18052 12044 18104 12096
rect 19524 12087 19576 12096
rect 19524 12053 19533 12087
rect 19533 12053 19567 12087
rect 19567 12053 19576 12087
rect 19524 12044 19576 12053
rect 20076 12087 20128 12096
rect 20076 12053 20085 12087
rect 20085 12053 20119 12087
rect 20119 12053 20128 12087
rect 20076 12044 20128 12053
rect 20536 12087 20588 12096
rect 20536 12053 20545 12087
rect 20545 12053 20579 12087
rect 20579 12053 20588 12087
rect 20536 12044 20588 12053
rect 22192 12044 22244 12096
rect 26332 12248 26384 12300
rect 24676 12112 24728 12164
rect 24492 12044 24544 12096
rect 25596 12087 25648 12096
rect 25596 12053 25605 12087
rect 25605 12053 25639 12087
rect 25639 12053 25648 12087
rect 25596 12044 25648 12053
rect 4250 11942 4302 11994
rect 4314 11942 4366 11994
rect 4378 11942 4430 11994
rect 4442 11942 4494 11994
rect 4506 11942 4558 11994
rect 11955 11942 12007 11994
rect 12019 11942 12071 11994
rect 12083 11942 12135 11994
rect 12147 11942 12199 11994
rect 12211 11942 12263 11994
rect 19660 11942 19712 11994
rect 19724 11942 19776 11994
rect 19788 11942 19840 11994
rect 19852 11942 19904 11994
rect 19916 11942 19968 11994
rect 27365 11942 27417 11994
rect 27429 11942 27481 11994
rect 27493 11942 27545 11994
rect 27557 11942 27609 11994
rect 27621 11942 27673 11994
rect 7748 11679 7800 11688
rect 7748 11645 7792 11679
rect 7792 11645 7800 11679
rect 7748 11636 7800 11645
rect 9220 11840 9272 11892
rect 10692 11840 10744 11892
rect 9404 11704 9456 11756
rect 9036 11636 9088 11688
rect 9680 11679 9732 11688
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 9680 11636 9732 11645
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 10048 11679 10100 11688
rect 10048 11645 10057 11679
rect 10057 11645 10091 11679
rect 10091 11645 10100 11679
rect 10048 11636 10100 11645
rect 11336 11840 11388 11892
rect 11704 11883 11756 11892
rect 11704 11849 11713 11883
rect 11713 11849 11747 11883
rect 11747 11849 11756 11883
rect 11704 11840 11756 11849
rect 13912 11840 13964 11892
rect 15200 11840 15252 11892
rect 15476 11840 15528 11892
rect 15660 11840 15712 11892
rect 14004 11704 14056 11756
rect 14096 11704 14148 11756
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 14924 11772 14976 11824
rect 17224 11840 17276 11892
rect 18512 11840 18564 11892
rect 20352 11840 20404 11892
rect 20536 11883 20588 11892
rect 20536 11849 20545 11883
rect 20545 11849 20579 11883
rect 20579 11849 20588 11883
rect 20536 11840 20588 11849
rect 20628 11840 20680 11892
rect 21088 11883 21140 11892
rect 21088 11849 21097 11883
rect 21097 11849 21131 11883
rect 21131 11849 21140 11883
rect 21088 11840 21140 11849
rect 13544 11568 13596 11620
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 15016 11679 15068 11688
rect 15016 11645 15025 11679
rect 15025 11645 15059 11679
rect 15059 11645 15068 11679
rect 15660 11747 15712 11756
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 15016 11636 15068 11645
rect 15476 11681 15528 11688
rect 15476 11647 15485 11681
rect 15485 11647 15519 11681
rect 15519 11647 15528 11681
rect 15476 11636 15528 11647
rect 15844 11636 15896 11688
rect 15292 11568 15344 11620
rect 9496 11500 9548 11552
rect 9588 11543 9640 11552
rect 9588 11509 9597 11543
rect 9597 11509 9631 11543
rect 9631 11509 9640 11543
rect 9588 11500 9640 11509
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 14832 11543 14884 11552
rect 14832 11509 14841 11543
rect 14841 11509 14875 11543
rect 14875 11509 14884 11543
rect 14832 11500 14884 11509
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 15476 11500 15528 11552
rect 16672 11772 16724 11824
rect 17040 11704 17092 11756
rect 18880 11704 18932 11756
rect 24768 11883 24820 11892
rect 24768 11849 24777 11883
rect 24777 11849 24811 11883
rect 24811 11849 24820 11883
rect 24768 11840 24820 11849
rect 21272 11772 21324 11824
rect 25504 11840 25556 11892
rect 25596 11840 25648 11892
rect 19708 11636 19760 11688
rect 20996 11636 21048 11688
rect 21548 11636 21600 11688
rect 21640 11636 21692 11688
rect 21824 11679 21876 11688
rect 21824 11645 21833 11679
rect 21833 11645 21867 11679
rect 21867 11645 21876 11679
rect 21824 11636 21876 11645
rect 22192 11679 22244 11688
rect 22192 11645 22201 11679
rect 22201 11645 22235 11679
rect 22235 11645 22244 11679
rect 22192 11636 22244 11645
rect 24308 11679 24360 11688
rect 24308 11645 24317 11679
rect 24317 11645 24351 11679
rect 24351 11645 24360 11679
rect 24308 11636 24360 11645
rect 24492 11636 24544 11688
rect 16672 11500 16724 11552
rect 19984 11500 20036 11552
rect 21548 11500 21600 11552
rect 24032 11568 24084 11620
rect 24124 11500 24176 11552
rect 24216 11543 24268 11552
rect 24216 11509 24225 11543
rect 24225 11509 24259 11543
rect 24259 11509 24268 11543
rect 24216 11500 24268 11509
rect 24676 11679 24728 11688
rect 24676 11645 24685 11679
rect 24685 11645 24719 11679
rect 24719 11645 24728 11679
rect 24676 11636 24728 11645
rect 25044 11636 25096 11688
rect 25964 11636 26016 11688
rect 25136 11500 25188 11552
rect 25412 11500 25464 11552
rect 25872 11568 25924 11620
rect 8102 11398 8154 11450
rect 8166 11398 8218 11450
rect 8230 11398 8282 11450
rect 8294 11398 8346 11450
rect 8358 11398 8410 11450
rect 15807 11398 15859 11450
rect 15871 11398 15923 11450
rect 15935 11398 15987 11450
rect 15999 11398 16051 11450
rect 16063 11398 16115 11450
rect 23512 11398 23564 11450
rect 23576 11398 23628 11450
rect 23640 11398 23692 11450
rect 23704 11398 23756 11450
rect 23768 11398 23820 11450
rect 31217 11398 31269 11450
rect 31281 11398 31333 11450
rect 31345 11398 31397 11450
rect 31409 11398 31461 11450
rect 31473 11398 31525 11450
rect 7748 11296 7800 11348
rect 10048 11296 10100 11348
rect 8116 11203 8168 11212
rect 8116 11169 8125 11203
rect 8125 11169 8159 11203
rect 8159 11169 8168 11203
rect 8116 11160 8168 11169
rect 6184 11092 6236 11144
rect 8484 11160 8536 11212
rect 10140 11228 10192 11280
rect 11612 11339 11664 11348
rect 11612 11305 11621 11339
rect 11621 11305 11655 11339
rect 11655 11305 11664 11339
rect 11612 11296 11664 11305
rect 12440 11296 12492 11348
rect 14372 11296 14424 11348
rect 15568 11296 15620 11348
rect 16304 11296 16356 11348
rect 16488 11296 16540 11348
rect 17224 11296 17276 11348
rect 18052 11296 18104 11348
rect 18236 11339 18288 11348
rect 18236 11305 18245 11339
rect 18245 11305 18279 11339
rect 18279 11305 18288 11339
rect 18236 11296 18288 11305
rect 19432 11339 19484 11348
rect 19432 11305 19441 11339
rect 19441 11305 19475 11339
rect 19475 11305 19484 11339
rect 19432 11296 19484 11305
rect 19524 11296 19576 11348
rect 19708 11339 19760 11348
rect 19708 11305 19717 11339
rect 19717 11305 19751 11339
rect 19751 11305 19760 11339
rect 19708 11296 19760 11305
rect 20076 11296 20128 11348
rect 8576 11092 8628 11144
rect 9220 11092 9272 11144
rect 10416 11092 10468 11144
rect 8944 11024 8996 11076
rect 9956 11024 10008 11076
rect 12532 11092 12584 11144
rect 11336 11067 11388 11076
rect 11336 11033 11345 11067
rect 11345 11033 11379 11067
rect 11379 11033 11388 11067
rect 11336 11024 11388 11033
rect 11612 11024 11664 11076
rect 11704 11024 11756 11076
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 9128 10956 9180 11008
rect 10140 10999 10192 11008
rect 10140 10965 10149 10999
rect 10149 10965 10183 10999
rect 10183 10965 10192 10999
rect 10140 10956 10192 10965
rect 10324 10956 10376 11008
rect 10692 10999 10744 11008
rect 10692 10965 10701 10999
rect 10701 10965 10735 10999
rect 10735 10965 10744 10999
rect 10692 10956 10744 10965
rect 11060 10999 11112 11008
rect 11060 10965 11069 10999
rect 11069 10965 11103 10999
rect 11103 10965 11112 10999
rect 11060 10956 11112 10965
rect 11244 10956 11296 11008
rect 13452 11203 13504 11212
rect 13452 11169 13475 11203
rect 13475 11169 13504 11203
rect 13452 11160 13504 11169
rect 14004 11160 14056 11212
rect 15292 11160 15344 11212
rect 15384 11203 15436 11212
rect 15384 11169 15393 11203
rect 15393 11169 15427 11203
rect 15427 11169 15436 11203
rect 15384 11160 15436 11169
rect 16120 11203 16172 11212
rect 16120 11169 16129 11203
rect 16129 11169 16163 11203
rect 16163 11169 16172 11203
rect 16120 11160 16172 11169
rect 16488 11160 16540 11212
rect 16856 11092 16908 11144
rect 12992 10999 13044 11008
rect 12992 10965 13001 10999
rect 13001 10965 13035 10999
rect 13035 10965 13044 10999
rect 12992 10956 13044 10965
rect 15476 11024 15528 11076
rect 14096 10956 14148 11008
rect 15844 10999 15896 11008
rect 15844 10965 15853 10999
rect 15853 10965 15887 10999
rect 15887 10965 15896 10999
rect 15844 10956 15896 10965
rect 16948 11024 17000 11076
rect 17776 11024 17828 11076
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 24216 11296 24268 11348
rect 24400 11296 24452 11348
rect 25044 11296 25096 11348
rect 25412 11296 25464 11348
rect 20260 11203 20312 11212
rect 20260 11169 20269 11203
rect 20269 11169 20303 11203
rect 20303 11169 20312 11203
rect 20996 11271 21048 11280
rect 20996 11237 21005 11271
rect 21005 11237 21039 11271
rect 21039 11237 21048 11271
rect 20996 11228 21048 11237
rect 21732 11228 21784 11280
rect 23296 11271 23348 11280
rect 23296 11237 23305 11271
rect 23305 11237 23339 11271
rect 23339 11237 23348 11271
rect 23296 11228 23348 11237
rect 20260 11160 20312 11169
rect 20720 11092 20772 11144
rect 21548 11160 21600 11212
rect 22192 11160 22244 11212
rect 23572 11160 23624 11212
rect 23848 11228 23900 11280
rect 24124 11228 24176 11280
rect 28264 11228 28316 11280
rect 24216 11160 24268 11212
rect 24492 11203 24544 11212
rect 24492 11169 24501 11203
rect 24501 11169 24535 11203
rect 24535 11169 24544 11203
rect 24492 11160 24544 11169
rect 24676 11160 24728 11212
rect 25228 11203 25280 11212
rect 25228 11169 25237 11203
rect 25237 11169 25271 11203
rect 25271 11169 25280 11203
rect 25228 11160 25280 11169
rect 25136 11092 25188 11144
rect 16764 10956 16816 11008
rect 17132 10956 17184 11008
rect 19340 11024 19392 11076
rect 21456 11024 21508 11076
rect 21548 11024 21600 11076
rect 23940 11024 23992 11076
rect 18052 10999 18104 11008
rect 18052 10965 18061 10999
rect 18061 10965 18095 10999
rect 18095 10965 18104 10999
rect 18052 10956 18104 10965
rect 18604 10999 18656 11008
rect 18604 10965 18613 10999
rect 18613 10965 18647 10999
rect 18647 10965 18656 10999
rect 18604 10956 18656 10965
rect 18880 10999 18932 11008
rect 18880 10965 18889 10999
rect 18889 10965 18923 10999
rect 18923 10965 18932 10999
rect 18880 10956 18932 10965
rect 21180 10956 21232 11008
rect 21640 10956 21692 11008
rect 23480 10999 23532 11008
rect 23480 10965 23489 10999
rect 23489 10965 23523 10999
rect 23523 10965 23532 10999
rect 23480 10956 23532 10965
rect 24032 10999 24084 11008
rect 24032 10965 24041 10999
rect 24041 10965 24075 10999
rect 24075 10965 24084 10999
rect 24032 10956 24084 10965
rect 24308 10999 24360 11008
rect 24308 10965 24317 10999
rect 24317 10965 24351 10999
rect 24351 10965 24360 10999
rect 24308 10956 24360 10965
rect 24584 10999 24636 11008
rect 24584 10965 24593 10999
rect 24593 10965 24627 10999
rect 24627 10965 24636 10999
rect 24584 10956 24636 10965
rect 24860 10999 24912 11008
rect 24860 10965 24869 10999
rect 24869 10965 24903 10999
rect 24903 10965 24912 10999
rect 24860 10956 24912 10965
rect 24952 10956 25004 11008
rect 25320 10956 25372 11008
rect 4250 10854 4302 10906
rect 4314 10854 4366 10906
rect 4378 10854 4430 10906
rect 4442 10854 4494 10906
rect 4506 10854 4558 10906
rect 11955 10854 12007 10906
rect 12019 10854 12071 10906
rect 12083 10854 12135 10906
rect 12147 10854 12199 10906
rect 12211 10854 12263 10906
rect 19660 10854 19712 10906
rect 19724 10854 19776 10906
rect 19788 10854 19840 10906
rect 19852 10854 19904 10906
rect 19916 10854 19968 10906
rect 27365 10854 27417 10906
rect 27429 10854 27481 10906
rect 27493 10854 27545 10906
rect 27557 10854 27609 10906
rect 27621 10854 27673 10906
rect 8116 10752 8168 10804
rect 8944 10752 8996 10804
rect 9128 10752 9180 10804
rect 11520 10752 11572 10804
rect 13268 10795 13320 10804
rect 13268 10761 13277 10795
rect 13277 10761 13311 10795
rect 13311 10761 13320 10795
rect 13268 10752 13320 10761
rect 15844 10752 15896 10804
rect 16212 10752 16264 10804
rect 16580 10752 16632 10804
rect 16856 10795 16908 10804
rect 16856 10761 16865 10795
rect 16865 10761 16899 10795
rect 16899 10761 16908 10795
rect 16856 10752 16908 10761
rect 19340 10795 19392 10804
rect 19340 10761 19349 10795
rect 19349 10761 19383 10795
rect 19383 10761 19392 10795
rect 19340 10752 19392 10761
rect 20904 10752 20956 10804
rect 24032 10752 24084 10804
rect 24676 10752 24728 10804
rect 24860 10752 24912 10804
rect 25228 10752 25280 10804
rect 7656 10548 7708 10600
rect 8024 10548 8076 10600
rect 8484 10616 8536 10668
rect 9680 10684 9732 10736
rect 8760 10548 8812 10600
rect 9220 10548 9272 10600
rect 9864 10548 9916 10600
rect 10692 10684 10744 10736
rect 19432 10684 19484 10736
rect 10140 10548 10192 10600
rect 11152 10548 11204 10600
rect 13820 10591 13872 10600
rect 13820 10557 13829 10591
rect 13829 10557 13863 10591
rect 13863 10557 13872 10591
rect 13820 10548 13872 10557
rect 14004 10548 14056 10600
rect 15660 10548 15712 10600
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 17132 10548 17184 10600
rect 18052 10548 18104 10600
rect 18880 10548 18932 10600
rect 9772 10480 9824 10532
rect 7840 10455 7892 10464
rect 7840 10421 7849 10455
rect 7849 10421 7883 10455
rect 7883 10421 7892 10455
rect 7840 10412 7892 10421
rect 8024 10412 8076 10464
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 9036 10455 9088 10464
rect 9036 10421 9045 10455
rect 9045 10421 9079 10455
rect 9079 10421 9088 10455
rect 9036 10412 9088 10421
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 10232 10412 10284 10464
rect 11520 10523 11572 10532
rect 11520 10489 11538 10523
rect 11538 10489 11572 10523
rect 11520 10480 11572 10489
rect 13360 10480 13412 10532
rect 15108 10480 15160 10532
rect 13728 10455 13780 10464
rect 13728 10421 13737 10455
rect 13737 10421 13771 10455
rect 13771 10421 13780 10455
rect 13728 10412 13780 10421
rect 16212 10412 16264 10464
rect 16672 10412 16724 10464
rect 17132 10412 17184 10464
rect 18144 10412 18196 10464
rect 20260 10548 20312 10600
rect 20352 10591 20404 10600
rect 20352 10557 20361 10591
rect 20361 10557 20395 10591
rect 20395 10557 20404 10591
rect 20352 10548 20404 10557
rect 19892 10455 19944 10464
rect 19892 10421 19901 10455
rect 19901 10421 19935 10455
rect 19935 10421 19944 10455
rect 19892 10412 19944 10421
rect 20720 10591 20772 10600
rect 20720 10557 20729 10591
rect 20729 10557 20763 10591
rect 20763 10557 20772 10591
rect 20720 10548 20772 10557
rect 21180 10591 21232 10600
rect 21180 10557 21189 10591
rect 21189 10557 21223 10591
rect 21223 10557 21232 10591
rect 21180 10548 21232 10557
rect 21364 10480 21416 10532
rect 21548 10548 21600 10600
rect 28264 10684 28316 10736
rect 22100 10548 22152 10600
rect 21916 10480 21968 10532
rect 23480 10548 23532 10600
rect 24308 10591 24360 10600
rect 24308 10557 24317 10591
rect 24317 10557 24351 10591
rect 24351 10557 24360 10591
rect 24308 10548 24360 10557
rect 24492 10616 24544 10668
rect 24584 10548 24636 10600
rect 25320 10548 25372 10600
rect 25688 10591 25740 10600
rect 25688 10557 25697 10591
rect 25697 10557 25731 10591
rect 25731 10557 25740 10591
rect 25688 10548 25740 10557
rect 21272 10412 21324 10464
rect 23572 10412 23624 10464
rect 24032 10412 24084 10464
rect 24216 10412 24268 10464
rect 31668 10412 31720 10464
rect 8102 10310 8154 10362
rect 8166 10310 8218 10362
rect 8230 10310 8282 10362
rect 8294 10310 8346 10362
rect 8358 10310 8410 10362
rect 15807 10310 15859 10362
rect 15871 10310 15923 10362
rect 15935 10310 15987 10362
rect 15999 10310 16051 10362
rect 16063 10310 16115 10362
rect 23512 10310 23564 10362
rect 23576 10310 23628 10362
rect 23640 10310 23692 10362
rect 23704 10310 23756 10362
rect 23768 10310 23820 10362
rect 31217 10310 31269 10362
rect 31281 10310 31333 10362
rect 31345 10310 31397 10362
rect 31409 10310 31461 10362
rect 31473 10310 31525 10362
rect 7932 10208 7984 10260
rect 8024 10251 8076 10260
rect 8024 10217 8033 10251
rect 8033 10217 8067 10251
rect 8067 10217 8076 10251
rect 8024 10208 8076 10217
rect 8576 10208 8628 10260
rect 8760 10208 8812 10260
rect 9036 10208 9088 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 9588 10208 9640 10260
rect 9864 10208 9916 10260
rect 11060 10208 11112 10260
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 12992 10208 13044 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 13728 10208 13780 10260
rect 13820 10208 13872 10260
rect 15200 10208 15252 10260
rect 15292 10208 15344 10260
rect 16212 10208 16264 10260
rect 16764 10251 16816 10260
rect 16764 10217 16773 10251
rect 16773 10217 16807 10251
rect 16807 10217 16816 10251
rect 16764 10208 16816 10217
rect 18696 10208 18748 10260
rect 19892 10208 19944 10260
rect 20352 10208 20404 10260
rect 28264 10208 28316 10260
rect 7196 10072 7248 10124
rect 7380 10115 7432 10124
rect 7380 10081 7389 10115
rect 7389 10081 7423 10115
rect 7423 10081 7432 10115
rect 7380 10072 7432 10081
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 8484 10072 8536 10124
rect 8668 10115 8720 10124
rect 8668 10081 8677 10115
rect 8677 10081 8711 10115
rect 8711 10081 8720 10115
rect 8668 10072 8720 10081
rect 9312 10072 9364 10124
rect 11612 10140 11664 10192
rect 6736 9936 6788 9988
rect 7840 9936 7892 9988
rect 11152 10072 11204 10124
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 11704 10072 11756 10124
rect 12348 10072 12400 10124
rect 13084 10004 13136 10056
rect 13912 10072 13964 10124
rect 14096 10115 14148 10124
rect 14096 10081 14105 10115
rect 14105 10081 14139 10115
rect 14139 10081 14148 10115
rect 14096 10072 14148 10081
rect 14372 10115 14424 10124
rect 14372 10081 14381 10115
rect 14381 10081 14415 10115
rect 14415 10081 14424 10115
rect 14372 10072 14424 10081
rect 14648 10072 14700 10124
rect 15108 10072 15160 10124
rect 15016 10004 15068 10056
rect 15568 10072 15620 10124
rect 13820 9936 13872 9988
rect 15844 10047 15896 10056
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 17040 10072 17092 10124
rect 17132 10115 17184 10124
rect 17132 10081 17141 10115
rect 17141 10081 17175 10115
rect 17175 10081 17184 10115
rect 17132 10072 17184 10081
rect 17316 10072 17368 10124
rect 18604 10072 18656 10124
rect 6644 9868 6696 9920
rect 7288 9868 7340 9920
rect 7472 9911 7524 9920
rect 7472 9877 7481 9911
rect 7481 9877 7515 9911
rect 7515 9877 7524 9911
rect 7472 9868 7524 9877
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 8300 9911 8352 9920
rect 8300 9877 8309 9911
rect 8309 9877 8343 9911
rect 8343 9877 8352 9911
rect 8300 9868 8352 9877
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 8668 9868 8720 9920
rect 9864 9868 9916 9920
rect 10324 9868 10376 9920
rect 11060 9868 11112 9920
rect 11704 9911 11756 9920
rect 11704 9877 11713 9911
rect 11713 9877 11747 9911
rect 11747 9877 11756 9911
rect 11704 9868 11756 9877
rect 11796 9868 11848 9920
rect 12900 9868 12952 9920
rect 12992 9868 13044 9920
rect 13912 9868 13964 9920
rect 14740 9911 14792 9920
rect 14740 9877 14749 9911
rect 14749 9877 14783 9911
rect 14783 9877 14792 9911
rect 14740 9868 14792 9877
rect 15752 9936 15804 9988
rect 15292 9911 15344 9920
rect 15292 9877 15301 9911
rect 15301 9877 15335 9911
rect 15335 9877 15344 9911
rect 15292 9868 15344 9877
rect 15384 9868 15436 9920
rect 16488 9911 16540 9920
rect 16488 9877 16497 9911
rect 16497 9877 16531 9911
rect 16531 9877 16540 9911
rect 16488 9868 16540 9877
rect 20168 9911 20220 9920
rect 20168 9877 20177 9911
rect 20177 9877 20211 9911
rect 20211 9877 20220 9911
rect 20168 9868 20220 9877
rect 20904 10183 20956 10192
rect 20904 10149 20913 10183
rect 20913 10149 20947 10183
rect 20947 10149 20956 10183
rect 20904 10140 20956 10149
rect 21272 10140 21324 10192
rect 21364 10115 21416 10124
rect 21364 10081 21373 10115
rect 21373 10081 21407 10115
rect 21407 10081 21416 10115
rect 21364 10072 21416 10081
rect 21732 10072 21784 10124
rect 21916 10072 21968 10124
rect 23388 10140 23440 10192
rect 24032 10115 24084 10124
rect 24032 10081 24041 10115
rect 24041 10081 24075 10115
rect 24075 10081 24084 10115
rect 24032 10072 24084 10081
rect 24952 10140 25004 10192
rect 24768 10072 24820 10124
rect 25044 10072 25096 10124
rect 25136 10115 25188 10124
rect 25136 10081 25145 10115
rect 25145 10081 25179 10115
rect 25179 10081 25188 10115
rect 25136 10072 25188 10081
rect 25320 10115 25372 10124
rect 25320 10081 25329 10115
rect 25329 10081 25363 10115
rect 25363 10081 25372 10115
rect 25320 10072 25372 10081
rect 26148 10140 26200 10192
rect 22100 9936 22152 9988
rect 26056 10004 26108 10056
rect 24860 9936 24912 9988
rect 25964 9936 26016 9988
rect 21364 9868 21416 9920
rect 21916 9868 21968 9920
rect 24308 9868 24360 9920
rect 24400 9911 24452 9920
rect 24400 9877 24409 9911
rect 24409 9877 24443 9911
rect 24443 9877 24452 9911
rect 24400 9868 24452 9877
rect 24676 9911 24728 9920
rect 24676 9877 24685 9911
rect 24685 9877 24719 9911
rect 24719 9877 24728 9911
rect 24676 9868 24728 9877
rect 25228 9911 25280 9920
rect 25228 9877 25237 9911
rect 25237 9877 25271 9911
rect 25271 9877 25280 9911
rect 25228 9868 25280 9877
rect 25504 9911 25556 9920
rect 25504 9877 25513 9911
rect 25513 9877 25547 9911
rect 25547 9877 25556 9911
rect 25504 9868 25556 9877
rect 26240 9868 26292 9920
rect 4250 9766 4302 9818
rect 4314 9766 4366 9818
rect 4378 9766 4430 9818
rect 4442 9766 4494 9818
rect 4506 9766 4558 9818
rect 11955 9766 12007 9818
rect 12019 9766 12071 9818
rect 12083 9766 12135 9818
rect 12147 9766 12199 9818
rect 12211 9766 12263 9818
rect 19660 9766 19712 9818
rect 19724 9766 19776 9818
rect 19788 9766 19840 9818
rect 19852 9766 19904 9818
rect 19916 9766 19968 9818
rect 27365 9766 27417 9818
rect 27429 9766 27481 9818
rect 27493 9766 27545 9818
rect 27557 9766 27609 9818
rect 27621 9766 27673 9818
rect 6184 9639 6236 9648
rect 6184 9605 6193 9639
rect 6193 9605 6227 9639
rect 6227 9605 6236 9639
rect 6184 9596 6236 9605
rect 6460 9503 6512 9512
rect 6460 9469 6469 9503
rect 6469 9469 6503 9503
rect 6503 9469 6512 9503
rect 6460 9460 6512 9469
rect 6736 9460 6788 9512
rect 7196 9664 7248 9716
rect 7472 9664 7524 9716
rect 7564 9664 7616 9716
rect 7380 9596 7432 9648
rect 9680 9664 9732 9716
rect 9772 9664 9824 9716
rect 8300 9596 8352 9648
rect 8668 9639 8720 9648
rect 8668 9605 8677 9639
rect 8677 9605 8711 9639
rect 8711 9605 8720 9639
rect 8668 9596 8720 9605
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 7288 9392 7340 9444
rect 7932 9503 7984 9512
rect 7932 9469 7949 9503
rect 7949 9469 7983 9503
rect 7983 9469 7984 9503
rect 7932 9460 7984 9469
rect 10692 9596 10744 9648
rect 11612 9664 11664 9716
rect 11704 9664 11756 9716
rect 11796 9664 11848 9716
rect 11336 9596 11388 9648
rect 11888 9639 11940 9648
rect 11888 9605 11897 9639
rect 11897 9605 11931 9639
rect 11931 9605 11940 9639
rect 11888 9596 11940 9605
rect 8484 9460 8536 9512
rect 8024 9392 8076 9444
rect 8576 9392 8628 9444
rect 6736 9367 6788 9376
rect 6736 9333 6745 9367
rect 6745 9333 6779 9367
rect 6779 9333 6788 9367
rect 6736 9324 6788 9333
rect 8760 9324 8812 9376
rect 9128 9324 9180 9376
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10048 9460 10100 9469
rect 9772 9435 9824 9444
rect 9772 9401 9790 9435
rect 9790 9401 9824 9435
rect 11060 9460 11112 9512
rect 11520 9503 11572 9512
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 11888 9460 11940 9512
rect 12348 9596 12400 9648
rect 12992 9528 13044 9580
rect 12624 9460 12676 9512
rect 13912 9707 13964 9716
rect 13912 9673 13921 9707
rect 13921 9673 13955 9707
rect 13955 9673 13964 9707
rect 13912 9664 13964 9673
rect 14372 9664 14424 9716
rect 14648 9596 14700 9648
rect 13912 9528 13964 9580
rect 9772 9392 9824 9401
rect 10232 9367 10284 9376
rect 10232 9333 10241 9367
rect 10241 9333 10275 9367
rect 10275 9333 10284 9367
rect 10232 9324 10284 9333
rect 10324 9324 10376 9376
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 11704 9367 11756 9376
rect 11704 9333 11713 9367
rect 11713 9333 11747 9367
rect 11747 9333 11756 9367
rect 11704 9324 11756 9333
rect 12900 9324 12952 9376
rect 13360 9324 13412 9376
rect 13728 9503 13780 9512
rect 13728 9469 13737 9503
rect 13737 9469 13771 9503
rect 13771 9469 13780 9503
rect 13728 9460 13780 9469
rect 14096 9503 14148 9512
rect 14096 9469 14105 9503
rect 14105 9469 14139 9503
rect 14139 9469 14148 9503
rect 14096 9460 14148 9469
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 14740 9460 14792 9512
rect 15568 9664 15620 9716
rect 20168 9664 20220 9716
rect 24216 9664 24268 9716
rect 24400 9664 24452 9716
rect 24676 9664 24728 9716
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 15752 9460 15804 9512
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 15200 9392 15252 9444
rect 16948 9392 17000 9444
rect 17592 9596 17644 9648
rect 17960 9639 18012 9648
rect 17960 9605 17969 9639
rect 17969 9605 18003 9639
rect 18003 9605 18012 9639
rect 17960 9596 18012 9605
rect 17868 9528 17920 9580
rect 23296 9596 23348 9648
rect 25136 9664 25188 9716
rect 25320 9664 25372 9716
rect 25688 9664 25740 9716
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 18236 9460 18288 9512
rect 19432 9460 19484 9512
rect 21364 9503 21416 9512
rect 21364 9469 21373 9503
rect 21373 9469 21407 9503
rect 21407 9469 21416 9503
rect 21364 9460 21416 9469
rect 21640 9503 21692 9512
rect 21640 9469 21649 9503
rect 21649 9469 21683 9503
rect 21683 9469 21692 9503
rect 21640 9460 21692 9469
rect 21732 9460 21784 9512
rect 21916 9503 21968 9512
rect 21916 9469 21925 9503
rect 21925 9469 21959 9503
rect 21959 9469 21968 9503
rect 21916 9460 21968 9469
rect 21088 9392 21140 9444
rect 15568 9324 15620 9376
rect 20076 9367 20128 9376
rect 20076 9333 20085 9367
rect 20085 9333 20119 9367
rect 20119 9333 20128 9367
rect 20076 9324 20128 9333
rect 20720 9324 20772 9376
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 21548 9367 21600 9376
rect 21548 9333 21557 9367
rect 21557 9333 21591 9367
rect 21591 9333 21600 9367
rect 21548 9324 21600 9333
rect 23848 9503 23900 9512
rect 23848 9469 23857 9503
rect 23857 9469 23891 9503
rect 23891 9469 23900 9503
rect 23848 9460 23900 9469
rect 22100 9392 22152 9444
rect 22192 9392 22244 9444
rect 24308 9460 24360 9512
rect 23940 9367 23992 9376
rect 23940 9333 23949 9367
rect 23949 9333 23983 9367
rect 23983 9333 23992 9367
rect 23940 9324 23992 9333
rect 24032 9324 24084 9376
rect 24584 9460 24636 9512
rect 25320 9503 25372 9512
rect 25320 9469 25329 9503
rect 25329 9469 25363 9503
rect 25363 9469 25372 9503
rect 25320 9460 25372 9469
rect 26056 9596 26108 9648
rect 26148 9596 26200 9648
rect 24768 9392 24820 9444
rect 25872 9503 25924 9512
rect 25872 9469 25881 9503
rect 25881 9469 25915 9503
rect 25915 9469 25924 9503
rect 25872 9460 25924 9469
rect 26240 9460 26292 9512
rect 26240 9324 26292 9376
rect 26976 9367 27028 9376
rect 26976 9333 26985 9367
rect 26985 9333 27019 9367
rect 27019 9333 27028 9367
rect 26976 9324 27028 9333
rect 8102 9222 8154 9274
rect 8166 9222 8218 9274
rect 8230 9222 8282 9274
rect 8294 9222 8346 9274
rect 8358 9222 8410 9274
rect 15807 9222 15859 9274
rect 15871 9222 15923 9274
rect 15935 9222 15987 9274
rect 15999 9222 16051 9274
rect 16063 9222 16115 9274
rect 23512 9222 23564 9274
rect 23576 9222 23628 9274
rect 23640 9222 23692 9274
rect 23704 9222 23756 9274
rect 23768 9222 23820 9274
rect 31217 9222 31269 9274
rect 31281 9222 31333 9274
rect 31345 9222 31397 9274
rect 31409 9222 31461 9274
rect 31473 9222 31525 9274
rect 6644 9163 6696 9172
rect 6644 9129 6653 9163
rect 6653 9129 6687 9163
rect 6687 9129 6696 9163
rect 6644 9120 6696 9129
rect 6736 9120 6788 9172
rect 7748 9120 7800 9172
rect 8392 9120 8444 9172
rect 7104 9052 7156 9104
rect 10232 9120 10284 9172
rect 10416 9163 10468 9172
rect 10416 9129 10425 9163
rect 10425 9129 10459 9163
rect 10459 9129 10468 9163
rect 10416 9120 10468 9129
rect 10508 9120 10560 9172
rect 10692 9163 10744 9172
rect 10692 9129 10701 9163
rect 10701 9129 10735 9163
rect 10735 9129 10744 9163
rect 10692 9120 10744 9129
rect 11704 9120 11756 9172
rect 13268 9120 13320 9172
rect 8760 9052 8812 9104
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7932 8984 7984 9036
rect 8116 9027 8168 9036
rect 8116 8993 8125 9027
rect 8125 8993 8159 9027
rect 8159 8993 8168 9027
rect 8116 8984 8168 8993
rect 8576 8984 8628 9036
rect 10140 9052 10192 9104
rect 7380 8916 7432 8925
rect 8300 8916 8352 8968
rect 9772 8984 9824 9036
rect 10324 8984 10376 9036
rect 11888 9052 11940 9104
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 13084 8984 13136 9036
rect 8576 8848 8628 8900
rect 10876 8916 10928 8968
rect 9680 8848 9732 8900
rect 11520 8848 11572 8900
rect 13544 9120 13596 9172
rect 13728 9120 13780 9172
rect 13912 9120 13964 9172
rect 15292 9120 15344 9172
rect 15660 9120 15712 9172
rect 16488 9120 16540 9172
rect 17316 9120 17368 9172
rect 15108 9027 15160 9036
rect 15108 8993 15117 9027
rect 15117 8993 15151 9027
rect 15151 8993 15160 9027
rect 15108 8984 15160 8993
rect 8024 8780 8076 8832
rect 8484 8823 8536 8832
rect 8484 8789 8493 8823
rect 8493 8789 8527 8823
rect 8527 8789 8536 8823
rect 8484 8780 8536 8789
rect 8760 8823 8812 8832
rect 8760 8789 8769 8823
rect 8769 8789 8803 8823
rect 8803 8789 8812 8823
rect 8760 8780 8812 8789
rect 8944 8780 8996 8832
rect 9036 8823 9088 8832
rect 9036 8789 9045 8823
rect 9045 8789 9079 8823
rect 9079 8789 9088 8823
rect 9036 8780 9088 8789
rect 9588 8823 9640 8832
rect 9588 8789 9597 8823
rect 9597 8789 9631 8823
rect 9631 8789 9640 8823
rect 9588 8780 9640 8789
rect 9772 8780 9824 8832
rect 9956 8780 10008 8832
rect 10324 8780 10376 8832
rect 13176 8780 13228 8832
rect 15016 8916 15068 8968
rect 15568 8984 15620 9036
rect 17776 9052 17828 9104
rect 18052 9163 18104 9172
rect 18052 9129 18061 9163
rect 18061 9129 18095 9163
rect 18095 9129 18104 9163
rect 18052 9120 18104 9129
rect 21088 9163 21140 9172
rect 21088 9129 21097 9163
rect 21097 9129 21131 9163
rect 21131 9129 21140 9163
rect 21088 9120 21140 9129
rect 21548 9120 21600 9172
rect 22192 9120 22244 9172
rect 16948 8984 17000 9036
rect 18144 9027 18196 9036
rect 18144 8993 18153 9027
rect 18153 8993 18187 9027
rect 18187 8993 18196 9027
rect 18144 8984 18196 8993
rect 20996 9052 21048 9104
rect 23848 9120 23900 9172
rect 23940 9120 23992 9172
rect 25044 9120 25096 9172
rect 25320 9120 25372 9172
rect 25872 9120 25924 9172
rect 25964 9163 26016 9172
rect 25964 9129 25973 9163
rect 25973 9129 26007 9163
rect 26007 9129 26016 9163
rect 25964 9120 26016 9129
rect 26976 9120 27028 9172
rect 22376 9095 22428 9104
rect 22376 9061 22385 9095
rect 22385 9061 22419 9095
rect 22419 9061 22428 9095
rect 22376 9052 22428 9061
rect 23480 9052 23532 9104
rect 24860 9052 24912 9104
rect 18788 8959 18840 8968
rect 18788 8925 18797 8959
rect 18797 8925 18831 8959
rect 18831 8925 18840 8959
rect 18788 8916 18840 8925
rect 20812 8916 20864 8968
rect 21272 9027 21324 9036
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 21272 8984 21324 8993
rect 21732 8984 21784 9036
rect 21916 8916 21968 8968
rect 20260 8848 20312 8900
rect 21640 8848 21692 8900
rect 22192 8984 22244 9036
rect 22928 8916 22980 8968
rect 26056 9027 26108 9036
rect 26056 8993 26065 9027
rect 26065 8993 26099 9027
rect 26099 8993 26108 9027
rect 26056 8984 26108 8993
rect 25412 8848 25464 8900
rect 26240 8848 26292 8900
rect 14096 8780 14148 8832
rect 14464 8780 14516 8832
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 15568 8823 15620 8832
rect 15568 8789 15577 8823
rect 15577 8789 15611 8823
rect 15611 8789 15620 8823
rect 15568 8780 15620 8789
rect 18328 8823 18380 8832
rect 18328 8789 18337 8823
rect 18337 8789 18371 8823
rect 18371 8789 18380 8823
rect 18328 8780 18380 8789
rect 20168 8780 20220 8832
rect 20352 8823 20404 8832
rect 20352 8789 20361 8823
rect 20361 8789 20395 8823
rect 20395 8789 20404 8823
rect 20352 8780 20404 8789
rect 21180 8780 21232 8832
rect 23020 8780 23072 8832
rect 23848 8823 23900 8832
rect 23848 8789 23857 8823
rect 23857 8789 23891 8823
rect 23891 8789 23900 8823
rect 23848 8780 23900 8789
rect 24584 8780 24636 8832
rect 25596 8823 25648 8832
rect 25596 8789 25605 8823
rect 25605 8789 25639 8823
rect 25639 8789 25648 8823
rect 25596 8780 25648 8789
rect 25964 8780 26016 8832
rect 4250 8678 4302 8730
rect 4314 8678 4366 8730
rect 4378 8678 4430 8730
rect 4442 8678 4494 8730
rect 4506 8678 4558 8730
rect 11955 8678 12007 8730
rect 12019 8678 12071 8730
rect 12083 8678 12135 8730
rect 12147 8678 12199 8730
rect 12211 8678 12263 8730
rect 19660 8678 19712 8730
rect 19724 8678 19776 8730
rect 19788 8678 19840 8730
rect 19852 8678 19904 8730
rect 19916 8678 19968 8730
rect 27365 8678 27417 8730
rect 27429 8678 27481 8730
rect 27493 8678 27545 8730
rect 27557 8678 27609 8730
rect 27621 8678 27673 8730
rect 6736 8415 6788 8424
rect 6736 8381 6745 8415
rect 6745 8381 6779 8415
rect 6779 8381 6788 8415
rect 6736 8372 6788 8381
rect 7656 8576 7708 8628
rect 8300 8576 8352 8628
rect 9036 8576 9088 8628
rect 10048 8576 10100 8628
rect 7196 8508 7248 8560
rect 7840 8508 7892 8560
rect 7656 8372 7708 8424
rect 7932 8304 7984 8356
rect 8484 8415 8536 8424
rect 8484 8381 8493 8415
rect 8493 8381 8527 8415
rect 8527 8381 8536 8415
rect 8484 8372 8536 8381
rect 8668 8508 8720 8560
rect 8668 8372 8720 8424
rect 8852 8551 8904 8560
rect 8852 8517 8861 8551
rect 8861 8517 8895 8551
rect 8895 8517 8904 8551
rect 8852 8508 8904 8517
rect 10692 8576 10744 8628
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 10416 8372 10468 8424
rect 10784 8508 10836 8560
rect 12624 8576 12676 8628
rect 15568 8576 15620 8628
rect 13176 8508 13228 8560
rect 14096 8551 14148 8560
rect 14096 8517 14105 8551
rect 14105 8517 14139 8551
rect 14139 8517 14148 8551
rect 14096 8508 14148 8517
rect 10600 8372 10652 8424
rect 11152 8372 11204 8424
rect 11336 8415 11388 8424
rect 11336 8381 11345 8415
rect 11345 8381 11379 8415
rect 11379 8381 11388 8415
rect 11336 8372 11388 8381
rect 11520 8372 11572 8424
rect 12900 8440 12952 8492
rect 11704 8372 11756 8424
rect 13268 8372 13320 8424
rect 13360 8372 13412 8424
rect 13820 8372 13872 8424
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 8944 8304 8996 8356
rect 9772 8304 9824 8356
rect 10140 8304 10192 8356
rect 7748 8236 7800 8288
rect 8116 8236 8168 8288
rect 10048 8236 10100 8288
rect 10600 8279 10652 8288
rect 10600 8245 10609 8279
rect 10609 8245 10643 8279
rect 10643 8245 10652 8279
rect 10600 8236 10652 8245
rect 11428 8347 11480 8356
rect 11428 8313 11437 8347
rect 11437 8313 11471 8347
rect 11471 8313 11480 8347
rect 11428 8304 11480 8313
rect 13084 8304 13136 8356
rect 13912 8304 13964 8356
rect 15292 8304 15344 8356
rect 16764 8576 16816 8628
rect 18236 8576 18288 8628
rect 18328 8576 18380 8628
rect 18788 8576 18840 8628
rect 16856 8372 16908 8424
rect 20352 8508 20404 8560
rect 17960 8415 18012 8424
rect 17960 8381 17969 8415
rect 17969 8381 18003 8415
rect 18003 8381 18012 8415
rect 18880 8440 18932 8492
rect 17960 8372 18012 8381
rect 17132 8304 17184 8356
rect 18512 8304 18564 8356
rect 12992 8279 13044 8288
rect 12992 8245 13001 8279
rect 13001 8245 13035 8279
rect 13035 8245 13044 8279
rect 12992 8236 13044 8245
rect 13728 8236 13780 8288
rect 17500 8279 17552 8288
rect 17500 8245 17509 8279
rect 17509 8245 17543 8279
rect 17543 8245 17552 8279
rect 17500 8236 17552 8245
rect 19432 8415 19484 8424
rect 19432 8381 19441 8415
rect 19441 8381 19475 8415
rect 19475 8381 19484 8415
rect 19432 8372 19484 8381
rect 20260 8415 20312 8424
rect 20260 8381 20269 8415
rect 20269 8381 20303 8415
rect 20303 8381 20312 8415
rect 20260 8372 20312 8381
rect 20536 8415 20588 8424
rect 20536 8381 20545 8415
rect 20545 8381 20579 8415
rect 20579 8381 20588 8415
rect 20536 8372 20588 8381
rect 21824 8576 21876 8628
rect 20904 8508 20956 8560
rect 22836 8551 22888 8560
rect 22836 8517 22845 8551
rect 22845 8517 22879 8551
rect 22879 8517 22888 8551
rect 22836 8508 22888 8517
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 21456 8440 21508 8449
rect 19156 8236 19208 8288
rect 19432 8236 19484 8288
rect 20260 8236 20312 8288
rect 21180 8415 21232 8424
rect 21180 8381 21189 8415
rect 21189 8381 21223 8415
rect 21223 8381 21232 8415
rect 21180 8372 21232 8381
rect 23020 8415 23072 8424
rect 23020 8381 23029 8415
rect 23029 8381 23063 8415
rect 23063 8381 23072 8415
rect 23020 8372 23072 8381
rect 24032 8576 24084 8628
rect 25228 8576 25280 8628
rect 25504 8576 25556 8628
rect 25688 8576 25740 8628
rect 23388 8551 23440 8560
rect 23388 8517 23397 8551
rect 23397 8517 23431 8551
rect 23431 8517 23440 8551
rect 23388 8508 23440 8517
rect 23480 8508 23532 8560
rect 24032 8372 24084 8424
rect 24124 8415 24176 8424
rect 24124 8381 24133 8415
rect 24133 8381 24167 8415
rect 24167 8381 24176 8415
rect 24124 8372 24176 8381
rect 21916 8304 21968 8356
rect 24584 8440 24636 8492
rect 26056 8508 26108 8560
rect 25228 8440 25280 8492
rect 25412 8415 25464 8424
rect 25412 8381 25421 8415
rect 25421 8381 25455 8415
rect 25455 8381 25464 8415
rect 25412 8372 25464 8381
rect 21180 8236 21232 8288
rect 24584 8304 24636 8356
rect 25872 8372 25924 8424
rect 26332 8415 26384 8424
rect 26332 8381 26341 8415
rect 26341 8381 26375 8415
rect 26375 8381 26384 8415
rect 26332 8372 26384 8381
rect 23020 8279 23072 8288
rect 23020 8245 23029 8279
rect 23029 8245 23063 8279
rect 23063 8245 23072 8279
rect 23020 8236 23072 8245
rect 24124 8236 24176 8288
rect 25044 8279 25096 8288
rect 25044 8245 25053 8279
rect 25053 8245 25087 8279
rect 25087 8245 25096 8279
rect 25044 8236 25096 8245
rect 25596 8279 25648 8288
rect 25596 8245 25605 8279
rect 25605 8245 25639 8279
rect 25639 8245 25648 8279
rect 25596 8236 25648 8245
rect 8102 8134 8154 8186
rect 8166 8134 8218 8186
rect 8230 8134 8282 8186
rect 8294 8134 8346 8186
rect 8358 8134 8410 8186
rect 15807 8134 15859 8186
rect 15871 8134 15923 8186
rect 15935 8134 15987 8186
rect 15999 8134 16051 8186
rect 16063 8134 16115 8186
rect 23512 8134 23564 8186
rect 23576 8134 23628 8186
rect 23640 8134 23692 8186
rect 23704 8134 23756 8186
rect 23768 8134 23820 8186
rect 31217 8134 31269 8186
rect 31281 8134 31333 8186
rect 31345 8134 31397 8186
rect 31409 8134 31461 8186
rect 31473 8134 31525 8186
rect 7656 8032 7708 8084
rect 7748 8032 7800 8084
rect 8484 8032 8536 8084
rect 8024 7939 8076 7948
rect 8024 7905 8033 7939
rect 8033 7905 8067 7939
rect 8067 7905 8076 7939
rect 8024 7896 8076 7905
rect 8300 7939 8352 7948
rect 8300 7905 8309 7939
rect 8309 7905 8343 7939
rect 8343 7905 8352 7939
rect 8300 7896 8352 7905
rect 8484 7896 8536 7948
rect 8760 8032 8812 8084
rect 9588 8032 9640 8084
rect 9680 8032 9732 8084
rect 9864 8032 9916 8084
rect 10600 8032 10652 8084
rect 10692 8032 10744 8084
rect 8576 7828 8628 7880
rect 7196 7692 7248 7744
rect 7656 7735 7708 7744
rect 7656 7701 7665 7735
rect 7665 7701 7699 7735
rect 7699 7701 7708 7735
rect 7656 7692 7708 7701
rect 8116 7760 8168 7812
rect 8852 7760 8904 7812
rect 10232 7939 10284 7948
rect 10232 7905 10241 7939
rect 10241 7905 10275 7939
rect 10275 7905 10284 7939
rect 10232 7896 10284 7905
rect 10324 7939 10376 7948
rect 10324 7905 10333 7939
rect 10333 7905 10367 7939
rect 10367 7905 10376 7939
rect 10324 7896 10376 7905
rect 11520 7964 11572 8016
rect 17592 8032 17644 8084
rect 12900 7964 12952 8016
rect 13728 7964 13780 8016
rect 10784 7896 10836 7948
rect 10048 7828 10100 7880
rect 9496 7760 9548 7812
rect 11152 7760 11204 7812
rect 11704 7760 11756 7812
rect 9128 7692 9180 7744
rect 9588 7735 9640 7744
rect 9588 7701 9597 7735
rect 9597 7701 9631 7735
rect 9631 7701 9640 7735
rect 9588 7692 9640 7701
rect 9864 7735 9916 7744
rect 9864 7701 9873 7735
rect 9873 7701 9907 7735
rect 9907 7701 9916 7735
rect 9864 7692 9916 7701
rect 12624 7692 12676 7744
rect 13268 7939 13320 7948
rect 13268 7905 13277 7939
rect 13277 7905 13311 7939
rect 13311 7905 13320 7939
rect 13268 7896 13320 7905
rect 14832 7896 14884 7948
rect 15292 8007 15344 8016
rect 15292 7973 15301 8007
rect 15301 7973 15335 8007
rect 15335 7973 15344 8007
rect 15292 7964 15344 7973
rect 15568 7760 15620 7812
rect 13176 7692 13228 7744
rect 14280 7692 14332 7744
rect 14372 7692 14424 7744
rect 18788 7964 18840 8016
rect 19340 7964 19392 8016
rect 23020 8032 23072 8084
rect 21456 7964 21508 8016
rect 21916 7964 21968 8016
rect 16212 7939 16264 7948
rect 16212 7905 16221 7939
rect 16221 7905 16255 7939
rect 16255 7905 16264 7939
rect 16212 7896 16264 7905
rect 16856 7896 16908 7948
rect 18512 7896 18564 7948
rect 20260 7828 20312 7880
rect 21732 7896 21784 7948
rect 22928 7896 22980 7948
rect 22100 7828 22152 7880
rect 25596 8032 25648 8084
rect 25504 7964 25556 8016
rect 15844 7735 15896 7744
rect 15844 7701 15853 7735
rect 15853 7701 15887 7735
rect 15887 7701 15896 7735
rect 15844 7692 15896 7701
rect 16304 7735 16356 7744
rect 16304 7701 16313 7735
rect 16313 7701 16347 7735
rect 16347 7701 16356 7735
rect 16304 7692 16356 7701
rect 16488 7692 16540 7744
rect 16672 7692 16724 7744
rect 19064 7760 19116 7812
rect 19524 7760 19576 7812
rect 25136 7896 25188 7948
rect 25228 7939 25280 7948
rect 25228 7905 25237 7939
rect 25237 7905 25271 7939
rect 25271 7905 25280 7939
rect 25228 7896 25280 7905
rect 25412 7896 25464 7948
rect 24768 7871 24820 7880
rect 24768 7837 24777 7871
rect 24777 7837 24811 7871
rect 24811 7837 24820 7871
rect 24768 7828 24820 7837
rect 25596 7828 25648 7880
rect 17960 7692 18012 7744
rect 18144 7735 18196 7744
rect 18144 7701 18153 7735
rect 18153 7701 18187 7735
rect 18187 7701 18196 7735
rect 18144 7692 18196 7701
rect 19984 7692 20036 7744
rect 21732 7692 21784 7744
rect 25504 7760 25556 7812
rect 24860 7692 24912 7744
rect 25688 7692 25740 7744
rect 25780 7692 25832 7744
rect 25872 7735 25924 7744
rect 25872 7701 25881 7735
rect 25881 7701 25915 7735
rect 25915 7701 25924 7735
rect 25872 7692 25924 7701
rect 26148 7735 26200 7744
rect 26148 7701 26157 7735
rect 26157 7701 26191 7735
rect 26191 7701 26200 7735
rect 26148 7692 26200 7701
rect 4250 7590 4302 7642
rect 4314 7590 4366 7642
rect 4378 7590 4430 7642
rect 4442 7590 4494 7642
rect 4506 7590 4558 7642
rect 11955 7590 12007 7642
rect 12019 7590 12071 7642
rect 12083 7590 12135 7642
rect 12147 7590 12199 7642
rect 12211 7590 12263 7642
rect 19660 7590 19712 7642
rect 19724 7590 19776 7642
rect 19788 7590 19840 7642
rect 19852 7590 19904 7642
rect 19916 7590 19968 7642
rect 27365 7590 27417 7642
rect 27429 7590 27481 7642
rect 27493 7590 27545 7642
rect 27557 7590 27609 7642
rect 27621 7590 27673 7642
rect 7012 7531 7064 7540
rect 7012 7497 7021 7531
rect 7021 7497 7055 7531
rect 7055 7497 7064 7531
rect 7012 7488 7064 7497
rect 7564 7488 7616 7540
rect 7840 7488 7892 7540
rect 8116 7488 8168 7540
rect 8300 7488 8352 7540
rect 9588 7488 9640 7540
rect 11336 7488 11388 7540
rect 9220 7420 9272 7472
rect 7012 7284 7064 7336
rect 7104 7327 7156 7336
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 7104 7284 7156 7293
rect 7288 7284 7340 7336
rect 7656 7327 7708 7336
rect 7656 7293 7657 7327
rect 7657 7293 7691 7327
rect 7691 7293 7708 7327
rect 7656 7284 7708 7293
rect 8760 7352 8812 7404
rect 6920 7148 6972 7200
rect 7104 7148 7156 7200
rect 7656 7148 7708 7200
rect 8116 7284 8168 7336
rect 8484 7216 8536 7268
rect 8944 7329 8996 7336
rect 8944 7295 8953 7329
rect 8953 7295 8987 7329
rect 8987 7295 8996 7329
rect 8944 7284 8996 7295
rect 9128 7352 9180 7404
rect 9588 7352 9640 7404
rect 9864 7352 9916 7404
rect 15292 7488 15344 7540
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 9496 7284 9548 7336
rect 9772 7327 9824 7336
rect 9772 7293 9781 7327
rect 9781 7293 9815 7327
rect 9815 7293 9824 7327
rect 9772 7284 9824 7293
rect 10140 7284 10192 7336
rect 14464 7420 14516 7472
rect 15844 7488 15896 7540
rect 16856 7488 16908 7540
rect 11244 7352 11296 7404
rect 11704 7352 11756 7404
rect 9864 7216 9916 7268
rect 10416 7216 10468 7268
rect 12532 7284 12584 7336
rect 12624 7284 12676 7336
rect 13268 7284 13320 7336
rect 13636 7284 13688 7336
rect 13728 7327 13780 7336
rect 13728 7293 13737 7327
rect 13737 7293 13771 7327
rect 13771 7293 13780 7327
rect 13728 7284 13780 7293
rect 13912 7284 13964 7336
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 12716 7216 12768 7268
rect 14648 7216 14700 7268
rect 15384 7216 15436 7268
rect 9220 7148 9272 7200
rect 10508 7148 10560 7200
rect 10876 7148 10928 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 11336 7148 11388 7200
rect 11520 7191 11572 7200
rect 11520 7157 11529 7191
rect 11529 7157 11563 7191
rect 11563 7157 11572 7191
rect 11520 7148 11572 7157
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 14096 7191 14148 7200
rect 14096 7157 14105 7191
rect 14105 7157 14139 7191
rect 14139 7157 14148 7191
rect 14096 7148 14148 7157
rect 14832 7148 14884 7200
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 15200 7191 15252 7200
rect 15200 7157 15209 7191
rect 15209 7157 15243 7191
rect 15243 7157 15252 7191
rect 15200 7148 15252 7157
rect 15568 7327 15620 7336
rect 15568 7293 15577 7327
rect 15577 7293 15611 7327
rect 15611 7293 15620 7327
rect 15568 7284 15620 7293
rect 16488 7420 16540 7472
rect 16304 7352 16356 7404
rect 16764 7352 16816 7404
rect 16672 7327 16724 7336
rect 16672 7293 16673 7327
rect 16673 7293 16707 7327
rect 16707 7293 16724 7327
rect 17776 7488 17828 7540
rect 18788 7488 18840 7540
rect 18604 7420 18656 7472
rect 19432 7420 19484 7472
rect 19800 7420 19852 7472
rect 15660 7216 15712 7268
rect 16672 7284 16724 7293
rect 17132 7284 17184 7336
rect 18696 7327 18748 7336
rect 18696 7293 18705 7327
rect 18705 7293 18739 7327
rect 18739 7293 18748 7327
rect 18696 7284 18748 7293
rect 18880 7284 18932 7336
rect 19064 7284 19116 7336
rect 19616 7395 19668 7404
rect 19616 7361 19625 7395
rect 19625 7361 19659 7395
rect 19659 7361 19668 7395
rect 19616 7352 19668 7361
rect 23388 7420 23440 7472
rect 20168 7284 20220 7336
rect 21916 7395 21968 7404
rect 21916 7361 21925 7395
rect 21925 7361 21959 7395
rect 21959 7361 21968 7395
rect 21916 7352 21968 7361
rect 23756 7420 23808 7472
rect 24492 7531 24544 7540
rect 24492 7497 24501 7531
rect 24501 7497 24535 7531
rect 24535 7497 24544 7531
rect 24492 7488 24544 7497
rect 24584 7488 24636 7540
rect 25596 7531 25648 7540
rect 25596 7497 25605 7531
rect 25605 7497 25639 7531
rect 25639 7497 25648 7531
rect 25596 7488 25648 7497
rect 25780 7488 25832 7540
rect 23940 7352 23992 7404
rect 18972 7216 19024 7268
rect 21364 7216 21416 7268
rect 24124 7284 24176 7336
rect 24216 7284 24268 7336
rect 24492 7284 24544 7336
rect 25228 7420 25280 7472
rect 24952 7327 25004 7336
rect 24952 7293 24961 7327
rect 24961 7293 24995 7327
rect 24995 7293 25004 7327
rect 24952 7284 25004 7293
rect 25044 7284 25096 7336
rect 25412 7327 25464 7336
rect 18328 7148 18380 7200
rect 18420 7191 18472 7200
rect 18420 7157 18429 7191
rect 18429 7157 18463 7191
rect 18463 7157 18472 7191
rect 18420 7148 18472 7157
rect 18512 7148 18564 7200
rect 19156 7148 19208 7200
rect 19800 7148 19852 7200
rect 19892 7191 19944 7200
rect 19892 7157 19901 7191
rect 19901 7157 19935 7191
rect 19935 7157 19944 7191
rect 19892 7148 19944 7157
rect 20168 7191 20220 7200
rect 20168 7157 20177 7191
rect 20177 7157 20211 7191
rect 20211 7157 20220 7191
rect 20168 7148 20220 7157
rect 20352 7148 20404 7200
rect 20996 7191 21048 7200
rect 20996 7157 21005 7191
rect 21005 7157 21039 7191
rect 21039 7157 21048 7191
rect 20996 7148 21048 7157
rect 21548 7191 21600 7200
rect 21548 7157 21557 7191
rect 21557 7157 21591 7191
rect 21591 7157 21600 7191
rect 21548 7148 21600 7157
rect 23112 7148 23164 7200
rect 23204 7148 23256 7200
rect 24124 7148 24176 7200
rect 25044 7148 25096 7200
rect 25412 7293 25421 7327
rect 25421 7293 25455 7327
rect 25455 7293 25464 7327
rect 25412 7284 25464 7293
rect 25504 7327 25556 7336
rect 25504 7293 25513 7327
rect 25513 7293 25547 7327
rect 25547 7293 25556 7327
rect 25504 7284 25556 7293
rect 25320 7191 25372 7200
rect 25320 7157 25329 7191
rect 25329 7157 25363 7191
rect 25363 7157 25372 7191
rect 25320 7148 25372 7157
rect 8102 7046 8154 7098
rect 8166 7046 8218 7098
rect 8230 7046 8282 7098
rect 8294 7046 8346 7098
rect 8358 7046 8410 7098
rect 15807 7046 15859 7098
rect 15871 7046 15923 7098
rect 15935 7046 15987 7098
rect 15999 7046 16051 7098
rect 16063 7046 16115 7098
rect 23512 7046 23564 7098
rect 23576 7046 23628 7098
rect 23640 7046 23692 7098
rect 23704 7046 23756 7098
rect 23768 7046 23820 7098
rect 31217 7046 31269 7098
rect 31281 7046 31333 7098
rect 31345 7046 31397 7098
rect 31409 7046 31461 7098
rect 31473 7046 31525 7098
rect 6920 6944 6972 6996
rect 7012 6944 7064 6996
rect 8024 6944 8076 6996
rect 8484 6944 8536 6996
rect 9680 6944 9732 6996
rect 9772 6944 9824 6996
rect 10508 6944 10560 6996
rect 11060 6944 11112 6996
rect 14556 6944 14608 6996
rect 15384 6944 15436 6996
rect 6552 6851 6604 6860
rect 6552 6817 6570 6851
rect 6570 6817 6604 6851
rect 6552 6808 6604 6817
rect 6828 6851 6880 6860
rect 6828 6817 6846 6851
rect 6846 6817 6880 6851
rect 6828 6808 6880 6817
rect 7196 6876 7248 6928
rect 7472 6851 7524 6860
rect 7472 6817 7480 6851
rect 7480 6817 7524 6851
rect 7472 6808 7524 6817
rect 7932 6808 7984 6860
rect 8208 6808 8260 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 8668 6876 8720 6928
rect 8760 6876 8812 6928
rect 8852 6851 8904 6860
rect 8852 6817 8861 6851
rect 8861 6817 8895 6851
rect 8895 6817 8904 6851
rect 8852 6808 8904 6817
rect 9220 6808 9272 6860
rect 11336 6876 11388 6928
rect 11704 6919 11756 6928
rect 11704 6885 11713 6919
rect 11713 6885 11747 6919
rect 11747 6885 11756 6919
rect 16764 6944 16816 6996
rect 18420 6944 18472 6996
rect 18880 6944 18932 6996
rect 19892 6944 19944 6996
rect 20168 6944 20220 6996
rect 20996 6944 21048 6996
rect 21088 6944 21140 6996
rect 11704 6876 11756 6885
rect 7380 6672 7432 6724
rect 6460 6604 6512 6656
rect 6736 6604 6788 6656
rect 7012 6604 7064 6656
rect 7196 6604 7248 6656
rect 7288 6604 7340 6656
rect 8392 6740 8444 6792
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 10416 6808 10468 6860
rect 9588 6672 9640 6724
rect 9772 6715 9824 6724
rect 9772 6681 9781 6715
rect 9781 6681 9815 6715
rect 9815 6681 9824 6715
rect 9772 6672 9824 6681
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 11428 6851 11480 6860
rect 11428 6817 11437 6851
rect 11437 6817 11471 6851
rect 11471 6817 11480 6851
rect 11428 6808 11480 6817
rect 16212 6876 16264 6928
rect 11152 6740 11204 6792
rect 12256 6808 12308 6860
rect 12532 6808 12584 6860
rect 14832 6808 14884 6860
rect 14924 6808 14976 6860
rect 10600 6672 10652 6724
rect 10692 6672 10744 6724
rect 11520 6672 11572 6724
rect 13636 6740 13688 6792
rect 12348 6672 12400 6724
rect 15476 6808 15528 6860
rect 17592 6876 17644 6928
rect 16764 6808 16816 6860
rect 18696 6808 18748 6860
rect 19708 6876 19760 6928
rect 23940 6944 23992 6996
rect 24584 6944 24636 6996
rect 25504 6944 25556 6996
rect 17868 6740 17920 6792
rect 18788 6740 18840 6792
rect 19340 6851 19392 6860
rect 19340 6817 19349 6851
rect 19349 6817 19383 6851
rect 19383 6817 19392 6851
rect 19340 6808 19392 6817
rect 20444 6851 20496 6860
rect 20444 6817 20453 6851
rect 20453 6817 20487 6851
rect 20487 6817 20496 6851
rect 20444 6808 20496 6817
rect 12256 6604 12308 6656
rect 13176 6604 13228 6656
rect 13728 6604 13780 6656
rect 15568 6647 15620 6656
rect 15568 6613 15577 6647
rect 15577 6613 15611 6647
rect 15611 6613 15620 6647
rect 15568 6604 15620 6613
rect 17960 6604 18012 6656
rect 19616 6672 19668 6724
rect 20536 6740 20588 6792
rect 21272 6851 21324 6860
rect 21272 6817 21281 6851
rect 21281 6817 21315 6851
rect 21315 6817 21324 6851
rect 21272 6808 21324 6817
rect 21824 6808 21876 6860
rect 21916 6808 21968 6860
rect 24032 6876 24084 6928
rect 22376 6740 22428 6792
rect 23572 6851 23624 6860
rect 23572 6817 23581 6851
rect 23581 6817 23615 6851
rect 23615 6817 23624 6851
rect 23572 6808 23624 6817
rect 23664 6851 23716 6860
rect 23664 6817 23673 6851
rect 23673 6817 23707 6851
rect 23707 6817 23716 6851
rect 23664 6808 23716 6817
rect 23296 6740 23348 6792
rect 24216 6851 24268 6860
rect 24216 6817 24225 6851
rect 24225 6817 24259 6851
rect 24259 6817 24268 6851
rect 24216 6808 24268 6817
rect 24400 6808 24452 6860
rect 24492 6851 24544 6860
rect 24492 6817 24501 6851
rect 24501 6817 24535 6851
rect 24535 6817 24544 6851
rect 24492 6808 24544 6817
rect 25228 6876 25280 6928
rect 24124 6740 24176 6792
rect 24952 6672 25004 6724
rect 18696 6604 18748 6656
rect 19524 6604 19576 6656
rect 20720 6604 20772 6656
rect 20904 6604 20956 6656
rect 21180 6604 21232 6656
rect 22192 6604 22244 6656
rect 22652 6647 22704 6656
rect 22652 6613 22661 6647
rect 22661 6613 22695 6647
rect 22695 6613 22704 6647
rect 22652 6604 22704 6613
rect 22744 6604 22796 6656
rect 23112 6604 23164 6656
rect 23480 6647 23532 6656
rect 23480 6613 23489 6647
rect 23489 6613 23523 6647
rect 23523 6613 23532 6647
rect 23480 6604 23532 6613
rect 23756 6647 23808 6656
rect 23756 6613 23765 6647
rect 23765 6613 23799 6647
rect 23799 6613 23808 6647
rect 23756 6604 23808 6613
rect 24308 6604 24360 6656
rect 24584 6647 24636 6656
rect 24584 6613 24593 6647
rect 24593 6613 24627 6647
rect 24627 6613 24636 6647
rect 24584 6604 24636 6613
rect 4250 6502 4302 6554
rect 4314 6502 4366 6554
rect 4378 6502 4430 6554
rect 4442 6502 4494 6554
rect 4506 6502 4558 6554
rect 11955 6502 12007 6554
rect 12019 6502 12071 6554
rect 12083 6502 12135 6554
rect 12147 6502 12199 6554
rect 12211 6502 12263 6554
rect 19660 6502 19712 6554
rect 19724 6502 19776 6554
rect 19788 6502 19840 6554
rect 19852 6502 19904 6554
rect 19916 6502 19968 6554
rect 27365 6502 27417 6554
rect 27429 6502 27481 6554
rect 27493 6502 27545 6554
rect 27557 6502 27609 6554
rect 27621 6502 27673 6554
rect 6460 6400 6512 6452
rect 7288 6400 7340 6452
rect 7472 6400 7524 6452
rect 8208 6400 8260 6452
rect 10140 6400 10192 6452
rect 10232 6400 10284 6452
rect 10600 6400 10652 6452
rect 11244 6400 11296 6452
rect 9496 6332 9548 6384
rect 9680 6375 9732 6384
rect 9680 6341 9689 6375
rect 9689 6341 9723 6375
rect 9723 6341 9732 6375
rect 9680 6332 9732 6341
rect 9864 6332 9916 6384
rect 10140 6307 10192 6316
rect 7104 6196 7156 6248
rect 7196 6196 7248 6248
rect 7840 6239 7892 6248
rect 7840 6205 7874 6239
rect 7874 6205 7892 6239
rect 7840 6196 7892 6205
rect 8024 6196 8076 6248
rect 8576 6128 8628 6180
rect 8944 6171 8996 6180
rect 8944 6137 8953 6171
rect 8953 6137 8987 6171
rect 8987 6137 8996 6171
rect 8944 6128 8996 6137
rect 9036 6128 9088 6180
rect 9312 6196 9364 6248
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 12716 6443 12768 6452
rect 12716 6409 12725 6443
rect 12725 6409 12759 6443
rect 12759 6409 12768 6443
rect 12716 6400 12768 6409
rect 15292 6332 15344 6384
rect 10692 6264 10744 6316
rect 11060 6307 11112 6316
rect 11060 6273 11069 6307
rect 11069 6273 11103 6307
rect 11103 6273 11112 6307
rect 11060 6264 11112 6273
rect 7380 6060 7432 6112
rect 8760 6103 8812 6112
rect 8760 6069 8769 6103
rect 8769 6069 8803 6103
rect 8803 6069 8812 6103
rect 8760 6060 8812 6069
rect 9220 6060 9272 6112
rect 10784 6239 10836 6248
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 11152 6196 11204 6248
rect 13912 6264 13964 6316
rect 11796 6128 11848 6180
rect 13176 6239 13228 6248
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 13820 6239 13872 6248
rect 13820 6205 13829 6239
rect 13829 6205 13863 6239
rect 13863 6205 13872 6239
rect 13820 6196 13872 6205
rect 15200 6196 15252 6248
rect 16764 6400 16816 6452
rect 18604 6400 18656 6452
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 19340 6400 19392 6452
rect 19524 6400 19576 6452
rect 20260 6400 20312 6452
rect 21732 6443 21784 6452
rect 21732 6409 21741 6443
rect 21741 6409 21775 6443
rect 21775 6409 21784 6443
rect 21732 6400 21784 6409
rect 21824 6400 21876 6452
rect 21916 6400 21968 6452
rect 23664 6400 23716 6452
rect 24492 6400 24544 6452
rect 18052 6332 18104 6384
rect 18328 6375 18380 6384
rect 18328 6341 18337 6375
rect 18337 6341 18371 6375
rect 18371 6341 18380 6375
rect 18328 6332 18380 6341
rect 19156 6332 19208 6384
rect 17960 6264 18012 6316
rect 10600 6060 10652 6112
rect 12256 6060 12308 6112
rect 12624 6060 12676 6112
rect 16856 6196 16908 6248
rect 18696 6264 18748 6316
rect 18328 6196 18380 6248
rect 13636 6060 13688 6112
rect 15200 6060 15252 6112
rect 15660 6060 15712 6112
rect 18880 6239 18932 6248
rect 18880 6205 18889 6239
rect 18889 6205 18923 6239
rect 18923 6205 18932 6239
rect 18880 6196 18932 6205
rect 19156 6196 19208 6248
rect 20812 6332 20864 6384
rect 21272 6264 21324 6316
rect 20904 6196 20956 6248
rect 20076 6128 20128 6180
rect 20352 6128 20404 6180
rect 19248 6060 19300 6112
rect 21272 6128 21324 6180
rect 21732 6196 21784 6248
rect 22008 6196 22060 6248
rect 22100 6239 22152 6248
rect 22100 6205 22109 6239
rect 22109 6205 22143 6239
rect 22143 6205 22152 6239
rect 22100 6196 22152 6205
rect 22192 6239 22244 6248
rect 22192 6205 22201 6239
rect 22201 6205 22235 6239
rect 22235 6205 22244 6239
rect 22192 6196 22244 6205
rect 22284 6196 22336 6248
rect 23756 6264 23808 6316
rect 21456 6103 21508 6112
rect 21456 6069 21465 6103
rect 21465 6069 21499 6103
rect 21499 6069 21508 6103
rect 21456 6060 21508 6069
rect 23204 6239 23256 6248
rect 23204 6205 23213 6239
rect 23213 6205 23247 6239
rect 23247 6205 23256 6239
rect 23204 6196 23256 6205
rect 22928 6128 22980 6180
rect 23020 6128 23072 6180
rect 23388 6196 23440 6248
rect 25320 6196 25372 6248
rect 23848 6128 23900 6180
rect 22284 6103 22336 6112
rect 22284 6069 22293 6103
rect 22293 6069 22327 6103
rect 22327 6069 22336 6103
rect 22284 6060 22336 6069
rect 22836 6060 22888 6112
rect 23296 6103 23348 6112
rect 23296 6069 23305 6103
rect 23305 6069 23339 6103
rect 23339 6069 23348 6103
rect 23296 6060 23348 6069
rect 8102 5958 8154 6010
rect 8166 5958 8218 6010
rect 8230 5958 8282 6010
rect 8294 5958 8346 6010
rect 8358 5958 8410 6010
rect 15807 5958 15859 6010
rect 15871 5958 15923 6010
rect 15935 5958 15987 6010
rect 15999 5958 16051 6010
rect 16063 5958 16115 6010
rect 23512 5958 23564 6010
rect 23576 5958 23628 6010
rect 23640 5958 23692 6010
rect 23704 5958 23756 6010
rect 23768 5958 23820 6010
rect 31217 5958 31269 6010
rect 31281 5958 31333 6010
rect 31345 5958 31397 6010
rect 31409 5958 31461 6010
rect 31473 5958 31525 6010
rect 6736 5856 6788 5908
rect 7012 5856 7064 5908
rect 7840 5856 7892 5908
rect 8484 5856 8536 5908
rect 8944 5856 8996 5908
rect 9220 5856 9272 5908
rect 9496 5856 9548 5908
rect 8576 5720 8628 5772
rect 9036 5720 9088 5772
rect 6552 5652 6604 5704
rect 6828 5652 6880 5704
rect 8668 5652 8720 5704
rect 10048 5856 10100 5908
rect 12348 5856 12400 5908
rect 13820 5856 13872 5908
rect 14464 5856 14516 5908
rect 9680 5763 9732 5772
rect 9680 5729 9714 5763
rect 9714 5729 9732 5763
rect 9680 5720 9732 5729
rect 11336 5720 11388 5772
rect 13636 5788 13688 5840
rect 17868 5856 17920 5908
rect 18788 5856 18840 5908
rect 20444 5856 20496 5908
rect 20536 5856 20588 5908
rect 21916 5856 21968 5908
rect 22560 5856 22612 5908
rect 23296 5856 23348 5908
rect 24124 5856 24176 5908
rect 13544 5720 13596 5772
rect 10876 5652 10928 5704
rect 11428 5652 11480 5704
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 15016 5720 15068 5772
rect 15660 5720 15712 5772
rect 10968 5584 11020 5636
rect 9680 5516 9732 5568
rect 19156 5720 19208 5772
rect 19340 5720 19392 5772
rect 20076 5652 20128 5704
rect 20352 5720 20404 5772
rect 20720 5788 20772 5840
rect 21364 5831 21416 5840
rect 21364 5797 21373 5831
rect 21373 5797 21407 5831
rect 21407 5797 21416 5831
rect 21364 5788 21416 5797
rect 19064 5627 19116 5636
rect 19064 5593 19073 5627
rect 19073 5593 19107 5627
rect 19107 5593 19116 5627
rect 19064 5584 19116 5593
rect 19248 5584 19300 5636
rect 20812 5763 20864 5772
rect 20812 5729 20821 5763
rect 20821 5729 20855 5763
rect 20855 5729 20864 5763
rect 20812 5720 20864 5729
rect 20904 5720 20956 5772
rect 21456 5763 21508 5772
rect 21456 5729 21465 5763
rect 21465 5729 21499 5763
rect 21499 5729 21508 5763
rect 21456 5720 21508 5729
rect 21640 5763 21692 5772
rect 21640 5729 21649 5763
rect 21649 5729 21683 5763
rect 21683 5729 21692 5763
rect 21640 5720 21692 5729
rect 21824 5720 21876 5772
rect 21916 5720 21968 5772
rect 20720 5652 20772 5704
rect 21364 5652 21416 5704
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 21548 5584 21600 5636
rect 22376 5584 22428 5636
rect 26148 5720 26200 5772
rect 25872 5652 25924 5704
rect 22928 5584 22980 5636
rect 24216 5584 24268 5636
rect 16304 5516 16356 5568
rect 17316 5516 17368 5568
rect 20536 5516 20588 5568
rect 21916 5559 21968 5568
rect 21916 5525 21925 5559
rect 21925 5525 21959 5559
rect 21959 5525 21968 5559
rect 21916 5516 21968 5525
rect 24860 5516 24912 5568
rect 4250 5414 4302 5466
rect 4314 5414 4366 5466
rect 4378 5414 4430 5466
rect 4442 5414 4494 5466
rect 4506 5414 4558 5466
rect 11955 5414 12007 5466
rect 12019 5414 12071 5466
rect 12083 5414 12135 5466
rect 12147 5414 12199 5466
rect 12211 5414 12263 5466
rect 19660 5414 19712 5466
rect 19724 5414 19776 5466
rect 19788 5414 19840 5466
rect 19852 5414 19904 5466
rect 19916 5414 19968 5466
rect 27365 5414 27417 5466
rect 27429 5414 27481 5466
rect 27493 5414 27545 5466
rect 27557 5414 27609 5466
rect 27621 5414 27673 5466
rect 9588 5312 9640 5364
rect 9680 5312 9732 5364
rect 8392 5151 8444 5160
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 9404 5176 9456 5228
rect 11060 5312 11112 5364
rect 12532 5355 12584 5364
rect 12532 5321 12541 5355
rect 12541 5321 12575 5355
rect 12575 5321 12584 5355
rect 12532 5312 12584 5321
rect 13084 5355 13136 5364
rect 13084 5321 13093 5355
rect 13093 5321 13127 5355
rect 13127 5321 13136 5355
rect 13084 5312 13136 5321
rect 14556 5312 14608 5364
rect 15476 5312 15528 5364
rect 19248 5355 19300 5364
rect 19248 5321 19257 5355
rect 19257 5321 19291 5355
rect 19291 5321 19300 5355
rect 19248 5312 19300 5321
rect 19340 5312 19392 5364
rect 20536 5312 20588 5364
rect 16028 5244 16080 5296
rect 20812 5312 20864 5364
rect 21456 5355 21508 5364
rect 21456 5321 21465 5355
rect 21465 5321 21499 5355
rect 21499 5321 21508 5355
rect 21456 5312 21508 5321
rect 22008 5312 22060 5364
rect 24584 5312 24636 5364
rect 9772 5015 9824 5024
rect 9772 4981 9781 5015
rect 9781 4981 9815 5015
rect 9815 4981 9824 5015
rect 9772 4972 9824 4981
rect 10048 5108 10100 5160
rect 10416 5040 10468 5092
rect 11520 5108 11572 5160
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 10876 5040 10928 5092
rect 10140 5015 10192 5024
rect 10140 4981 10149 5015
rect 10149 4981 10183 5015
rect 10183 4981 10192 5015
rect 10140 4972 10192 4981
rect 11612 4972 11664 5024
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 13912 5151 13964 5160
rect 13912 5117 13921 5151
rect 13921 5117 13955 5151
rect 13955 5117 13964 5151
rect 13912 5108 13964 5117
rect 14464 5151 14516 5160
rect 14464 5117 14473 5151
rect 14473 5117 14507 5151
rect 14507 5117 14516 5151
rect 14464 5108 14516 5117
rect 15476 5176 15528 5228
rect 14924 5151 14976 5160
rect 14924 5117 14933 5151
rect 14933 5117 14967 5151
rect 14967 5117 14976 5151
rect 14924 5108 14976 5117
rect 15292 5108 15344 5160
rect 15384 5108 15436 5160
rect 16028 5108 16080 5160
rect 16856 5176 16908 5228
rect 17316 5151 17368 5160
rect 17316 5117 17350 5151
rect 17350 5117 17368 5151
rect 17316 5108 17368 5117
rect 19156 5151 19208 5160
rect 19156 5117 19157 5151
rect 19157 5117 19191 5151
rect 19191 5117 19208 5151
rect 14096 5040 14148 5092
rect 15108 5040 15160 5092
rect 16212 5040 16264 5092
rect 19156 5108 19208 5117
rect 19708 5108 19760 5160
rect 20260 5176 20312 5228
rect 20904 5244 20956 5296
rect 19984 5151 20036 5160
rect 19984 5117 19993 5151
rect 19993 5117 20027 5151
rect 20027 5117 20036 5151
rect 19984 5108 20036 5117
rect 20628 5108 20680 5160
rect 21916 5244 21968 5296
rect 22100 5244 22152 5296
rect 25688 5244 25740 5296
rect 14556 4972 14608 5024
rect 15200 4972 15252 5024
rect 15384 4972 15436 5024
rect 16028 4972 16080 5024
rect 16396 4972 16448 5024
rect 16488 5015 16540 5024
rect 16488 4981 16497 5015
rect 16497 4981 16531 5015
rect 16531 4981 16540 5015
rect 16488 4972 16540 4981
rect 16672 5015 16724 5024
rect 16672 4981 16699 5015
rect 16699 4981 16724 5015
rect 16672 4972 16724 4981
rect 16764 4972 16816 5024
rect 19524 4972 19576 5024
rect 20076 5015 20128 5024
rect 20076 4981 20085 5015
rect 20085 4981 20119 5015
rect 20119 4981 20128 5015
rect 20076 4972 20128 4981
rect 20536 4972 20588 5024
rect 21088 5040 21140 5092
rect 21548 5151 21600 5160
rect 21548 5117 21557 5151
rect 21557 5117 21591 5151
rect 21591 5117 21600 5151
rect 21548 5108 21600 5117
rect 21916 5108 21968 5160
rect 22100 5151 22152 5160
rect 22100 5117 22109 5151
rect 22109 5117 22143 5151
rect 22143 5117 22152 5151
rect 22100 5108 22152 5117
rect 22928 5176 22980 5228
rect 23388 5176 23440 5228
rect 22744 4972 22796 5024
rect 8102 4870 8154 4922
rect 8166 4870 8218 4922
rect 8230 4870 8282 4922
rect 8294 4870 8346 4922
rect 8358 4870 8410 4922
rect 15807 4870 15859 4922
rect 15871 4870 15923 4922
rect 15935 4870 15987 4922
rect 15999 4870 16051 4922
rect 16063 4870 16115 4922
rect 23512 4870 23564 4922
rect 23576 4870 23628 4922
rect 23640 4870 23692 4922
rect 23704 4870 23756 4922
rect 23768 4870 23820 4922
rect 31217 4870 31269 4922
rect 31281 4870 31333 4922
rect 31345 4870 31397 4922
rect 31409 4870 31461 4922
rect 31473 4870 31525 4922
rect 9312 4768 9364 4820
rect 10140 4768 10192 4820
rect 10324 4768 10376 4820
rect 10876 4768 10928 4820
rect 11336 4768 11388 4820
rect 9772 4700 9824 4752
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 10048 4632 10100 4684
rect 10140 4675 10192 4684
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 10508 4632 10560 4684
rect 10600 4632 10652 4684
rect 10692 4632 10744 4684
rect 11520 4700 11572 4752
rect 8760 4564 8812 4616
rect 9312 4471 9364 4480
rect 9312 4437 9321 4471
rect 9321 4437 9355 4471
rect 9355 4437 9364 4471
rect 9312 4428 9364 4437
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 11428 4632 11480 4641
rect 11796 4811 11848 4820
rect 11796 4777 11805 4811
rect 11805 4777 11839 4811
rect 11839 4777 11848 4811
rect 11796 4768 11848 4777
rect 13084 4768 13136 4820
rect 13268 4768 13320 4820
rect 13544 4768 13596 4820
rect 14096 4768 14148 4820
rect 14648 4768 14700 4820
rect 16212 4768 16264 4820
rect 16488 4768 16540 4820
rect 16764 4768 16816 4820
rect 19892 4768 19944 4820
rect 20076 4768 20128 4820
rect 21180 4768 21232 4820
rect 21916 4768 21968 4820
rect 23848 4768 23900 4820
rect 12992 4632 13044 4684
rect 14188 4700 14240 4752
rect 14096 4675 14148 4684
rect 14096 4641 14105 4675
rect 14105 4641 14139 4675
rect 14139 4641 14148 4675
rect 14096 4632 14148 4641
rect 14280 4675 14332 4684
rect 14280 4641 14289 4675
rect 14289 4641 14323 4675
rect 14323 4641 14332 4675
rect 14280 4632 14332 4641
rect 13820 4564 13872 4616
rect 14832 4632 14884 4684
rect 15476 4632 15528 4684
rect 15844 4675 15896 4684
rect 15844 4641 15853 4675
rect 15853 4641 15887 4675
rect 15887 4641 15896 4675
rect 15844 4632 15896 4641
rect 15936 4675 15988 4684
rect 15936 4641 15945 4675
rect 15945 4641 15979 4675
rect 15979 4641 15988 4675
rect 15936 4632 15988 4641
rect 16672 4700 16724 4752
rect 16488 4675 16540 4684
rect 16488 4641 16497 4675
rect 16497 4641 16531 4675
rect 16531 4641 16540 4675
rect 16488 4632 16540 4641
rect 10600 4496 10652 4548
rect 11428 4496 11480 4548
rect 12716 4496 12768 4548
rect 15660 4496 15712 4548
rect 16856 4632 16908 4684
rect 20444 4675 20496 4684
rect 20444 4641 20453 4675
rect 20453 4641 20487 4675
rect 20487 4641 20496 4675
rect 20444 4632 20496 4641
rect 11796 4428 11848 4480
rect 14188 4428 14240 4480
rect 15844 4428 15896 4480
rect 16396 4428 16448 4480
rect 19340 4564 19392 4616
rect 20168 4564 20220 4616
rect 20996 4675 21048 4684
rect 20996 4641 21005 4675
rect 21005 4641 21039 4675
rect 21039 4641 21048 4675
rect 20996 4632 21048 4641
rect 22836 4564 22888 4616
rect 21364 4496 21416 4548
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 18328 4428 18380 4437
rect 4250 4326 4302 4378
rect 4314 4326 4366 4378
rect 4378 4326 4430 4378
rect 4442 4326 4494 4378
rect 4506 4326 4558 4378
rect 11955 4326 12007 4378
rect 12019 4326 12071 4378
rect 12083 4326 12135 4378
rect 12147 4326 12199 4378
rect 12211 4326 12263 4378
rect 19660 4326 19712 4378
rect 19724 4326 19776 4378
rect 19788 4326 19840 4378
rect 19852 4326 19904 4378
rect 19916 4326 19968 4378
rect 27365 4326 27417 4378
rect 27429 4326 27481 4378
rect 27493 4326 27545 4378
rect 27557 4326 27609 4378
rect 27621 4326 27673 4378
rect 9312 4224 9364 4276
rect 9496 4156 9548 4208
rect 9864 4156 9916 4208
rect 8484 4088 8536 4140
rect 11796 4224 11848 4276
rect 15292 4267 15344 4276
rect 15292 4233 15301 4267
rect 15301 4233 15335 4267
rect 15335 4233 15344 4267
rect 15292 4224 15344 4233
rect 15844 4224 15896 4276
rect 18328 4224 18380 4276
rect 21916 4224 21968 4276
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 19524 4156 19576 4208
rect 20628 4156 20680 4208
rect 10140 4020 10192 4072
rect 10508 4020 10560 4072
rect 11428 4020 11480 4072
rect 14924 4088 14976 4140
rect 14188 4063 14240 4072
rect 14188 4029 14222 4063
rect 14222 4029 14240 4063
rect 14188 4020 14240 4029
rect 16396 3952 16448 4004
rect 10232 3884 10284 3936
rect 10600 3884 10652 3936
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 17040 3927 17092 3936
rect 17040 3893 17049 3927
rect 17049 3893 17083 3927
rect 17083 3893 17092 3927
rect 17040 3884 17092 3893
rect 8102 3782 8154 3834
rect 8166 3782 8218 3834
rect 8230 3782 8282 3834
rect 8294 3782 8346 3834
rect 8358 3782 8410 3834
rect 15807 3782 15859 3834
rect 15871 3782 15923 3834
rect 15935 3782 15987 3834
rect 15999 3782 16051 3834
rect 16063 3782 16115 3834
rect 23512 3782 23564 3834
rect 23576 3782 23628 3834
rect 23640 3782 23692 3834
rect 23704 3782 23756 3834
rect 23768 3782 23820 3834
rect 31217 3782 31269 3834
rect 31281 3782 31333 3834
rect 31345 3782 31397 3834
rect 31409 3782 31461 3834
rect 31473 3782 31525 3834
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 10140 3680 10192 3732
rect 8760 3612 8812 3664
rect 10232 3655 10284 3664
rect 10232 3621 10241 3655
rect 10241 3621 10275 3655
rect 10275 3621 10284 3655
rect 10232 3612 10284 3621
rect 8484 3544 8536 3596
rect 9036 3544 9088 3596
rect 14280 3680 14332 3732
rect 16396 3680 16448 3732
rect 10508 3408 10560 3460
rect 12808 3544 12860 3596
rect 12992 3544 13044 3596
rect 14096 3612 14148 3664
rect 15384 3655 15436 3664
rect 15384 3621 15393 3655
rect 15393 3621 15427 3655
rect 15427 3621 15436 3655
rect 15384 3612 15436 3621
rect 16212 3612 16264 3664
rect 17040 3612 17092 3664
rect 15016 3587 15068 3596
rect 15016 3553 15033 3587
rect 15033 3553 15067 3587
rect 15067 3553 15068 3587
rect 15016 3544 15068 3553
rect 16120 3544 16172 3596
rect 16488 3544 16540 3596
rect 16856 3544 16908 3596
rect 15292 3408 15344 3460
rect 10324 3340 10376 3392
rect 16120 3340 16172 3392
rect 23204 3340 23256 3392
rect 4250 3238 4302 3290
rect 4314 3238 4366 3290
rect 4378 3238 4430 3290
rect 4442 3238 4494 3290
rect 4506 3238 4558 3290
rect 11955 3238 12007 3290
rect 12019 3238 12071 3290
rect 12083 3238 12135 3290
rect 12147 3238 12199 3290
rect 12211 3238 12263 3290
rect 19660 3238 19712 3290
rect 19724 3238 19776 3290
rect 19788 3238 19840 3290
rect 19852 3238 19904 3290
rect 19916 3238 19968 3290
rect 27365 3238 27417 3290
rect 27429 3238 27481 3290
rect 27493 3238 27545 3290
rect 27557 3238 27609 3290
rect 27621 3238 27673 3290
rect 9680 2796 9732 2848
rect 11704 2796 11756 2848
rect 8102 2694 8154 2746
rect 8166 2694 8218 2746
rect 8230 2694 8282 2746
rect 8294 2694 8346 2746
rect 8358 2694 8410 2746
rect 15807 2694 15859 2746
rect 15871 2694 15923 2746
rect 15935 2694 15987 2746
rect 15999 2694 16051 2746
rect 16063 2694 16115 2746
rect 23512 2694 23564 2746
rect 23576 2694 23628 2746
rect 23640 2694 23692 2746
rect 23704 2694 23756 2746
rect 23768 2694 23820 2746
rect 31217 2694 31269 2746
rect 31281 2694 31333 2746
rect 31345 2694 31397 2746
rect 31409 2694 31461 2746
rect 31473 2694 31525 2746
rect 4250 2150 4302 2202
rect 4314 2150 4366 2202
rect 4378 2150 4430 2202
rect 4442 2150 4494 2202
rect 4506 2150 4558 2202
rect 11955 2150 12007 2202
rect 12019 2150 12071 2202
rect 12083 2150 12135 2202
rect 12147 2150 12199 2202
rect 12211 2150 12263 2202
rect 19660 2150 19712 2202
rect 19724 2150 19776 2202
rect 19788 2150 19840 2202
rect 19852 2150 19904 2202
rect 19916 2150 19968 2202
rect 27365 2150 27417 2202
rect 27429 2150 27481 2202
rect 27493 2150 27545 2202
rect 27557 2150 27609 2202
rect 27621 2150 27673 2202
rect 8102 1606 8154 1658
rect 8166 1606 8218 1658
rect 8230 1606 8282 1658
rect 8294 1606 8346 1658
rect 8358 1606 8410 1658
rect 15807 1606 15859 1658
rect 15871 1606 15923 1658
rect 15935 1606 15987 1658
rect 15999 1606 16051 1658
rect 16063 1606 16115 1658
rect 23512 1606 23564 1658
rect 23576 1606 23628 1658
rect 23640 1606 23692 1658
rect 23704 1606 23756 1658
rect 23768 1606 23820 1658
rect 31217 1606 31269 1658
rect 31281 1606 31333 1658
rect 31345 1606 31397 1658
rect 31409 1606 31461 1658
rect 31473 1606 31525 1658
rect 4250 1062 4302 1114
rect 4314 1062 4366 1114
rect 4378 1062 4430 1114
rect 4442 1062 4494 1114
rect 4506 1062 4558 1114
rect 11955 1062 12007 1114
rect 12019 1062 12071 1114
rect 12083 1062 12135 1114
rect 12147 1062 12199 1114
rect 12211 1062 12263 1114
rect 19660 1062 19712 1114
rect 19724 1062 19776 1114
rect 19788 1062 19840 1114
rect 19852 1062 19904 1114
rect 19916 1062 19968 1114
rect 27365 1062 27417 1114
rect 27429 1062 27481 1114
rect 27493 1062 27545 1114
rect 27557 1062 27609 1114
rect 27621 1062 27673 1114
rect 8668 960 8720 1012
rect 7840 799 7892 808
rect 7840 765 7849 799
rect 7849 765 7883 799
rect 7883 765 7892 799
rect 7840 756 7892 765
rect 8102 518 8154 570
rect 8166 518 8218 570
rect 8230 518 8282 570
rect 8294 518 8346 570
rect 8358 518 8410 570
rect 15807 518 15859 570
rect 15871 518 15923 570
rect 15935 518 15987 570
rect 15999 518 16051 570
rect 16063 518 16115 570
rect 23512 518 23564 570
rect 23576 518 23628 570
rect 23640 518 23692 570
rect 23704 518 23756 570
rect 23768 518 23820 570
rect 31217 518 31269 570
rect 31281 518 31333 570
rect 31345 518 31397 570
rect 31409 518 31461 570
rect 31473 518 31525 570
rect 16028 416 16080 468
rect 16304 416 16356 468
<< metal2 >>
rect 8390 19600 8446 20000
rect 9034 19600 9090 20000
rect 9678 19600 9734 20000
rect 10322 19600 10378 20000
rect 10966 19600 11022 20000
rect 11610 19600 11666 20000
rect 12254 19600 12310 20000
rect 12898 19600 12954 20000
rect 13004 19638 13308 19666
rect 8404 19258 8432 19600
rect 8404 19230 8524 19258
rect 8102 19068 8410 19077
rect 8102 19066 8108 19068
rect 8164 19066 8188 19068
rect 8244 19066 8268 19068
rect 8324 19066 8348 19068
rect 8404 19066 8410 19068
rect 8164 19014 8166 19066
rect 8346 19014 8348 19066
rect 8102 19012 8108 19014
rect 8164 19012 8188 19014
rect 8244 19012 8268 19014
rect 8324 19012 8348 19014
rect 8404 19012 8410 19014
rect 8102 19003 8410 19012
rect 4250 18524 4558 18533
rect 4250 18522 4256 18524
rect 4312 18522 4336 18524
rect 4392 18522 4416 18524
rect 4472 18522 4496 18524
rect 4552 18522 4558 18524
rect 4312 18470 4314 18522
rect 4494 18470 4496 18522
rect 4250 18468 4256 18470
rect 4312 18468 4336 18470
rect 4392 18468 4416 18470
rect 4472 18468 4496 18470
rect 4552 18468 4558 18470
rect 4250 18459 4558 18468
rect 8102 17980 8410 17989
rect 8102 17978 8108 17980
rect 8164 17978 8188 17980
rect 8244 17978 8268 17980
rect 8324 17978 8348 17980
rect 8404 17978 8410 17980
rect 8164 17926 8166 17978
rect 8346 17926 8348 17978
rect 8102 17924 8108 17926
rect 8164 17924 8188 17926
rect 8244 17924 8268 17926
rect 8324 17924 8348 17926
rect 8404 17924 8410 17926
rect 8102 17915 8410 17924
rect 4250 17436 4558 17445
rect 4250 17434 4256 17436
rect 4312 17434 4336 17436
rect 4392 17434 4416 17436
rect 4472 17434 4496 17436
rect 4552 17434 4558 17436
rect 4312 17382 4314 17434
rect 4494 17382 4496 17434
rect 4250 17380 4256 17382
rect 4312 17380 4336 17382
rect 4392 17380 4416 17382
rect 4472 17380 4496 17382
rect 4552 17380 4558 17382
rect 4250 17371 4558 17380
rect 8102 16892 8410 16901
rect 8102 16890 8108 16892
rect 8164 16890 8188 16892
rect 8244 16890 8268 16892
rect 8324 16890 8348 16892
rect 8404 16890 8410 16892
rect 8164 16838 8166 16890
rect 8346 16838 8348 16890
rect 8102 16836 8108 16838
rect 8164 16836 8188 16838
rect 8244 16836 8268 16838
rect 8324 16836 8348 16838
rect 8404 16836 8410 16838
rect 8102 16827 8410 16836
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 4250 16348 4558 16357
rect 4250 16346 4256 16348
rect 4312 16346 4336 16348
rect 4392 16346 4416 16348
rect 4472 16346 4496 16348
rect 4552 16346 4558 16348
rect 4312 16294 4314 16346
rect 4494 16294 4496 16346
rect 4250 16292 4256 16294
rect 4312 16292 4336 16294
rect 4392 16292 4416 16294
rect 4472 16292 4496 16294
rect 4552 16292 4558 16294
rect 4250 16283 4558 16292
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7378 15328 7434 15337
rect 4250 15260 4558 15269
rect 7378 15263 7434 15272
rect 4250 15258 4256 15260
rect 4312 15258 4336 15260
rect 4392 15258 4416 15260
rect 4472 15258 4496 15260
rect 4552 15258 4558 15260
rect 4312 15206 4314 15258
rect 4494 15206 4496 15258
rect 4250 15204 4256 15206
rect 4312 15204 4336 15206
rect 4392 15204 4416 15206
rect 4472 15204 4496 15206
rect 4552 15204 4558 15206
rect 4250 15195 4558 15204
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 4250 14172 4558 14181
rect 4250 14170 4256 14172
rect 4312 14170 4336 14172
rect 4392 14170 4416 14172
rect 4472 14170 4496 14172
rect 4552 14170 4558 14172
rect 4312 14118 4314 14170
rect 4494 14118 4496 14170
rect 4250 14116 4256 14118
rect 4312 14116 4336 14118
rect 4392 14116 4416 14118
rect 4472 14116 4496 14118
rect 4552 14116 4558 14118
rect 4250 14107 4558 14116
rect 7116 13870 7144 14214
rect 7208 14006 7236 14758
rect 7196 14000 7248 14006
rect 7196 13942 7248 13948
rect 7392 13870 7420 15263
rect 7484 13938 7512 16186
rect 7838 16008 7894 16017
rect 7760 15966 7838 15994
rect 7564 14544 7616 14550
rect 7654 14512 7710 14521
rect 7616 14492 7654 14498
rect 7564 14486 7654 14492
rect 7576 14470 7654 14486
rect 7654 14447 7710 14456
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7668 13870 7696 14447
rect 7760 13954 7788 15966
rect 7838 15943 7894 15952
rect 7838 15192 7894 15201
rect 7838 15127 7894 15136
rect 7852 14618 7880 15127
rect 7944 14618 7972 16730
rect 8496 16153 8524 19230
rect 9048 17354 9076 19600
rect 9048 17326 9168 17354
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 8482 16144 8538 16153
rect 8482 16079 8538 16088
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8036 14482 8064 15846
rect 8102 15804 8410 15813
rect 8102 15802 8108 15804
rect 8164 15802 8188 15804
rect 8244 15802 8268 15804
rect 8324 15802 8348 15804
rect 8404 15802 8410 15804
rect 8164 15750 8166 15802
rect 8346 15750 8348 15802
rect 8102 15748 8108 15750
rect 8164 15748 8188 15750
rect 8244 15748 8268 15750
rect 8324 15748 8348 15750
rect 8404 15748 8410 15750
rect 8102 15739 8410 15748
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8312 14822 8340 15302
rect 8496 14958 8524 15438
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8102 14716 8410 14725
rect 8102 14714 8108 14716
rect 8164 14714 8188 14716
rect 8244 14714 8268 14716
rect 8324 14714 8348 14716
rect 8404 14714 8410 14716
rect 8164 14662 8166 14714
rect 8346 14662 8348 14714
rect 8102 14660 8108 14662
rect 8164 14660 8188 14662
rect 8244 14660 8268 14662
rect 8324 14660 8348 14662
rect 8404 14660 8410 14662
rect 8102 14651 8410 14660
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 7852 14074 7880 14418
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 7944 13954 7972 14010
rect 7760 13926 7972 13954
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 4250 13084 4558 13093
rect 4250 13082 4256 13084
rect 4312 13082 4336 13084
rect 4392 13082 4416 13084
rect 4472 13082 4496 13084
rect 4552 13082 4558 13084
rect 4312 13030 4314 13082
rect 4494 13030 4496 13082
rect 4250 13028 4256 13030
rect 4312 13028 4336 13030
rect 4392 13028 4416 13030
rect 4472 13028 4496 13030
rect 4552 13028 4558 13030
rect 4250 13019 4558 13028
rect 7392 12306 7420 13126
rect 7576 12986 7604 13738
rect 7944 13530 7972 13806
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7656 13456 7708 13462
rect 7654 13424 7656 13433
rect 7708 13424 7710 13433
rect 7654 13359 7710 13368
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 8036 13376 8064 14214
rect 8128 13938 8156 14418
rect 8496 14396 8524 14894
rect 8404 14368 8524 14396
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8312 13938 8340 14282
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8208 13864 8260 13870
rect 8404 13818 8432 14368
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8260 13812 8432 13818
rect 8208 13806 8432 13812
rect 8220 13790 8432 13806
rect 8102 13628 8410 13637
rect 8102 13626 8108 13628
rect 8164 13626 8188 13628
rect 8244 13626 8268 13628
rect 8324 13626 8348 13628
rect 8404 13626 8410 13628
rect 8164 13574 8166 13626
rect 8346 13574 8348 13626
rect 8102 13572 8108 13574
rect 8164 13572 8188 13574
rect 8244 13572 8268 13574
rect 8324 13572 8348 13574
rect 8404 13572 8410 13574
rect 8102 13563 8410 13572
rect 8496 13530 8524 14214
rect 8588 14074 8616 15370
rect 8680 15162 8708 17002
rect 8760 16720 8812 16726
rect 8760 16662 8812 16668
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8772 14958 8800 16662
rect 9140 15881 9168 17326
rect 9586 16280 9642 16289
rect 9586 16215 9642 16224
rect 9126 15872 9182 15881
rect 9126 15807 9182 15816
rect 9494 15600 9550 15609
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 9416 15544 9494 15552
rect 9600 15586 9628 16215
rect 9692 15745 9720 19600
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9784 16182 9812 17070
rect 10230 16688 10286 16697
rect 10152 16646 10230 16674
rect 10048 16584 10100 16590
rect 10046 16552 10048 16561
rect 10100 16552 10102 16561
rect 10046 16487 10102 16496
rect 10046 16416 10102 16425
rect 10046 16351 10102 16360
rect 9772 16176 9824 16182
rect 9772 16118 9824 16124
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9678 15736 9734 15745
rect 9784 15706 9812 15982
rect 9678 15671 9734 15680
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9600 15570 9720 15586
rect 9600 15564 9732 15570
rect 9600 15558 9680 15564
rect 9416 15524 9496 15544
rect 8760 14952 8812 14958
rect 8666 14920 8722 14929
rect 8760 14894 8812 14900
rect 8666 14855 8722 14864
rect 8680 14482 8708 14855
rect 8956 14618 8984 15506
rect 9310 15464 9366 15473
rect 9232 15422 9310 15450
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 9140 14482 9168 15302
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8944 14408 8996 14414
rect 9232 14362 9260 15422
rect 9310 15399 9366 15408
rect 9312 14952 9364 14958
rect 9310 14920 9312 14929
rect 9364 14920 9366 14929
rect 9310 14855 9366 14864
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 8944 14350 8996 14356
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8116 13388 8168 13394
rect 8036 13348 8116 13376
rect 7944 13297 7972 13330
rect 7930 13288 7986 13297
rect 8036 13258 8064 13348
rect 8116 13330 8168 13336
rect 7930 13223 7986 13232
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12986 7788 13126
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 8036 12434 8064 13194
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12782 8156 13126
rect 8404 12782 8432 13466
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8102 12540 8410 12549
rect 8102 12538 8108 12540
rect 8164 12538 8188 12540
rect 8244 12538 8268 12540
rect 8324 12538 8348 12540
rect 8404 12538 8410 12540
rect 8164 12486 8166 12538
rect 8346 12486 8348 12538
rect 8102 12484 8108 12486
rect 8164 12484 8188 12486
rect 8244 12484 8268 12486
rect 8324 12484 8348 12486
rect 8404 12484 8410 12486
rect 8102 12475 8410 12484
rect 8496 12442 8524 12582
rect 8588 12442 8616 13806
rect 8668 13524 8720 13530
rect 8772 13512 8800 13806
rect 8720 13484 8800 13512
rect 8668 13466 8720 13472
rect 8864 13410 8892 14350
rect 8956 14074 8984 14350
rect 9140 14334 9260 14362
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 9140 13462 9168 14334
rect 9324 13870 9352 14758
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 8680 13382 8892 13410
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 9232 13394 9260 13670
rect 9310 13560 9366 13569
rect 9310 13495 9366 13504
rect 9220 13388 9272 13394
rect 8484 12436 8536 12442
rect 8036 12406 8156 12434
rect 8128 12306 8156 12406
rect 8484 12378 8536 12384
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8680 12238 8708 13382
rect 9220 13330 9272 13336
rect 9232 13297 9260 13330
rect 9324 13326 9352 13495
rect 9312 13320 9364 13326
rect 9218 13288 9274 13297
rect 9312 13262 9364 13268
rect 9218 13223 9274 13232
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8956 12889 8984 12922
rect 9036 12912 9088 12918
rect 8942 12880 8998 12889
rect 8852 12844 8904 12850
rect 9036 12854 9088 12860
rect 8942 12815 8998 12824
rect 8852 12786 8904 12792
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8772 12442 8800 12650
rect 8864 12442 8892 12786
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 9048 12322 9076 12854
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 8864 12294 9076 12322
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 4250 11996 4558 12005
rect 4250 11994 4256 11996
rect 4312 11994 4336 11996
rect 4392 11994 4416 11996
rect 4472 11994 4496 11996
rect 4552 11994 4558 11996
rect 4312 11942 4314 11994
rect 4494 11942 4496 11994
rect 4250 11940 4256 11942
rect 4312 11940 4336 11942
rect 4392 11940 4416 11942
rect 4472 11940 4496 11942
rect 4552 11940 4558 11942
rect 4250 11931 4558 11940
rect 8864 11914 8892 12294
rect 8944 12096 8996 12102
rect 9140 12050 9168 12650
rect 9232 12306 9260 13223
rect 9416 12986 9444 15524
rect 9548 15535 9550 15544
rect 9496 15506 9548 15512
rect 9680 15506 9732 15512
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9600 15026 9628 15370
rect 9772 15156 9824 15162
rect 9876 15144 9904 16118
rect 9956 15700 10008 15706
rect 10060 15688 10088 16351
rect 10152 16046 10180 16646
rect 10230 16623 10286 16632
rect 10336 16561 10364 19600
rect 10980 16969 11008 19600
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11072 17156 11284 17184
rect 10966 16960 11022 16969
rect 10966 16895 11022 16904
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 10966 16688 11022 16697
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10322 16552 10378 16561
rect 10322 16487 10378 16496
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 10600 16516 10652 16522
rect 10600 16458 10652 16464
rect 10520 16046 10548 16458
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10140 15904 10192 15910
rect 10324 15904 10376 15910
rect 10192 15864 10272 15892
rect 10140 15846 10192 15852
rect 10008 15660 10088 15688
rect 9956 15642 10008 15648
rect 10048 15564 10100 15570
rect 10244 15552 10272 15864
rect 10324 15846 10376 15852
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10336 15706 10364 15846
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10324 15564 10376 15570
rect 10244 15524 10281 15552
rect 10048 15506 10100 15512
rect 10060 15178 10088 15506
rect 10253 15484 10281 15524
rect 10324 15506 10376 15512
rect 10152 15456 10281 15484
rect 10152 15337 10180 15456
rect 10138 15328 10194 15337
rect 10138 15263 10194 15272
rect 10138 15192 10194 15201
rect 10060 15150 10138 15178
rect 9824 15116 9904 15144
rect 10138 15127 10194 15136
rect 10232 15156 10284 15162
rect 9772 15098 9824 15104
rect 10232 15098 10284 15104
rect 9862 15056 9918 15065
rect 9588 15020 9640 15026
rect 10138 15056 10194 15065
rect 9862 14991 9918 15000
rect 9968 15014 10138 15042
rect 9588 14962 9640 14968
rect 9680 14952 9732 14958
rect 9732 14929 9812 14940
rect 9732 14920 9826 14929
rect 9732 14912 9770 14920
rect 9680 14894 9732 14900
rect 9496 14884 9548 14890
rect 9770 14855 9826 14864
rect 9496 14826 9548 14832
rect 9508 14278 9536 14826
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9784 14482 9812 14758
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9876 14074 9904 14991
rect 9968 14958 9996 15014
rect 10138 14991 10194 15000
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9586 13696 9642 13705
rect 9586 13631 9642 13640
rect 9600 13530 9628 13631
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9784 12782 9812 14010
rect 10152 14006 10180 14894
rect 10244 14618 10272 15098
rect 10336 14958 10364 15506
rect 10414 15192 10470 15201
rect 10520 15162 10548 15846
rect 10612 15706 10640 16458
rect 10704 16046 10732 16594
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10704 15570 10732 15982
rect 10888 15706 10916 16662
rect 11072 16658 11100 17156
rect 11256 17066 11284 17156
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 10966 16623 10968 16632
rect 11020 16623 11022 16632
rect 11060 16652 11112 16658
rect 10968 16594 11020 16600
rect 11060 16594 11112 16600
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10980 16250 11008 16458
rect 11164 16266 11192 17002
rect 11348 16658 11376 17274
rect 11520 17128 11572 17134
rect 11440 17088 11520 17116
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11256 16425 11284 16594
rect 11440 16538 11468 17088
rect 11520 17070 11572 17076
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11348 16510 11468 16538
rect 11242 16416 11298 16425
rect 11242 16351 11298 16360
rect 11348 16266 11376 16510
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 11060 16244 11112 16250
rect 11164 16238 11376 16266
rect 11060 16186 11112 16192
rect 10968 16040 11020 16046
rect 10966 16008 10968 16017
rect 11020 16008 11022 16017
rect 10966 15943 11022 15952
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10980 15450 11008 15846
rect 11072 15638 11100 16186
rect 11256 16046 11284 16238
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11334 16008 11390 16017
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15745 11192 15846
rect 11150 15736 11206 15745
rect 11150 15671 11206 15680
rect 11060 15632 11112 15638
rect 11058 15600 11060 15609
rect 11112 15600 11114 15609
rect 11058 15535 11114 15544
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10888 15422 11008 15450
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 10598 15328 10654 15337
rect 10654 15286 10732 15314
rect 10598 15263 10654 15272
rect 10414 15127 10470 15136
rect 10508 15156 10560 15162
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10428 14822 10456 15127
rect 10508 15098 10560 15104
rect 10704 14958 10732 15286
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10690 14784 10746 14793
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10428 14521 10456 14758
rect 10414 14512 10470 14521
rect 10414 14447 10470 14456
rect 10612 14396 10640 14758
rect 10690 14719 10746 14728
rect 10704 14618 10732 14719
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10520 14368 10640 14396
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10060 13394 10088 13670
rect 10152 13530 10180 13738
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9416 12442 9444 12582
rect 9876 12442 9904 13126
rect 10060 12442 10088 13330
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10046 12336 10102 12345
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9404 12300 9456 12306
rect 10046 12271 10048 12280
rect 9404 12242 9456 12248
rect 10100 12271 10102 12280
rect 10048 12242 10100 12248
rect 8996 12044 9168 12050
rect 8944 12038 9168 12044
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 8956 12022 9168 12038
rect 8864 11886 9076 11914
rect 9232 11898 9260 12038
rect 9048 11694 9076 11886
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9416 11762 9444 12242
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 10048 11688 10100 11694
rect 10152 11676 10180 12582
rect 10244 12442 10272 14010
rect 10520 14006 10548 14368
rect 10796 14090 10824 15370
rect 10888 14521 10916 15422
rect 10966 15328 11022 15337
rect 10966 15263 11022 15272
rect 10980 14890 11008 15263
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 11072 14550 11100 15438
rect 11150 14920 11206 14929
rect 11256 14906 11284 15982
rect 11334 15943 11390 15952
rect 11348 15552 11376 15943
rect 11440 15706 11468 16390
rect 11532 16289 11560 16934
rect 11518 16280 11574 16289
rect 11518 16215 11574 16224
rect 11532 16114 11560 16215
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11428 15564 11480 15570
rect 11348 15524 11428 15552
rect 11428 15506 11480 15512
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11206 14878 11284 14906
rect 11334 14920 11390 14929
rect 11150 14855 11206 14864
rect 11334 14855 11390 14864
rect 11348 14822 11376 14855
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11060 14544 11112 14550
rect 10874 14512 10930 14521
rect 11060 14486 11112 14492
rect 10874 14447 10930 14456
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10612 14062 10824 14090
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10508 13388 10560 13394
rect 10612 13376 10640 14062
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10704 13530 10732 13806
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10560 13348 10640 13376
rect 10508 13330 10560 13336
rect 10612 12850 10640 13348
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10324 12300 10376 12306
rect 10428 12288 10456 12718
rect 10796 12374 10824 13942
rect 10888 13870 10916 14350
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10966 13832 11022 13841
rect 10966 13767 11022 13776
rect 10980 12986 11008 13767
rect 11072 13530 11100 14214
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 11348 13444 11376 14554
rect 11256 13416 11376 13444
rect 11256 13258 11284 13416
rect 11440 13376 11468 15302
rect 11532 14958 11560 15846
rect 11624 14958 11652 19600
rect 12268 18737 12296 19600
rect 12912 19530 12940 19600
rect 13004 19530 13032 19638
rect 12912 19502 13032 19530
rect 12254 18728 12310 18737
rect 12254 18663 12310 18672
rect 11955 18524 12263 18533
rect 11955 18522 11961 18524
rect 12017 18522 12041 18524
rect 12097 18522 12121 18524
rect 12177 18522 12201 18524
rect 12257 18522 12263 18524
rect 12017 18470 12019 18522
rect 12199 18470 12201 18522
rect 11955 18468 11961 18470
rect 12017 18468 12041 18470
rect 12097 18468 12121 18470
rect 12177 18468 12201 18470
rect 12257 18468 12263 18470
rect 11955 18459 12263 18468
rect 11955 17436 12263 17445
rect 11955 17434 11961 17436
rect 12017 17434 12041 17436
rect 12097 17434 12121 17436
rect 12177 17434 12201 17436
rect 12257 17434 12263 17436
rect 12017 17382 12019 17434
rect 12199 17382 12201 17434
rect 11955 17380 11961 17382
rect 12017 17380 12041 17382
rect 12097 17380 12121 17382
rect 12177 17380 12201 17382
rect 12257 17380 12263 17382
rect 11955 17371 12263 17380
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 11888 17128 11940 17134
rect 11808 17088 11888 17116
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 15570 11744 16526
rect 11808 15570 11836 17088
rect 11888 17070 11940 17076
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12084 16658 12112 17070
rect 12360 16810 12388 17206
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12360 16782 12480 16810
rect 12452 16658 12480 16782
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 11955 16348 12263 16357
rect 11955 16346 11961 16348
rect 12017 16346 12041 16348
rect 12097 16346 12121 16348
rect 12177 16346 12201 16348
rect 12257 16346 12263 16348
rect 12017 16294 12019 16346
rect 12199 16294 12201 16346
rect 11955 16292 11961 16294
rect 12017 16292 12041 16294
rect 12097 16292 12121 16294
rect 12177 16292 12201 16294
rect 12257 16292 12263 16294
rect 11955 16283 12263 16292
rect 12360 16250 12388 16594
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11900 15638 11928 16118
rect 12452 16114 12480 16390
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 11980 15496 12032 15502
rect 11978 15464 11980 15473
rect 12032 15464 12034 15473
rect 11978 15399 12034 15408
rect 12176 15348 12204 15506
rect 11716 15320 12204 15348
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11716 14464 11744 15320
rect 11955 15260 12263 15269
rect 11955 15258 11961 15260
rect 12017 15258 12041 15260
rect 12097 15258 12121 15260
rect 12177 15258 12201 15260
rect 12257 15258 12263 15260
rect 12017 15206 12019 15258
rect 12199 15206 12201 15258
rect 11955 15204 11961 15206
rect 12017 15204 12041 15206
rect 12097 15204 12121 15206
rect 12177 15204 12201 15206
rect 12257 15204 12263 15206
rect 11955 15195 12263 15204
rect 11796 14884 11848 14890
rect 11796 14826 11848 14832
rect 11532 14436 11744 14464
rect 11532 13734 11560 14436
rect 11612 14340 11664 14346
rect 11612 14282 11664 14288
rect 11624 13870 11652 14282
rect 11808 14090 11836 14826
rect 11955 14172 12263 14181
rect 11955 14170 11961 14172
rect 12017 14170 12041 14172
rect 12097 14170 12121 14172
rect 12177 14170 12201 14172
rect 12257 14170 12263 14172
rect 12017 14118 12019 14170
rect 12199 14118 12201 14170
rect 11955 14116 11961 14118
rect 12017 14116 12041 14118
rect 12097 14116 12121 14118
rect 12177 14116 12201 14118
rect 12257 14116 12263 14118
rect 11955 14107 12263 14116
rect 11704 14068 11756 14074
rect 11808 14062 11928 14090
rect 11704 14010 11756 14016
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11624 13394 11652 13806
rect 11348 13348 11468 13376
rect 11612 13388 11664 13394
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11348 13190 11376 13348
rect 11612 13330 11664 13336
rect 11716 13274 11744 14010
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11440 13246 11744 13274
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11334 13016 11390 13025
rect 10968 12980 11020 12986
rect 11334 12951 11390 12960
rect 10968 12922 11020 12928
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 11072 12306 11100 12854
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 10376 12260 10456 12288
rect 11060 12300 11112 12306
rect 10324 12242 10376 12248
rect 11060 12242 11112 12248
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11898 10732 12038
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10100 11648 10180 11676
rect 10048 11630 10100 11636
rect 7760 11354 7788 11630
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 8102 11452 8410 11461
rect 8102 11450 8108 11452
rect 8164 11450 8188 11452
rect 8244 11450 8268 11452
rect 8324 11450 8348 11452
rect 8404 11450 8410 11452
rect 8164 11398 8166 11450
rect 8346 11398 8348 11450
rect 8102 11396 8108 11398
rect 8164 11396 8188 11398
rect 8244 11396 8268 11398
rect 8324 11396 8348 11398
rect 8404 11396 8410 11398
rect 8102 11387 8410 11396
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 9508 11257 9536 11494
rect 9494 11248 9550 11257
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8484 11212 8536 11218
rect 9494 11183 9550 11192
rect 8484 11154 8536 11160
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 4250 10908 4558 10917
rect 4250 10906 4256 10908
rect 4312 10906 4336 10908
rect 4392 10906 4416 10908
rect 4472 10906 4496 10908
rect 4552 10906 4558 10908
rect 4312 10854 4314 10906
rect 4494 10854 4496 10906
rect 4250 10852 4256 10854
rect 4312 10852 4336 10854
rect 4392 10852 4416 10854
rect 4472 10852 4496 10854
rect 4552 10852 4558 10854
rect 4250 10843 4558 10852
rect 4250 9820 4558 9829
rect 4250 9818 4256 9820
rect 4312 9818 4336 9820
rect 4392 9818 4416 9820
rect 4472 9818 4496 9820
rect 4552 9818 4558 9820
rect 4312 9766 4314 9818
rect 4494 9766 4496 9818
rect 4250 9764 4256 9766
rect 4312 9764 4336 9766
rect 4392 9764 4416 9766
rect 4472 9764 4496 9766
rect 4552 9764 4558 9766
rect 4250 9755 4558 9764
rect 6196 9654 6224 11086
rect 8128 10810 8156 11154
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8496 10674 8524 11154
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 7656 10600 7708 10606
rect 8024 10600 8076 10606
rect 7656 10542 7708 10548
rect 7944 10548 8024 10554
rect 7944 10542 8076 10548
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6460 9512 6512 9518
rect 6458 9480 6460 9489
rect 6512 9480 6514 9489
rect 6458 9415 6514 9424
rect 6656 9178 6684 9862
rect 6748 9518 6776 9930
rect 7208 9722 7236 10066
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7208 9518 7236 9658
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 9178 6776 9318
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 7116 9110 7144 9454
rect 7300 9450 7328 9862
rect 7392 9654 7420 10066
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9722 7512 9862
rect 7576 9722 7604 10066
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7104 9104 7156 9110
rect 7156 9064 7236 9092
rect 7104 9046 7156 9052
rect 4250 8732 4558 8741
rect 4250 8730 4256 8732
rect 4312 8730 4336 8732
rect 4392 8730 4416 8732
rect 4472 8730 4496 8732
rect 4552 8730 4558 8732
rect 4312 8678 4314 8730
rect 4494 8678 4496 8730
rect 4250 8676 4256 8678
rect 4312 8676 4336 8678
rect 4392 8676 4416 8678
rect 4472 8676 4496 8678
rect 4552 8676 4558 8678
rect 4250 8667 4558 8676
rect 7208 8566 7236 9064
rect 7300 8956 7328 9386
rect 7380 8968 7432 8974
rect 7300 8928 7380 8956
rect 7380 8910 7432 8916
rect 7668 8634 7696 10542
rect 7944 10526 8064 10542
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7852 9994 7880 10406
rect 7944 10266 7972 10526
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 10266 8064 10406
rect 8102 10364 8410 10373
rect 8102 10362 8108 10364
rect 8164 10362 8188 10364
rect 8244 10362 8268 10364
rect 8324 10362 8348 10364
rect 8404 10362 8410 10364
rect 8164 10310 8166 10362
rect 8346 10310 8348 10362
rect 8102 10308 8108 10310
rect 8164 10308 8188 10310
rect 8244 10308 8268 10310
rect 8324 10308 8348 10310
rect 8404 10308 8410 10310
rect 8102 10299 8410 10308
rect 8588 10266 8616 11086
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8772 10606 8800 10950
rect 8956 10810 8984 11018
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9140 10810 9168 10950
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9232 10606 9260 11086
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 8772 10266 8800 10406
rect 9048 10266 9076 10406
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9140 10169 9168 10202
rect 9126 10160 9182 10169
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8668 10124 8720 10130
rect 9324 10130 9352 10406
rect 9600 10266 9628 11494
rect 9692 10742 9720 11630
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9126 10095 9182 10104
rect 9312 10124 9364 10130
rect 8668 10066 8720 10072
rect 9312 10066 9364 10072
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 7760 9178 7788 9862
rect 8312 9654 8340 9862
rect 8300 9648 8352 9654
rect 8496 9602 8524 10066
rect 8680 9926 8708 10066
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8300 9590 8352 9596
rect 8404 9574 8524 9602
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7944 9042 7972 9454
rect 8024 9444 8076 9450
rect 8404 9432 8432 9574
rect 8496 9518 8524 9574
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8588 9450 8616 9862
rect 9692 9722 9720 10678
rect 9876 10606 9904 11494
rect 9968 11082 9996 11630
rect 10060 11354 10088 11630
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10140 11280 10192 11286
rect 10060 11228 10140 11234
rect 10060 11222 10192 11228
rect 10060 11206 10180 11222
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 10060 10962 10088 11206
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 9968 10934 10088 10962
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9784 9722 9812 10474
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10266 9904 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 8668 9648 8720 9654
rect 8666 9616 8668 9625
rect 8720 9616 8722 9625
rect 8666 9551 8722 9560
rect 8076 9404 8432 9432
rect 8576 9444 8628 9450
rect 8024 9386 8076 9392
rect 8576 9386 8628 9392
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 8102 9276 8410 9285
rect 8102 9274 8108 9276
rect 8164 9274 8188 9276
rect 8244 9274 8268 9276
rect 8324 9274 8348 9276
rect 8404 9274 8410 9276
rect 8164 9222 8166 9274
rect 8346 9222 8348 9274
rect 8102 9220 8108 9222
rect 8164 9220 8188 9222
rect 8244 9220 8268 9222
rect 8324 9220 8348 9222
rect 8404 9220 8410 9222
rect 8102 9211 8410 9220
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7196 8560 7248 8566
rect 7248 8520 7328 8548
rect 7196 8502 7248 8508
rect 6736 8424 6788 8430
rect 6734 8392 6736 8401
rect 6788 8392 6790 8401
rect 6734 8327 6790 8336
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 4250 7644 4558 7653
rect 4250 7642 4256 7644
rect 4312 7642 4336 7644
rect 4392 7642 4416 7644
rect 4472 7642 4496 7644
rect 4552 7642 4558 7644
rect 4312 7590 4314 7642
rect 4494 7590 4496 7642
rect 4250 7588 4256 7590
rect 4312 7588 4336 7590
rect 4392 7588 4416 7590
rect 4472 7588 4496 7590
rect 4552 7588 4558 7590
rect 4250 7579 4558 7588
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7024 7449 7052 7482
rect 7010 7440 7066 7449
rect 7010 7375 7066 7384
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7104 7336 7156 7342
rect 7208 7324 7236 7686
rect 7300 7342 7328 8520
rect 7668 8430 7696 8570
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7668 8090 7696 8366
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 8090 7788 8230
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7156 7296 7236 7324
rect 7104 7278 7156 7284
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 7002 6960 7142
rect 7024 7002 7052 7278
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 4250 6556 4558 6565
rect 4250 6554 4256 6556
rect 4312 6554 4336 6556
rect 4392 6554 4416 6556
rect 4472 6554 4496 6556
rect 4552 6554 4558 6556
rect 4312 6502 4314 6554
rect 4494 6502 4496 6554
rect 4250 6500 4256 6502
rect 4312 6500 4336 6502
rect 4392 6500 4416 6502
rect 4472 6500 4496 6502
rect 4552 6500 4558 6502
rect 4250 6491 4558 6500
rect 6472 6458 6500 6598
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6564 5710 6592 6802
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 5914 6776 6598
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6840 5710 6868 6802
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 5914 7052 6598
rect 7116 6254 7144 7142
rect 7208 6934 7236 7296
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7208 6254 7236 6598
rect 7300 6458 7328 6598
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7392 6118 7420 6666
rect 7484 6458 7512 6802
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7576 6338 7604 7482
rect 7668 7342 7696 7686
rect 7852 7546 7880 8502
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 6905 7696 7142
rect 7654 6896 7710 6905
rect 7654 6831 7710 6840
rect 7852 6746 7880 7482
rect 7944 6866 7972 8298
rect 8036 8072 8064 8774
rect 8128 8294 8156 8978
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8634 8340 8910
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8116 8288 8168 8294
rect 8404 8276 8432 9114
rect 8772 9110 8800 9318
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8576 9036 8628 9042
rect 8628 8996 8708 9024
rect 8576 8978 8628 8984
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8496 8430 8524 8774
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8404 8248 8524 8276
rect 8116 8230 8168 8236
rect 8102 8188 8410 8197
rect 8102 8186 8108 8188
rect 8164 8186 8188 8188
rect 8244 8186 8268 8188
rect 8324 8186 8348 8188
rect 8404 8186 8410 8188
rect 8164 8134 8166 8186
rect 8346 8134 8348 8186
rect 8102 8132 8108 8134
rect 8164 8132 8188 8134
rect 8244 8132 8268 8134
rect 8324 8132 8348 8134
rect 8404 8132 8410 8134
rect 8102 8123 8410 8132
rect 8496 8090 8524 8248
rect 8484 8084 8536 8090
rect 8036 8044 8156 8072
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8036 7002 8064 7890
rect 8128 7818 8156 8044
rect 8484 8026 8536 8032
rect 8588 7970 8616 8842
rect 8680 8566 8708 8996
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8496 7954 8616 7970
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8484 7948 8616 7954
rect 8536 7942 8616 7948
rect 8484 7890 8536 7896
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8312 7546 8340 7890
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8128 7342 8156 7482
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8102 7100 8410 7109
rect 8102 7098 8108 7100
rect 8164 7098 8188 7100
rect 8244 7098 8268 7100
rect 8324 7098 8348 7100
rect 8404 7098 8410 7100
rect 8164 7046 8166 7098
rect 8346 7046 8348 7098
rect 8102 7044 8108 7046
rect 8164 7044 8188 7046
rect 8244 7044 8268 7046
rect 8324 7044 8348 7046
rect 8404 7044 8410 7046
rect 8102 7035 8410 7044
rect 8496 7002 8524 7210
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8484 6860 8536 6866
rect 8588 6848 8616 7822
rect 8680 6934 8708 8366
rect 8772 8090 8800 8774
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8864 7993 8892 8502
rect 8956 8362 8984 8774
rect 9048 8634 9076 8774
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9140 8514 9168 9318
rect 9692 8906 9720 9658
rect 9770 9480 9826 9489
rect 9770 9415 9772 9424
rect 9824 9415 9826 9424
rect 9772 9386 9824 9392
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9048 8486 9168 8514
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8850 7984 8906 7993
rect 8850 7919 8906 7928
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8772 6934 8800 7346
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8864 6866 8892 7754
rect 8944 7336 8996 7342
rect 9048 7324 9076 8486
rect 9600 8090 9628 8774
rect 9692 8090 9720 8842
rect 9784 8838 9812 8978
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9770 8392 9826 8401
rect 9770 8327 9772 8336
rect 9824 8327 9826 8336
rect 9772 8298 9824 8304
rect 9876 8090 9904 9862
rect 9968 8838 9996 10934
rect 10152 10606 10180 10950
rect 10230 10704 10286 10713
rect 10230 10639 10286 10648
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10244 10470 10272 10639
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10336 9926 10364 10950
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 10060 8634 10088 9454
rect 10336 9382 10364 9862
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10244 9178 10272 9318
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10152 8362 10180 9046
rect 10336 9042 10364 9318
rect 10428 9178 10456 11086
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 10704 10742 10732 10950
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 11072 10266 11100 10950
rect 11164 10606 11192 12650
rect 11256 12442 11284 12718
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11348 11898 11376 12951
rect 11440 12442 11468 13246
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11532 12306 11560 13126
rect 11624 12714 11652 13126
rect 11702 13016 11758 13025
rect 11702 12951 11758 12960
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11624 11354 11652 12242
rect 11716 11898 11744 12951
rect 11808 12434 11836 13942
rect 11900 13938 11928 14062
rect 12360 14056 12388 15846
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12268 14028 12388 14056
rect 12162 13968 12218 13977
rect 11888 13932 11940 13938
rect 12162 13903 12218 13912
rect 11888 13874 11940 13880
rect 12072 13864 12124 13870
rect 12070 13832 12072 13841
rect 12124 13832 12126 13841
rect 12176 13802 12204 13903
rect 12070 13767 12126 13776
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12268 13462 12296 14028
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 11955 13084 12263 13093
rect 11955 13082 11961 13084
rect 12017 13082 12041 13084
rect 12097 13082 12121 13084
rect 12177 13082 12201 13084
rect 12257 13082 12263 13084
rect 12017 13030 12019 13082
rect 12199 13030 12201 13082
rect 11955 13028 11961 13030
rect 12017 13028 12041 13030
rect 12097 13028 12121 13030
rect 12177 13028 12201 13030
rect 12257 13028 12263 13030
rect 11955 13019 12263 13028
rect 11980 12436 12032 12442
rect 11808 12406 11980 12434
rect 12360 12434 12388 13874
rect 12452 13569 12480 15506
rect 12544 15450 12572 16934
rect 12636 16794 12664 17070
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12636 16697 12664 16730
rect 12622 16688 12678 16697
rect 12622 16623 12678 16632
rect 12636 16250 12664 16623
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12820 16046 12848 16390
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12808 16040 12860 16046
rect 13004 16017 13032 17070
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13096 16046 13124 16390
rect 13084 16040 13136 16046
rect 12808 15982 12860 15988
rect 12990 16008 13046 16017
rect 12636 15706 12664 15982
rect 13084 15982 13136 15988
rect 12990 15943 13046 15952
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12544 15422 12664 15450
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12438 13560 12494 13569
rect 12544 13530 12572 15302
rect 12636 15201 12664 15422
rect 12622 15192 12678 15201
rect 12728 15162 12756 15846
rect 12622 15127 12678 15136
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12820 15042 12848 15846
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12992 15564 13044 15570
rect 13188 15552 13216 16390
rect 13280 15892 13308 19638
rect 13542 19600 13598 20000
rect 14186 19600 14242 20000
rect 14830 19600 14886 20000
rect 15474 19600 15530 20000
rect 16118 19600 16174 20000
rect 16762 19600 16818 20000
rect 17406 19600 17462 20000
rect 18050 19600 18106 20000
rect 18694 19600 18750 20000
rect 19338 19600 19394 20000
rect 19982 19600 20038 20000
rect 20626 19600 20682 20000
rect 20732 19638 21220 19666
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13372 16046 13400 16390
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13280 15864 13400 15892
rect 13268 15564 13320 15570
rect 13188 15524 13268 15552
rect 12992 15506 13044 15512
rect 13268 15506 13320 15512
rect 12636 15014 12848 15042
rect 12636 13734 12664 15014
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12438 13495 12494 13504
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12636 12646 12664 12854
rect 12728 12782 12756 13330
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 12434 12664 12582
rect 11980 12378 12032 12384
rect 12084 12406 12388 12434
rect 12452 12406 12664 12434
rect 12716 12436 12768 12442
rect 12084 12306 12112 12406
rect 12452 12306 12480 12406
rect 12716 12378 12768 12384
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 11955 11996 12263 12005
rect 11955 11994 11961 11996
rect 12017 11994 12041 11996
rect 12097 11994 12121 11996
rect 12177 11994 12201 11996
rect 12257 11994 12263 11996
rect 12017 11942 12019 11994
rect 12199 11942 12201 11994
rect 11955 11940 11961 11942
rect 12017 11940 12041 11942
rect 12097 11940 12121 11942
rect 12177 11940 12201 11942
rect 12257 11940 12263 11942
rect 11955 11931 12263 11940
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 12452 11354 12480 12242
rect 12728 12084 12756 12378
rect 12820 12238 12848 14350
rect 12912 13705 12940 15506
rect 13004 14929 13032 15506
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13084 14952 13136 14958
rect 12990 14920 13046 14929
rect 13084 14894 13136 14900
rect 12990 14855 13046 14864
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13004 13870 13032 14758
rect 13096 14618 13124 14894
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 12898 13696 12954 13705
rect 13188 13682 13216 14758
rect 13280 14482 13308 15302
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 12898 13631 12954 13640
rect 13096 13654 13216 13682
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12912 12170 12940 12718
rect 13004 12714 13032 13126
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 12728 12056 12848 12084
rect 12820 12050 12848 12056
rect 13004 12050 13032 12378
rect 13096 12345 13124 13654
rect 13372 13530 13400 15864
rect 13464 14482 13492 16390
rect 13556 16017 13584 19600
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 16658 13768 16934
rect 13832 16794 13860 17070
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13740 16522 13768 16594
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13924 16250 13952 16934
rect 14016 16794 14044 17070
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 14016 16250 14044 16730
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 14094 16144 14150 16153
rect 14094 16079 14150 16088
rect 13542 16008 13598 16017
rect 13542 15943 13598 15952
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13634 15872 13690 15881
rect 13634 15807 13690 15816
rect 13648 15162 13676 15807
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13740 15162 13768 15506
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13832 14958 13860 15914
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13924 15162 13952 15506
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 14108 15042 14136 16079
rect 14200 16028 14228 19600
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 14476 16046 14504 16458
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14464 16040 14516 16046
rect 14200 16000 14412 16028
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 13924 15014 14136 15042
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13556 14346 13584 14758
rect 13648 14482 13860 14498
rect 13648 14476 13872 14482
rect 13648 14470 13820 14476
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13464 12986 13492 13942
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13188 12442 13216 12718
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13082 12336 13138 12345
rect 13280 12306 13308 12582
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13082 12271 13138 12280
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13188 12186 13216 12242
rect 13372 12186 13400 12378
rect 13188 12158 13400 12186
rect 12820 12022 13032 12050
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 13464 11218 13492 12038
rect 13556 11626 13584 13874
rect 13648 13802 13676 14470
rect 13820 14418 13872 14424
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13740 13870 13768 14214
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13648 12918 13676 13738
rect 13832 13394 13860 14282
rect 13924 14006 13952 15014
rect 14004 14884 14056 14890
rect 14004 14826 14056 14832
rect 14016 14414 14044 14826
rect 14200 14482 14228 15302
rect 14292 14822 14320 15370
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14292 14482 14320 14758
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 13530 13952 13670
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 14016 13326 14044 14350
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13636 12912 13688 12918
rect 13636 12854 13688 12860
rect 13924 12306 13952 13194
rect 14016 12714 14044 13262
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13832 11694 13860 12106
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11898 13952 12038
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 14016 11762 14044 12650
rect 14200 12374 14228 14010
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14292 12374 14320 13126
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14108 11762 14136 12242
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 14016 11218 14044 11698
rect 14384 11354 14412 16000
rect 14464 15982 14516 15988
rect 14464 13796 14516 13802
rect 14568 13784 14596 16186
rect 14660 14482 14688 16594
rect 14844 16182 14872 19600
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14936 16794 14964 16934
rect 14924 16788 14976 16794
rect 14924 16730 14976 16736
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14936 16454 14964 16594
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14832 16176 14884 16182
rect 14832 16118 14884 16124
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14752 15638 14780 15846
rect 14844 15706 14872 15846
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14740 15632 14792 15638
rect 14740 15574 14792 15580
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 15028 13977 15056 16458
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15212 14822 15240 16390
rect 15292 16040 15344 16046
rect 15488 15994 15516 19600
rect 16132 19258 16160 19600
rect 16132 19230 16252 19258
rect 15807 19068 16115 19077
rect 15807 19066 15813 19068
rect 15869 19066 15893 19068
rect 15949 19066 15973 19068
rect 16029 19066 16053 19068
rect 16109 19066 16115 19068
rect 15869 19014 15871 19066
rect 16051 19014 16053 19066
rect 15807 19012 15813 19014
rect 15869 19012 15893 19014
rect 15949 19012 15973 19014
rect 16029 19012 16053 19014
rect 16109 19012 16115 19014
rect 15807 19003 16115 19012
rect 15807 17980 16115 17989
rect 15807 17978 15813 17980
rect 15869 17978 15893 17980
rect 15949 17978 15973 17980
rect 16029 17978 16053 17980
rect 16109 17978 16115 17980
rect 15869 17926 15871 17978
rect 16051 17926 16053 17978
rect 15807 17924 15813 17926
rect 15869 17924 15893 17926
rect 15949 17924 15973 17926
rect 16029 17924 16053 17926
rect 16109 17924 16115 17926
rect 15807 17915 16115 17924
rect 15807 16892 16115 16901
rect 15807 16890 15813 16892
rect 15869 16890 15893 16892
rect 15949 16890 15973 16892
rect 16029 16890 16053 16892
rect 16109 16890 16115 16892
rect 15869 16838 15871 16890
rect 16051 16838 16053 16890
rect 15807 16836 15813 16838
rect 15869 16836 15893 16838
rect 15949 16836 15973 16838
rect 16029 16836 16053 16838
rect 16109 16836 16115 16838
rect 15807 16827 16115 16836
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15292 15982 15344 15988
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15014 13968 15070 13977
rect 15014 13903 15070 13912
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14516 13756 14596 13784
rect 14464 13738 14516 13744
rect 14660 13326 14688 13806
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14752 12306 14780 13670
rect 15212 12782 15240 14486
rect 15304 13870 15332 15982
rect 15396 15966 15516 15994
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15304 12918 15332 13806
rect 15396 12986 15424 15966
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 15706 15516 15846
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15488 14618 15516 15370
rect 15580 14890 15608 16662
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15764 16250 15792 16594
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 16132 16046 16160 16526
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 15672 15706 15700 15982
rect 15807 15804 16115 15813
rect 15807 15802 15813 15804
rect 15869 15802 15893 15804
rect 15949 15802 15973 15804
rect 16029 15802 16053 15804
rect 16109 15802 16115 15804
rect 15869 15750 15871 15802
rect 16051 15750 16053 15802
rect 15807 15748 15813 15750
rect 15869 15748 15893 15750
rect 15949 15748 15973 15750
rect 16029 15748 16053 15750
rect 16109 15748 16115 15750
rect 15807 15739 16115 15748
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15807 14716 16115 14725
rect 15807 14714 15813 14716
rect 15869 14714 15893 14716
rect 15949 14714 15973 14716
rect 16029 14714 16053 14716
rect 16109 14714 16115 14716
rect 15869 14662 15871 14714
rect 16051 14662 16053 14714
rect 15807 14660 15813 14662
rect 15869 14660 15893 14662
rect 15949 14660 15973 14662
rect 16029 14660 16053 14662
rect 16109 14660 16115 14662
rect 15807 14651 16115 14660
rect 16224 14618 16252 19230
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 15936 13864 15988 13870
rect 15672 13824 15936 13852
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13190 15516 13670
rect 15672 13530 15700 13824
rect 15936 13806 15988 13812
rect 15807 13628 16115 13637
rect 15807 13626 15813 13628
rect 15869 13626 15893 13628
rect 15949 13626 15973 13628
rect 16029 13626 16053 13628
rect 16109 13626 16115 13628
rect 15869 13574 15871 13626
rect 16051 13574 16053 13626
rect 15807 13572 15813 13574
rect 15869 13572 15893 13574
rect 15949 13572 15973 13574
rect 16029 13572 16053 13574
rect 16109 13572 16115 13574
rect 15807 13563 16115 13572
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 16224 13394 16252 14214
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15016 12232 15068 12238
rect 14936 12180 15016 12186
rect 14936 12174 15068 12180
rect 14936 12158 15056 12174
rect 15108 12164 15160 12170
rect 14936 11830 14964 12158
rect 15108 12106 15160 12112
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 15028 11694 15056 12038
rect 14924 11688 14976 11694
rect 14922 11656 14924 11665
rect 15016 11688 15068 11694
rect 14976 11656 14978 11665
rect 15016 11630 15068 11636
rect 14922 11591 14978 11600
rect 15120 11558 15148 12106
rect 15212 11898 15240 12242
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15198 11792 15254 11801
rect 15198 11727 15254 11736
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11164 10130 11192 10542
rect 11256 10130 11284 10950
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 9178 10548 9318
rect 10704 9178 10732 9590
rect 11072 9518 11100 9862
rect 11348 9654 11376 11018
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11532 10538 11560 10746
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 11624 10198 11652 11018
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11624 9722 11652 10134
rect 11716 10130 11744 11018
rect 11955 10908 12263 10917
rect 11955 10906 11961 10908
rect 12017 10906 12041 10908
rect 12097 10906 12121 10908
rect 12177 10906 12201 10908
rect 12257 10906 12263 10908
rect 12017 10854 12019 10906
rect 12199 10854 12201 10906
rect 11955 10852 11961 10854
rect 12017 10852 12041 10854
rect 12097 10852 12121 10854
rect 12177 10852 12201 10854
rect 12257 10852 12263 10854
rect 11955 10843 12263 10852
rect 12544 10266 12572 11086
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 13266 10976 13322 10985
rect 13004 10266 13032 10950
rect 13266 10911 13322 10920
rect 13280 10810 13308 10911
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 14016 10606 14044 11154
rect 14844 11121 14872 11494
rect 14830 11112 14886 11121
rect 14830 11047 14886 11056
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13372 10266 13400 10474
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10266 13768 10406
rect 13832 10266 13860 10542
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 14108 10130 14136 10950
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15120 10130 15148 10474
rect 15212 10266 15240 11727
rect 15304 11626 15332 12854
rect 15807 12540 16115 12549
rect 15807 12538 15813 12540
rect 15869 12538 15893 12540
rect 15949 12538 15973 12540
rect 16029 12538 16053 12540
rect 16109 12538 16115 12540
rect 15869 12486 15871 12538
rect 16051 12486 16053 12538
rect 15807 12484 15813 12486
rect 15869 12484 15893 12486
rect 15949 12484 15973 12486
rect 16029 12484 16053 12486
rect 16109 12484 16115 12486
rect 15807 12475 16115 12484
rect 16316 12434 16344 16118
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 15570 16712 15846
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16684 14618 16712 15302
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16408 14006 16436 14418
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16408 13802 16436 13942
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16776 13530 16804 19600
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16868 15570 16896 16526
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16868 14618 16896 15506
rect 17144 14890 17172 15846
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17328 14618 17356 15302
rect 17420 15162 17448 19600
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17972 15570 18000 15982
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 16856 14612 16908 14618
rect 17316 14612 17368 14618
rect 16908 14572 16988 14600
rect 16856 14554 16908 14560
rect 16960 14482 16988 14572
rect 17316 14554 17368 14560
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 17512 14278 17540 15370
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17328 14074 17356 14214
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 16948 13796 17000 13802
rect 16948 13738 17000 13744
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16868 12986 16896 13126
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16868 12434 16896 12922
rect 16960 12782 16988 13738
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16224 12406 16344 12434
rect 16408 12406 16896 12434
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15382 11928 15438 11937
rect 15488 11898 15516 12310
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15382 11863 15438 11872
rect 15476 11892 15528 11898
rect 15396 11676 15424 11863
rect 15476 11834 15528 11840
rect 15476 11688 15528 11694
rect 15396 11648 15476 11676
rect 15476 11630 15528 11636
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15384 11212 15436 11218
rect 15488 11200 15516 11494
rect 15580 11354 15608 12038
rect 15672 11898 15700 12242
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15658 11792 15714 11801
rect 15658 11727 15660 11736
rect 15712 11727 15714 11736
rect 15660 11698 15712 11704
rect 15764 11642 15792 12242
rect 15856 11801 15884 12242
rect 15842 11792 15898 11801
rect 15842 11727 15898 11736
rect 15844 11688 15896 11694
rect 15764 11636 15844 11642
rect 15764 11630 15896 11636
rect 15764 11614 15884 11630
rect 15856 11540 15884 11614
rect 15672 11512 15884 11540
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15488 11172 15608 11200
rect 15384 11154 15436 11160
rect 15304 10266 15332 11154
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 13912 10124 13964 10130
rect 14096 10124 14148 10130
rect 13964 10084 14044 10112
rect 13912 10066 13964 10072
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11716 9722 11744 9862
rect 11808 9722 11836 9862
rect 11955 9820 12263 9829
rect 11955 9818 11961 9820
rect 12017 9818 12041 9820
rect 12097 9818 12121 9820
rect 12177 9818 12201 9820
rect 12257 9818 12263 9820
rect 12017 9766 12019 9818
rect 12199 9766 12201 9818
rect 11955 9764 11961 9766
rect 12017 9764 12041 9766
rect 12097 9764 12121 9766
rect 12177 9764 12201 9766
rect 12257 9764 12263 9766
rect 11955 9755 12263 9764
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11624 9602 11652 9658
rect 12360 9654 12388 10066
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 11888 9648 11940 9654
rect 11624 9596 11888 9602
rect 11624 9590 11940 9596
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 11624 9574 11928 9590
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 9217 11376 9318
rect 11334 9208 11390 9217
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10692 9172 10744 9178
rect 11334 9143 11390 9152
rect 10692 9114 10744 9120
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7410 9168 7686
rect 9220 7472 9272 7478
rect 9272 7420 9444 7426
rect 9220 7414 9444 7420
rect 9128 7404 9180 7410
rect 9232 7398 9444 7414
rect 9128 7346 9180 7352
rect 8996 7296 9076 7324
rect 9220 7336 9272 7342
rect 9218 7304 9220 7313
rect 9312 7336 9364 7342
rect 9272 7304 9274 7313
rect 8944 7278 8996 7284
rect 9312 7278 9364 7284
rect 9218 7239 9274 7248
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 6866 9260 7142
rect 8536 6820 8616 6848
rect 8852 6860 8904 6866
rect 8484 6802 8536 6808
rect 8852 6802 8904 6808
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 8220 6746 8248 6802
rect 7852 6718 8248 6746
rect 8392 6792 8444 6798
rect 8760 6792 8812 6798
rect 8444 6740 8760 6746
rect 8392 6734 8812 6740
rect 8404 6718 8800 6734
rect 8220 6458 8248 6718
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 7576 6310 8064 6338
rect 8036 6254 8064 6310
rect 9324 6254 9352 7278
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 8024 6248 8076 6254
rect 9312 6248 9364 6254
rect 8024 6190 8076 6196
rect 9034 6216 9090 6225
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7852 5914 7880 6190
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8944 6180 8996 6186
rect 9312 6190 9364 6196
rect 9034 6151 9036 6160
rect 8944 6122 8996 6128
rect 9088 6151 9090 6160
rect 9036 6122 9088 6128
rect 8102 6012 8410 6021
rect 8102 6010 8108 6012
rect 8164 6010 8188 6012
rect 8244 6010 8268 6012
rect 8324 6010 8348 6012
rect 8404 6010 8410 6012
rect 8164 5958 8166 6010
rect 8346 5958 8348 6010
rect 8102 5956 8108 5958
rect 8164 5956 8188 5958
rect 8244 5956 8268 5958
rect 8324 5956 8348 5958
rect 8404 5956 8410 5958
rect 8102 5947 8410 5956
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 4250 5468 4558 5477
rect 4250 5466 4256 5468
rect 4312 5466 4336 5468
rect 4392 5466 4416 5468
rect 4472 5466 4496 5468
rect 4552 5466 4558 5468
rect 4312 5414 4314 5466
rect 4494 5414 4496 5466
rect 4250 5412 4256 5414
rect 4312 5412 4336 5414
rect 4392 5412 4416 5414
rect 4472 5412 4496 5414
rect 4552 5412 4558 5414
rect 4250 5403 4558 5412
rect 8392 5160 8444 5166
rect 8496 5148 8524 5850
rect 8588 5778 8616 6122
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8444 5120 8524 5148
rect 8392 5102 8444 5108
rect 8102 4924 8410 4933
rect 8102 4922 8108 4924
rect 8164 4922 8188 4924
rect 8244 4922 8268 4924
rect 8324 4922 8348 4924
rect 8404 4922 8410 4924
rect 8164 4870 8166 4922
rect 8346 4870 8348 4922
rect 8102 4868 8108 4870
rect 8164 4868 8188 4870
rect 8244 4868 8268 4870
rect 8324 4868 8348 4870
rect 8404 4868 8410 4870
rect 8102 4859 8410 4868
rect 4250 4380 4558 4389
rect 4250 4378 4256 4380
rect 4312 4378 4336 4380
rect 4392 4378 4416 4380
rect 4472 4378 4496 4380
rect 4552 4378 4558 4380
rect 4312 4326 4314 4378
rect 4494 4326 4496 4378
rect 4250 4324 4256 4326
rect 4312 4324 4336 4326
rect 4392 4324 4416 4326
rect 4472 4324 4496 4326
rect 4552 4324 4558 4326
rect 4250 4315 4558 4324
rect 8496 4146 8524 5120
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8102 3836 8410 3845
rect 8102 3834 8108 3836
rect 8164 3834 8188 3836
rect 8244 3834 8268 3836
rect 8324 3834 8348 3836
rect 8404 3834 8410 3836
rect 8164 3782 8166 3834
rect 8346 3782 8348 3834
rect 8102 3780 8108 3782
rect 8164 3780 8188 3782
rect 8244 3780 8268 3782
rect 8324 3780 8348 3782
rect 8404 3780 8410 3782
rect 8102 3771 8410 3780
rect 8496 3602 8524 4082
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 4250 3292 4558 3301
rect 4250 3290 4256 3292
rect 4312 3290 4336 3292
rect 4392 3290 4416 3292
rect 4472 3290 4496 3292
rect 4552 3290 4558 3292
rect 4312 3238 4314 3290
rect 4494 3238 4496 3290
rect 4250 3236 4256 3238
rect 4312 3236 4336 3238
rect 4392 3236 4416 3238
rect 4472 3236 4496 3238
rect 4552 3236 4558 3238
rect 4250 3227 4558 3236
rect 8102 2748 8410 2757
rect 8102 2746 8108 2748
rect 8164 2746 8188 2748
rect 8244 2746 8268 2748
rect 8324 2746 8348 2748
rect 8404 2746 8410 2748
rect 8164 2694 8166 2746
rect 8346 2694 8348 2746
rect 8102 2692 8108 2694
rect 8164 2692 8188 2694
rect 8244 2692 8268 2694
rect 8324 2692 8348 2694
rect 8404 2692 8410 2694
rect 8102 2683 8410 2692
rect 4250 2204 4558 2213
rect 4250 2202 4256 2204
rect 4312 2202 4336 2204
rect 4392 2202 4416 2204
rect 4472 2202 4496 2204
rect 4552 2202 4558 2204
rect 4312 2150 4314 2202
rect 4494 2150 4496 2202
rect 4250 2148 4256 2150
rect 4312 2148 4336 2150
rect 4392 2148 4416 2150
rect 4472 2148 4496 2150
rect 4552 2148 4558 2150
rect 4250 2139 4558 2148
rect 8102 1660 8410 1669
rect 8102 1658 8108 1660
rect 8164 1658 8188 1660
rect 8244 1658 8268 1660
rect 8324 1658 8348 1660
rect 8404 1658 8410 1660
rect 8164 1606 8166 1658
rect 8346 1606 8348 1658
rect 8102 1604 8108 1606
rect 8164 1604 8188 1606
rect 8244 1604 8268 1606
rect 8324 1604 8348 1606
rect 8404 1604 8410 1606
rect 8102 1595 8410 1604
rect 4250 1116 4558 1125
rect 4250 1114 4256 1116
rect 4312 1114 4336 1116
rect 4392 1114 4416 1116
rect 4472 1114 4496 1116
rect 4552 1114 4558 1116
rect 4312 1062 4314 1114
rect 4494 1062 4496 1114
rect 4250 1060 4256 1062
rect 4312 1060 4336 1062
rect 4392 1060 4416 1062
rect 4472 1060 4496 1062
rect 4552 1060 4558 1062
rect 4250 1051 4558 1060
rect 8680 1018 8708 5646
rect 8772 4622 8800 6054
rect 8956 5914 8984 6122
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9048 5778 9076 6122
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9232 5914 9260 6054
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9324 4826 9352 6190
rect 9416 5234 9444 7398
rect 9508 7342 9536 7754
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7546 9628 7686
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9496 7336 9548 7342
rect 9600 7313 9628 7346
rect 9496 7278 9548 7284
rect 9586 7304 9642 7313
rect 9586 7239 9642 7248
rect 9692 7002 9720 8026
rect 10060 7886 10088 8230
rect 10336 7954 10364 8774
rect 10888 8634 10916 8910
rect 11532 8906 11560 9454
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11716 9178 11744 9318
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11900 9110 11928 9454
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11955 8732 12263 8741
rect 11955 8730 11961 8732
rect 12017 8730 12041 8732
rect 12097 8730 12121 8732
rect 12177 8730 12201 8732
rect 12257 8730 12263 8732
rect 12017 8678 12019 8730
rect 12199 8678 12201 8730
rect 11955 8676 11961 8678
rect 12017 8676 12041 8678
rect 12097 8676 12121 8678
rect 12177 8676 12201 8678
rect 12257 8676 12263 8678
rect 11955 8667 12263 8676
rect 12636 8634 12664 9454
rect 12912 9382 12940 9862
rect 13004 9586 13032 9862
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12714 9072 12770 9081
rect 13096 9042 13124 9998
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 12714 9007 12716 9016
rect 12768 9007 12770 9016
rect 13084 9036 13136 9042
rect 12716 8978 12768 8984
rect 13084 8978 13136 8984
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 10416 8424 10468 8430
rect 10600 8424 10652 8430
rect 10468 8384 10600 8412
rect 10416 8366 10468 8372
rect 10600 8366 10652 8372
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10612 8090 10640 8230
rect 10704 8090 10732 8570
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9876 7410 9904 7686
rect 10138 7440 10194 7449
rect 9864 7404 9916 7410
rect 10138 7375 10194 7384
rect 9864 7346 9916 7352
rect 10152 7342 10180 7375
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 9784 7002 9812 7278
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9508 5914 9536 6326
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9600 5370 9628 6666
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9692 5778 9720 6326
rect 9784 6225 9812 6666
rect 9876 6390 9904 7210
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10152 6458 10180 6734
rect 10244 6458 10272 7890
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10322 6896 10378 6905
rect 10428 6866 10456 7210
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 7002 10548 7142
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10322 6831 10378 6840
rect 10416 6860 10468 6866
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10232 6452 10284 6458
rect 10336 6440 10364 6831
rect 10416 6802 10468 6808
rect 10704 6730 10732 8026
rect 10796 7954 10824 8502
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10612 6458 10640 6666
rect 10600 6452 10652 6458
rect 10336 6412 10456 6440
rect 10232 6394 10284 6400
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10048 6248 10100 6254
rect 9770 6216 9826 6225
rect 10048 6190 10100 6196
rect 9770 6151 9826 6160
rect 10060 5914 10088 6190
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9680 5568 9732 5574
rect 10152 5534 10180 6258
rect 9680 5510 9732 5516
rect 9692 5370 9720 5510
rect 10060 5506 10180 5534
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 10060 5166 10088 5506
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9324 4729 9352 4762
rect 9784 4758 9812 4966
rect 9772 4752 9824 4758
rect 9310 4720 9366 4729
rect 9772 4694 9824 4700
rect 10060 4690 10088 5102
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10152 4826 10180 4966
rect 10336 4826 10364 6258
rect 10428 5098 10456 6412
rect 10600 6394 10652 6400
rect 10704 6322 10732 6666
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10796 6254 10824 7890
rect 11164 7818 11192 8366
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10612 4690 10640 6054
rect 10888 5710 10916 7142
rect 11072 7002 11100 7142
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11164 6798 11192 7754
rect 11348 7546 11376 8366
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10876 5092 10928 5098
rect 10876 5034 10928 5040
rect 10888 4826 10916 5034
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10690 4720 10746 4729
rect 9310 4655 9366 4664
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10600 4684 10652 4690
rect 10690 4655 10692 4664
rect 10600 4626 10652 4632
rect 10744 4655 10746 4664
rect 10692 4626 10744 4632
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4282 9352 4422
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9508 4214 9536 4626
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8772 3670 8800 3878
rect 9876 3738 9904 4150
rect 10152 4078 10180 4626
rect 10520 4078 10548 4626
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10152 3738 10180 4014
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10244 3670 10272 3878
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8668 1012 8720 1018
rect 8668 954 8720 960
rect 7840 808 7892 814
rect 7840 750 7892 756
rect 7852 490 7880 750
rect 8102 572 8410 581
rect 8102 570 8108 572
rect 8164 570 8188 572
rect 8244 570 8268 572
rect 8324 570 8348 572
rect 8404 570 8410 572
rect 8164 518 8166 570
rect 8346 518 8348 570
rect 8102 516 8108 518
rect 8164 516 8188 518
rect 8244 516 8268 518
rect 8324 516 8348 518
rect 8404 516 8410 518
rect 8102 507 8410 516
rect 7760 462 7880 490
rect 7760 400 7788 462
rect 8312 428 8432 456
rect 7746 0 7802 400
rect 8312 377 8340 428
rect 8404 400 8432 428
rect 9048 400 9076 3538
rect 10520 3466 10548 4014
rect 10612 3942 10640 4490
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9692 400 9720 2790
rect 10336 400 10364 3334
rect 10980 400 11008 5578
rect 11072 5370 11100 6258
rect 11164 6254 11192 6734
rect 11256 6458 11284 7346
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 6934 11376 7142
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11440 6866 11468 8298
rect 11532 8022 11560 8366
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11716 7818 11744 8366
rect 12912 8022 12940 8434
rect 13096 8362 13124 8978
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13188 8566 13216 8774
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 13280 8430 13308 9114
rect 13372 8430 13400 9318
rect 13450 9208 13506 9217
rect 13506 9178 13584 9194
rect 13740 9178 13768 9454
rect 13506 9172 13596 9178
rect 13506 9166 13544 9172
rect 13450 9143 13506 9152
rect 13544 9114 13596 9120
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13832 8430 13860 9930
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13924 9722 13952 9862
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14016 9674 14044 10084
rect 14372 10124 14424 10130
rect 14148 10084 14228 10112
rect 14096 10066 14148 10072
rect 14016 9646 14136 9674
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13924 9178 13952 9522
rect 14108 9518 14136 9646
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14200 9330 14228 10084
rect 14372 10066 14424 10072
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 14384 9722 14412 10066
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14660 9654 14688 10066
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14660 9518 14688 9590
rect 14752 9518 14780 9862
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14108 9302 14228 9330
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 14108 8838 14136 9302
rect 15028 8974 15056 9998
rect 15120 9042 15148 10066
rect 15396 9926 15424 11154
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15488 10033 15516 11018
rect 15580 10282 15608 11172
rect 15672 10606 15700 11512
rect 15807 11452 16115 11461
rect 15807 11450 15813 11452
rect 15869 11450 15893 11452
rect 15949 11450 15973 11452
rect 16029 11450 16053 11452
rect 16109 11450 16115 11452
rect 15869 11398 15871 11450
rect 16051 11398 16053 11450
rect 15807 11396 15813 11398
rect 15869 11396 15893 11398
rect 15949 11396 15973 11398
rect 16029 11396 16053 11398
rect 16109 11396 16115 11398
rect 15807 11387 16115 11396
rect 16118 11248 16174 11257
rect 16118 11183 16120 11192
rect 16172 11183 16174 11192
rect 16120 11154 16172 11160
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15856 10810 15884 10950
rect 16224 10810 16252 12406
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16316 11354 16344 12106
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 10441 15700 10542
rect 16212 10464 16264 10470
rect 15658 10432 15714 10441
rect 16212 10406 16264 10412
rect 15658 10367 15714 10376
rect 15807 10364 16115 10373
rect 15807 10362 15813 10364
rect 15869 10362 15893 10364
rect 15949 10362 15973 10364
rect 16029 10362 16053 10364
rect 16109 10362 16115 10364
rect 15869 10310 15871 10362
rect 16051 10310 16053 10362
rect 15807 10308 15813 10310
rect 15869 10308 15893 10310
rect 15949 10308 15973 10310
rect 16029 10308 16053 10310
rect 16109 10308 16115 10310
rect 15807 10299 16115 10308
rect 15580 10254 15700 10282
rect 16224 10266 16252 10406
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15474 10024 15530 10033
rect 15474 9959 15530 9968
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14108 8566 14136 8774
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14476 8430 14504 8774
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 11955 7644 12263 7653
rect 11955 7642 11961 7644
rect 12017 7642 12041 7644
rect 12097 7642 12121 7644
rect 12177 7642 12201 7644
rect 12257 7642 12263 7644
rect 12017 7590 12019 7642
rect 12199 7590 12201 7642
rect 11955 7588 11961 7590
rect 12017 7588 12041 7590
rect 12097 7588 12121 7590
rect 12177 7588 12201 7590
rect 12257 7588 12263 7590
rect 11955 7579 12263 7588
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11532 7041 11560 7142
rect 11518 7032 11574 7041
rect 11518 6967 11574 6976
rect 11716 6934 11744 7346
rect 12636 7342 12664 7686
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11348 4826 11376 5714
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11440 4690 11468 5646
rect 11532 5166 11560 6666
rect 11808 6338 11836 7142
rect 12544 7018 12572 7278
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12544 6990 12664 7018
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12268 6662 12296 6802
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 11955 6556 12263 6565
rect 11955 6554 11961 6556
rect 12017 6554 12041 6556
rect 12097 6554 12121 6556
rect 12177 6554 12201 6556
rect 12257 6554 12263 6556
rect 12017 6502 12019 6554
rect 12199 6502 12201 6554
rect 11955 6500 11961 6502
rect 12017 6500 12041 6502
rect 12097 6500 12121 6502
rect 12177 6500 12201 6502
rect 12257 6500 12263 6502
rect 11955 6491 12263 6500
rect 11716 6310 11836 6338
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 4758 11560 5102
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11440 4078 11468 4490
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11624 400 11652 4966
rect 11716 2854 11744 6310
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11808 4826 11836 6122
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12268 5658 12296 6054
rect 12360 5914 12388 6666
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12268 5630 12388 5658
rect 11955 5468 12263 5477
rect 11955 5466 11961 5468
rect 12017 5466 12041 5468
rect 12097 5466 12121 5468
rect 12177 5466 12201 5468
rect 12257 5466 12263 5468
rect 12017 5414 12019 5466
rect 12199 5414 12201 5466
rect 11955 5412 11961 5414
rect 12017 5412 12041 5414
rect 12097 5412 12121 5414
rect 12177 5412 12201 5414
rect 12257 5412 12263 5414
rect 11955 5403 12263 5412
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11808 4282 11836 4422
rect 11955 4380 12263 4389
rect 11955 4378 11961 4380
rect 12017 4378 12041 4380
rect 12097 4378 12121 4380
rect 12177 4378 12201 4380
rect 12257 4378 12263 4380
rect 12017 4326 12019 4378
rect 12199 4326 12201 4378
rect 11955 4324 11961 4326
rect 12017 4324 12041 4326
rect 12097 4324 12121 4326
rect 12177 4324 12201 4326
rect 12257 4324 12263 4326
rect 11955 4315 12263 4324
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11955 3292 12263 3301
rect 11955 3290 11961 3292
rect 12017 3290 12041 3292
rect 12097 3290 12121 3292
rect 12177 3290 12201 3292
rect 12257 3290 12263 3292
rect 12017 3238 12019 3290
rect 12199 3238 12201 3290
rect 11955 3236 11961 3238
rect 12017 3236 12041 3238
rect 12097 3236 12121 3238
rect 12177 3236 12201 3238
rect 12257 3236 12263 3238
rect 11955 3227 12263 3236
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11955 2204 12263 2213
rect 11955 2202 11961 2204
rect 12017 2202 12041 2204
rect 12097 2202 12121 2204
rect 12177 2202 12201 2204
rect 12257 2202 12263 2204
rect 12017 2150 12019 2202
rect 12199 2150 12201 2202
rect 11955 2148 11961 2150
rect 12017 2148 12041 2150
rect 12097 2148 12121 2150
rect 12177 2148 12201 2150
rect 12257 2148 12263 2150
rect 11955 2139 12263 2148
rect 11955 1116 12263 1125
rect 11955 1114 11961 1116
rect 12017 1114 12041 1116
rect 12097 1114 12121 1116
rect 12177 1114 12201 1116
rect 12257 1114 12263 1116
rect 12017 1062 12019 1114
rect 12199 1062 12201 1114
rect 11955 1060 11961 1062
rect 12017 1060 12041 1062
rect 12097 1060 12121 1062
rect 12177 1060 12201 1062
rect 12257 1060 12263 1062
rect 11955 1051 12263 1060
rect 12360 898 12388 5630
rect 12544 5370 12572 6802
rect 12636 6118 12664 6990
rect 12728 6458 12756 7210
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12728 4554 12756 5102
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12820 3602 12848 5646
rect 13004 5534 13032 8230
rect 13280 7954 13308 8366
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13740 8022 13768 8230
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13188 6662 13216 7686
rect 13280 7342 13308 7890
rect 13740 7342 13768 7958
rect 13924 7342 13952 8298
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14292 7342 14320 7686
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13728 7336 13780 7342
rect 13912 7336 13964 7342
rect 13780 7296 13860 7324
rect 13728 7278 13780 7284
rect 13648 6798 13676 7278
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13188 6254 13216 6598
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13648 6118 13676 6734
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5846 13676 6054
rect 13636 5840 13688 5846
rect 13636 5782 13688 5788
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 12912 5506 13032 5534
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12268 870 12388 898
rect 12268 400 12296 870
rect 12912 400 12940 5506
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13096 4826 13124 5306
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4826 13308 4966
rect 13556 4826 13584 5714
rect 13740 5534 13768 6598
rect 13832 6254 13860 7296
rect 13912 7278 13964 7284
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 13924 6322 13952 7278
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13648 5506 13768 5534
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 13004 3942 13032 4626
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3602 13032 3878
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13648 2258 13676 5506
rect 13832 4622 13860 5850
rect 14108 5534 14136 7142
rect 14108 5506 14228 5534
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13924 4672 13952 5102
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14108 4826 14136 5034
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14200 4758 14228 5506
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14096 4684 14148 4690
rect 13924 4644 14096 4672
rect 14096 4626 14148 4632
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 14108 3670 14136 4626
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14200 4078 14228 4422
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14292 3738 14320 4626
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 14384 2802 14412 7686
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14476 6066 14504 7414
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14568 7002 14596 7278
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14476 6038 14596 6066
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14476 5166 14504 5850
rect 14568 5545 14596 6038
rect 14554 5536 14610 5545
rect 14554 5471 14610 5480
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14568 5030 14596 5306
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14660 4826 14688 7210
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 13556 2230 13676 2258
rect 14200 2774 14412 2802
rect 14752 2802 14780 8774
rect 15212 8401 15240 9386
rect 15304 9178 15332 9862
rect 15580 9722 15608 10066
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15566 9616 15622 9625
rect 15566 9551 15568 9560
rect 15620 9551 15622 9560
rect 15568 9522 15620 9528
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15580 9042 15608 9318
rect 15672 9178 15700 10254
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 15934 10160 15990 10169
rect 15934 10095 15990 10104
rect 16304 10124 16356 10130
rect 15844 10056 15896 10062
rect 15842 10024 15844 10033
rect 15896 10024 15898 10033
rect 15752 9988 15804 9994
rect 15842 9959 15898 9968
rect 15752 9930 15804 9936
rect 15764 9518 15792 9930
rect 15948 9518 15976 10095
rect 16408 10112 16436 12406
rect 16868 12102 16896 12406
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16500 11354 16528 12038
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 16684 11642 16712 11766
rect 16592 11614 16712 11642
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16500 11121 16528 11154
rect 16486 11112 16542 11121
rect 16486 11047 16542 11056
rect 16592 10810 16620 11614
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16684 10470 16712 11494
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16776 10266 16804 10950
rect 16868 10810 16896 11086
rect 16960 11082 16988 12718
rect 17052 11762 17080 12718
rect 17144 12714 17172 13670
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 17144 11937 17172 12106
rect 17130 11928 17186 11937
rect 17236 11898 17264 13806
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17604 12306 17632 13398
rect 17696 12986 17724 13806
rect 17788 13394 17816 14894
rect 17972 14482 18000 15506
rect 18064 14634 18092 19600
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18248 15552 18276 16186
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18340 15706 18368 15982
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18432 15638 18460 15846
rect 18420 15632 18472 15638
rect 18420 15574 18472 15580
rect 18328 15564 18380 15570
rect 18248 15524 18328 15552
rect 18328 15506 18380 15512
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18156 14958 18184 15302
rect 18340 15162 18368 15506
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18064 14606 18184 14634
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18064 14074 18092 14418
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17972 13394 18000 14010
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 13530 18092 13806
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17788 12782 17816 13330
rect 18156 12986 18184 14606
rect 18340 14482 18368 15098
rect 18604 15088 18656 15094
rect 18602 15056 18604 15065
rect 18656 15056 18658 15065
rect 18602 14991 18658 15000
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18328 14476 18380 14482
rect 18248 14436 18328 14464
rect 18248 13870 18276 14436
rect 18328 14418 18380 14424
rect 18432 14396 18460 14486
rect 18604 14408 18656 14414
rect 18432 14368 18552 14396
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 18340 13870 18368 14282
rect 18524 14278 18552 14368
rect 18604 14350 18656 14356
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18432 13530 18460 14214
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17788 12442 17816 12718
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 18616 12374 18644 14350
rect 18604 12368 18656 12374
rect 18510 12336 18566 12345
rect 17592 12300 17644 12306
rect 18604 12310 18656 12316
rect 18510 12271 18566 12280
rect 17592 12242 17644 12248
rect 17130 11863 17186 11872
rect 17224 11892 17276 11898
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 17052 10674 17080 11698
rect 17144 11014 17172 11863
rect 17224 11834 17276 11840
rect 17236 11354 17264 11834
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 17052 10130 17080 10610
rect 17144 10606 17172 10950
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17144 10130 17172 10406
rect 16356 10084 16436 10112
rect 17040 10124 17092 10130
rect 16304 10066 16356 10072
rect 17040 10066 17092 10072
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15807 9276 16115 9285
rect 15807 9274 15813 9276
rect 15869 9274 15893 9276
rect 15949 9274 15973 9276
rect 16029 9274 16053 9276
rect 16109 9274 16115 9276
rect 15869 9222 15871 9274
rect 16051 9222 16053 9274
rect 15807 9220 15813 9222
rect 15869 9220 15893 9222
rect 15949 9220 15973 9222
rect 16029 9220 16053 9222
rect 16109 9220 16115 9222
rect 15807 9211 16115 9220
rect 16500 9178 16528 9862
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16960 9042 16988 9386
rect 17328 9178 17356 10066
rect 17604 9654 17632 12242
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 18064 11354 18092 12038
rect 18524 11898 18552 12271
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18234 11792 18290 11801
rect 18234 11727 18290 11736
rect 18248 11354 18276 11727
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15580 8634 15608 8774
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 16764 8628 16816 8634
rect 16816 8588 16988 8616
rect 16764 8570 16816 8576
rect 16856 8424 16908 8430
rect 15198 8392 15254 8401
rect 16856 8366 16908 8372
rect 15198 8327 15254 8336
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15304 8022 15332 8298
rect 15807 8188 16115 8197
rect 15807 8186 15813 8188
rect 15869 8186 15893 8188
rect 15949 8186 15973 8188
rect 16029 8186 16053 8188
rect 16109 8186 16115 8188
rect 15869 8134 15871 8186
rect 16051 8134 16053 8186
rect 15807 8132 15813 8134
rect 15869 8132 15893 8134
rect 15949 8132 15973 8134
rect 16029 8132 16053 8134
rect 16109 8132 16115 8134
rect 15807 8123 16115 8132
rect 15292 8016 15344 8022
rect 15292 7958 15344 7964
rect 16868 7954 16896 8366
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 14844 7290 14872 7890
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 14844 7262 15056 7290
rect 14832 7200 14884 7206
rect 14830 7168 14832 7177
rect 14924 7200 14976 7206
rect 14884 7168 14886 7177
rect 14924 7142 14976 7148
rect 14830 7103 14886 7112
rect 14936 6866 14964 7142
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14844 4690 14872 6802
rect 15028 6474 15056 7262
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 14936 6446 15056 6474
rect 14936 5166 14964 6446
rect 15212 6254 15240 7142
rect 15304 6474 15332 7482
rect 15580 7342 15608 7754
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15856 7546 15884 7686
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 15396 7002 15424 7210
rect 15474 7168 15530 7177
rect 15474 7103 15530 7112
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15382 6896 15438 6905
rect 15488 6866 15516 7103
rect 15382 6831 15438 6840
rect 15476 6860 15528 6866
rect 15396 6610 15424 6831
rect 15476 6802 15528 6808
rect 15568 6656 15620 6662
rect 15396 6582 15516 6610
rect 15568 6598 15620 6604
rect 15304 6446 15424 6474
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 15028 5409 15056 5714
rect 15106 5536 15162 5545
rect 15106 5471 15162 5480
rect 15014 5400 15070 5409
rect 15014 5335 15070 5344
rect 15120 5216 15148 5471
rect 15028 5188 15148 5216
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14922 4992 14978 5001
rect 14922 4927 14978 4936
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14936 4146 14964 4927
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 15028 3602 15056 5188
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 15120 4842 15148 5034
rect 15212 5030 15240 6054
rect 15304 5166 15332 6326
rect 15396 5166 15424 6446
rect 15488 5370 15516 6582
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15396 4842 15424 4966
rect 15120 4814 15424 4842
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15304 3466 15332 4218
rect 15396 3670 15424 4814
rect 15488 4690 15516 5170
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15292 3460 15344 3466
rect 15292 3402 15344 3408
rect 14752 2774 14872 2802
rect 15580 2774 15608 6598
rect 15672 6118 15700 7210
rect 15807 7100 16115 7109
rect 15807 7098 15813 7100
rect 15869 7098 15893 7100
rect 15949 7098 15973 7100
rect 16029 7098 16053 7100
rect 16109 7098 16115 7100
rect 15869 7046 15871 7098
rect 16051 7046 16053 7098
rect 15807 7044 15813 7046
rect 15869 7044 15893 7046
rect 15949 7044 15973 7046
rect 16029 7044 16053 7046
rect 16109 7044 16115 7046
rect 15807 7035 16115 7044
rect 16224 6934 16252 7890
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16316 7410 16344 7686
rect 16500 7478 16528 7686
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16684 7342 16712 7686
rect 16868 7546 16896 7890
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16776 7002 16804 7346
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16776 6458 16804 6802
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16868 6254 16896 7482
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15807 6012 16115 6021
rect 15807 6010 15813 6012
rect 15869 6010 15893 6012
rect 15949 6010 15973 6012
rect 16029 6010 16053 6012
rect 16109 6010 16115 6012
rect 15869 5958 15871 6010
rect 16051 5958 16053 6010
rect 15807 5956 15813 5958
rect 15869 5956 15893 5958
rect 15949 5956 15973 5958
rect 16029 5956 16053 5958
rect 16109 5956 16115 5958
rect 15807 5947 16115 5956
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15672 4554 15700 5714
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 16040 5166 16068 5238
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 16040 5030 16068 5102
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 15807 4924 16115 4933
rect 15807 4922 15813 4924
rect 15869 4922 15893 4924
rect 15949 4922 15973 4924
rect 16029 4922 16053 4924
rect 16109 4922 16115 4924
rect 15869 4870 15871 4922
rect 16051 4870 16053 4922
rect 15807 4868 15813 4870
rect 15869 4868 15893 4870
rect 15949 4868 15973 4870
rect 16029 4868 16053 4870
rect 16109 4868 16115 4870
rect 15807 4859 16115 4868
rect 16224 4826 16252 5034
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15856 4486 15884 4626
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15856 4282 15884 4422
rect 15948 4298 15976 4626
rect 15844 4276 15896 4282
rect 15948 4270 16252 4298
rect 15844 4218 15896 4224
rect 15807 3836 16115 3845
rect 15807 3834 15813 3836
rect 15869 3834 15893 3836
rect 15949 3834 15973 3836
rect 16029 3834 16053 3836
rect 16109 3834 16115 3836
rect 15869 3782 15871 3834
rect 16051 3782 16053 3834
rect 15807 3780 15813 3782
rect 15869 3780 15893 3782
rect 15949 3780 15973 3782
rect 16029 3780 16053 3782
rect 16109 3780 16115 3782
rect 15807 3771 16115 3780
rect 16224 3670 16252 4270
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16132 3398 16160 3538
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 13556 400 13584 2230
rect 14200 400 14228 2774
rect 14844 400 14872 2774
rect 15488 2746 15608 2774
rect 15807 2748 16115 2757
rect 15807 2746 15813 2748
rect 15869 2746 15893 2748
rect 15949 2746 15973 2748
rect 16029 2746 16053 2748
rect 16109 2746 16115 2748
rect 15488 400 15516 2746
rect 15869 2694 15871 2746
rect 16051 2694 16053 2746
rect 15807 2692 15813 2694
rect 15869 2692 15893 2694
rect 15949 2692 15973 2694
rect 16029 2692 16053 2694
rect 16109 2692 16115 2694
rect 15807 2683 16115 2692
rect 15807 1660 16115 1669
rect 15807 1658 15813 1660
rect 15869 1658 15893 1660
rect 15949 1658 15973 1660
rect 16029 1658 16053 1660
rect 16109 1658 16115 1660
rect 15869 1606 15871 1658
rect 16051 1606 16053 1658
rect 15807 1604 15813 1606
rect 15869 1604 15893 1606
rect 15949 1604 15973 1606
rect 16029 1604 16053 1606
rect 16109 1604 16115 1606
rect 15807 1595 16115 1604
rect 15807 572 16115 581
rect 15807 570 15813 572
rect 15869 570 15893 572
rect 15949 570 15973 572
rect 16029 570 16053 572
rect 16109 570 16115 572
rect 15869 518 15871 570
rect 16051 518 16053 570
rect 15807 516 15813 518
rect 15869 516 15893 518
rect 15949 516 15973 518
rect 16029 516 16053 518
rect 16109 516 16115 518
rect 15807 507 16115 516
rect 16316 474 16344 5510
rect 16868 5234 16896 6190
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16408 4486 16436 4966
rect 16500 4826 16528 4966
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16684 4758 16712 4966
rect 16776 4826 16804 4966
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16868 4690 16896 5170
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16408 3738 16436 3946
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16500 3602 16528 4626
rect 16868 3602 16896 4626
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16960 2774 16988 8588
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17144 7342 17172 8298
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17328 5166 17356 5510
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17052 3670 17080 3878
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 17512 2774 17540 8230
rect 17604 8090 17632 9590
rect 17788 9110 17816 11018
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18064 10606 18092 10950
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 17960 9648 18012 9654
rect 17958 9616 17960 9625
rect 18012 9616 18014 9625
rect 17868 9580 17920 9586
rect 17958 9551 18014 9560
rect 17868 9522 17920 9528
rect 17776 9104 17828 9110
rect 17774 9072 17776 9081
rect 17828 9072 17830 9081
rect 17774 9007 17830 9016
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17604 6934 17632 8026
rect 17880 7562 17908 9522
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 9178 18092 9454
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 18156 9042 18184 10406
rect 18616 10130 18644 10950
rect 18708 10266 18736 19600
rect 19352 17105 19380 19600
rect 19660 18524 19968 18533
rect 19660 18522 19666 18524
rect 19722 18522 19746 18524
rect 19802 18522 19826 18524
rect 19882 18522 19906 18524
rect 19962 18522 19968 18524
rect 19722 18470 19724 18522
rect 19904 18470 19906 18522
rect 19660 18468 19666 18470
rect 19722 18468 19746 18470
rect 19802 18468 19826 18470
rect 19882 18468 19906 18470
rect 19962 18468 19968 18470
rect 19660 18459 19968 18468
rect 19660 17436 19968 17445
rect 19660 17434 19666 17436
rect 19722 17434 19746 17436
rect 19802 17434 19826 17436
rect 19882 17434 19906 17436
rect 19962 17434 19968 17436
rect 19722 17382 19724 17434
rect 19904 17382 19906 17434
rect 19660 17380 19666 17382
rect 19722 17380 19746 17382
rect 19802 17380 19826 17382
rect 19882 17380 19906 17382
rect 19962 17380 19968 17382
rect 19660 17371 19968 17380
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19338 17096 19394 17105
rect 19338 17031 19394 17040
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19260 16658 19288 16934
rect 19536 16658 19564 17138
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18800 14346 18828 16050
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19076 15706 19104 15846
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 18984 15552 19012 15642
rect 19064 15564 19116 15570
rect 18984 15524 19064 15552
rect 19168 15552 19196 15846
rect 19116 15524 19288 15552
rect 19064 15506 19116 15512
rect 18880 15496 18932 15502
rect 18932 15444 19196 15450
rect 18880 15438 19196 15444
rect 18892 15422 19196 15438
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 19076 14618 19104 15302
rect 19168 14618 19196 15422
rect 19260 15314 19288 15524
rect 19352 15434 19380 16594
rect 19996 16538 20024 19600
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20364 16969 20392 17070
rect 20444 17060 20496 17066
rect 20444 17002 20496 17008
rect 20350 16960 20406 16969
rect 20350 16895 20406 16904
rect 20350 16824 20406 16833
rect 20350 16759 20406 16768
rect 20260 16720 20312 16726
rect 20260 16662 20312 16668
rect 19996 16510 20208 16538
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19444 16130 19472 16390
rect 19536 16250 19564 16390
rect 19660 16348 19968 16357
rect 19660 16346 19666 16348
rect 19722 16346 19746 16348
rect 19802 16346 19826 16348
rect 19882 16346 19906 16348
rect 19962 16346 19968 16348
rect 19722 16294 19724 16346
rect 19904 16294 19906 16346
rect 19660 16292 19666 16294
rect 19722 16292 19746 16294
rect 19802 16292 19826 16294
rect 19882 16292 19906 16294
rect 19962 16292 19968 16294
rect 19660 16283 19968 16292
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19800 16176 19852 16182
rect 19444 16114 19656 16130
rect 19800 16118 19852 16124
rect 19444 16108 19668 16114
rect 19444 16102 19616 16108
rect 19616 16050 19668 16056
rect 19432 16040 19484 16046
rect 19484 16000 19564 16028
rect 19432 15982 19484 15988
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19444 15570 19472 15846
rect 19536 15706 19564 16000
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19812 15638 19840 16118
rect 19996 16046 20024 16390
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 20088 15638 20116 16390
rect 19800 15632 19852 15638
rect 19800 15574 19852 15580
rect 20076 15632 20128 15638
rect 20076 15574 20128 15580
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19432 15360 19484 15366
rect 19260 15286 19380 15314
rect 19432 15302 19484 15308
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19352 15162 19380 15286
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19444 14482 19472 15302
rect 19536 14482 19564 15302
rect 19660 15260 19968 15269
rect 19660 15258 19666 15260
rect 19722 15258 19746 15260
rect 19802 15258 19826 15260
rect 19882 15258 19906 15260
rect 19962 15258 19968 15260
rect 19722 15206 19724 15258
rect 19904 15206 19906 15258
rect 19660 15204 19666 15206
rect 19722 15204 19746 15206
rect 19802 15204 19826 15206
rect 19882 15204 19906 15206
rect 19962 15204 19968 15206
rect 19660 15195 19968 15204
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 18788 14340 18840 14346
rect 18788 14282 18840 14288
rect 18800 13938 18828 14282
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 14074 19288 14214
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19536 14006 19564 14418
rect 19660 14172 19968 14181
rect 19660 14170 19666 14172
rect 19722 14170 19746 14172
rect 19802 14170 19826 14172
rect 19882 14170 19906 14172
rect 19962 14170 19968 14172
rect 19722 14118 19724 14170
rect 19904 14118 19906 14170
rect 19660 14116 19666 14118
rect 19722 14116 19746 14118
rect 19802 14116 19826 14118
rect 19882 14116 19906 14118
rect 19962 14116 19968 14118
rect 19660 14107 19968 14116
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 19340 13728 19392 13734
rect 19062 13696 19118 13705
rect 19340 13670 19392 13676
rect 19062 13631 19118 13640
rect 19076 13530 19104 13631
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19352 12186 19380 13670
rect 19660 13084 19968 13093
rect 19660 13082 19666 13084
rect 19722 13082 19746 13084
rect 19802 13082 19826 13084
rect 19882 13082 19906 13084
rect 19962 13082 19968 13084
rect 19722 13030 19724 13082
rect 19904 13030 19906 13082
rect 19660 13028 19666 13030
rect 19722 13028 19746 13030
rect 19802 13028 19826 13030
rect 19882 13028 19906 13030
rect 19962 13028 19968 13030
rect 19660 13019 19968 13028
rect 20180 12986 20208 16510
rect 20272 16250 20300 16662
rect 20364 16590 20392 16759
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20456 16289 20484 17002
rect 20536 16448 20588 16454
rect 20536 16390 20588 16396
rect 20442 16280 20498 16289
rect 20260 16244 20312 16250
rect 20442 16215 20498 16224
rect 20260 16186 20312 16192
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20272 14958 20300 15846
rect 20364 15366 20392 15982
rect 20548 15706 20576 16390
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20640 15586 20668 19600
rect 20732 15688 20760 19638
rect 21192 19530 21220 19638
rect 21270 19600 21326 20000
rect 21914 19600 21970 20000
rect 22558 19600 22614 20000
rect 23202 19600 23258 20000
rect 23846 19600 23902 20000
rect 24490 19600 24546 20000
rect 25134 19600 25190 20000
rect 25240 19638 25452 19666
rect 21284 19530 21312 19600
rect 21192 19502 21312 19530
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 21008 17134 21036 17546
rect 21180 17536 21232 17542
rect 21928 17490 21956 19600
rect 21180 17478 21232 17484
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20824 16250 20852 16934
rect 21100 16726 21128 17002
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 20916 16250 20944 16662
rect 21192 16561 21220 17478
rect 21744 17462 21956 17490
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21284 16726 21312 17274
rect 21456 17128 21508 17134
rect 21640 17128 21692 17134
rect 21456 17070 21508 17076
rect 21546 17096 21602 17105
rect 21468 16794 21496 17070
rect 21640 17070 21692 17076
rect 21744 17082 21772 17462
rect 21836 17338 22232 17354
rect 21824 17332 22232 17338
rect 21876 17326 22232 17332
rect 21824 17274 21876 17280
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 22008 17128 22060 17134
rect 21546 17031 21602 17040
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21272 16720 21324 16726
rect 21272 16662 21324 16668
rect 21272 16584 21324 16590
rect 21178 16552 21234 16561
rect 21272 16526 21324 16532
rect 21178 16487 21234 16496
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 21192 16046 21220 16390
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 20732 15660 20852 15688
rect 20548 15558 20668 15586
rect 20720 15564 20772 15570
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20364 15094 20392 15302
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 20364 14770 20392 15030
rect 20272 14742 20392 14770
rect 20272 13802 20300 14742
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20364 13462 20392 14214
rect 20456 13841 20484 14214
rect 20442 13832 20498 13841
rect 20442 13767 20498 13776
rect 20548 13530 20576 15558
rect 20720 15506 20772 15512
rect 20732 14550 20760 15506
rect 20824 15162 20852 15660
rect 20916 15337 20944 15982
rect 21284 15910 21312 16526
rect 21376 16250 21404 16730
rect 21456 16652 21508 16658
rect 21560 16640 21588 17031
rect 21652 16998 21680 17070
rect 21744 17054 21864 17082
rect 22008 17070 22060 17076
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21730 16960 21786 16969
rect 21508 16612 21588 16640
rect 21456 16594 21508 16600
rect 21454 16552 21510 16561
rect 21454 16487 21510 16496
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21272 15904 21324 15910
rect 21376 15881 21404 15982
rect 21272 15846 21324 15852
rect 21362 15872 21418 15881
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 20902 15328 20958 15337
rect 20902 15263 20958 15272
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20720 14340 20772 14346
rect 20720 14282 20772 14288
rect 20732 14074 20760 14282
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 21008 13870 21036 15370
rect 21100 14618 21128 15846
rect 21284 15570 21312 15846
rect 21362 15807 21418 15816
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21192 14822 21220 15302
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20352 13456 20404 13462
rect 20352 13398 20404 13404
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20732 12782 20760 13126
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20824 12434 20852 12650
rect 20732 12406 20852 12434
rect 20732 12306 20760 12406
rect 20916 12306 20944 13126
rect 21100 12850 21128 13262
rect 21192 13161 21220 14214
rect 21284 13326 21312 15506
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21178 13152 21234 13161
rect 21178 13087 21234 13096
rect 21376 12918 21404 15302
rect 21468 15201 21496 16487
rect 21548 15904 21600 15910
rect 21652 15881 21680 16934
rect 21730 16895 21786 16904
rect 21744 16658 21772 16895
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21836 15994 21864 17054
rect 21916 16992 21968 16998
rect 22020 16969 22048 17070
rect 21916 16934 21968 16940
rect 22006 16960 22062 16969
rect 21744 15966 21864 15994
rect 21548 15846 21600 15852
rect 21638 15872 21694 15881
rect 21454 15192 21510 15201
rect 21454 15127 21510 15136
rect 21560 14657 21588 15846
rect 21638 15807 21694 15816
rect 21640 15360 21692 15366
rect 21640 15302 21692 15308
rect 21546 14648 21602 14657
rect 21546 14583 21602 14592
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 21468 13938 21496 14214
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21456 13796 21508 13802
rect 21456 13738 21508 13744
rect 21468 13394 21496 13738
rect 21560 13530 21588 14418
rect 21652 13977 21680 15302
rect 21744 14890 21772 15966
rect 21928 15910 21956 16934
rect 22006 16895 22062 16904
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 22020 15858 22048 16594
rect 22112 16250 22140 17206
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22204 16046 22232 17326
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22296 16658 22324 17206
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22282 16280 22338 16289
rect 22282 16215 22338 16224
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 21836 15745 21864 15846
rect 22020 15830 22140 15858
rect 21822 15736 21878 15745
rect 22112 15706 22140 15830
rect 22296 15706 22324 16215
rect 22388 16153 22416 17070
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22480 16250 22508 16390
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 22374 16144 22430 16153
rect 22374 16079 22376 16088
rect 22428 16079 22430 16088
rect 22376 16050 22428 16056
rect 22468 16040 22520 16046
rect 22572 16017 22600 19600
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22664 16794 22692 16934
rect 22756 16794 22784 17138
rect 23020 16992 23072 16998
rect 22834 16960 22890 16969
rect 23020 16934 23072 16940
rect 22834 16895 22890 16904
rect 22848 16794 22876 16895
rect 22926 16824 22982 16833
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22836 16788 22888 16794
rect 22926 16759 22982 16768
rect 22836 16730 22888 16736
rect 22744 16584 22796 16590
rect 22744 16526 22796 16532
rect 22756 16402 22784 16526
rect 22834 16416 22890 16425
rect 22756 16374 22834 16402
rect 22834 16351 22890 16360
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22468 15982 22520 15988
rect 22558 16008 22614 16017
rect 21822 15671 21878 15680
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 21914 15600 21970 15609
rect 21914 15535 21916 15544
rect 21968 15535 21970 15544
rect 22008 15564 22060 15570
rect 21916 15506 21968 15512
rect 22008 15506 22060 15512
rect 21732 14884 21784 14890
rect 21732 14826 21784 14832
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21744 14346 21772 14554
rect 21824 14476 21876 14482
rect 21876 14436 21956 14464
rect 21824 14418 21876 14424
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 21638 13968 21694 13977
rect 21638 13903 21694 13912
rect 21732 13864 21784 13870
rect 21652 13824 21732 13852
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21364 12912 21416 12918
rect 21364 12854 21416 12860
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 19536 12186 19564 12242
rect 18880 12164 18932 12170
rect 19352 12158 19564 12186
rect 18880 12106 18932 12112
rect 18892 11762 18920 12106
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 20076 12096 20128 12102
rect 20536 12096 20588 12102
rect 20076 12038 20128 12044
rect 20350 12064 20406 12073
rect 19338 11792 19394 11801
rect 18880 11756 18932 11762
rect 19338 11727 19394 11736
rect 18880 11698 18932 11704
rect 19352 11200 19380 11727
rect 19430 11656 19486 11665
rect 19430 11591 19486 11600
rect 19444 11354 19472 11591
rect 19536 11354 19564 12038
rect 19660 11996 19968 12005
rect 19660 11994 19666 11996
rect 19722 11994 19746 11996
rect 19802 11994 19826 11996
rect 19882 11994 19906 11996
rect 19962 11994 19968 11996
rect 19722 11942 19724 11994
rect 19904 11942 19906 11994
rect 19660 11940 19666 11942
rect 19722 11940 19746 11942
rect 19802 11940 19826 11942
rect 19882 11940 19906 11942
rect 19962 11940 19968 11942
rect 19660 11931 19968 11940
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19720 11354 19748 11630
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19996 11218 20024 11494
rect 20088 11354 20116 12038
rect 20536 12038 20588 12044
rect 20350 11999 20406 12008
rect 20364 11898 20392 11999
rect 20548 11898 20576 12038
rect 20640 11898 20668 12242
rect 20904 12164 20956 12170
rect 20904 12106 20956 12112
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20916 11676 20944 12106
rect 21008 11778 21036 12718
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 21100 11898 21128 12582
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21272 11824 21324 11830
rect 21008 11772 21272 11778
rect 21008 11766 21324 11772
rect 21008 11750 21312 11766
rect 20996 11688 21048 11694
rect 20916 11648 20996 11676
rect 20996 11630 21048 11636
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 21008 11286 21036 11630
rect 20996 11280 21048 11286
rect 20996 11222 21048 11228
rect 19984 11212 20036 11218
rect 19352 11172 19472 11200
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18892 10606 18920 10950
rect 19352 10810 19380 11018
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19444 10742 19472 11172
rect 19984 11154 20036 11160
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 19660 10908 19968 10917
rect 19660 10906 19666 10908
rect 19722 10906 19746 10908
rect 19802 10906 19826 10908
rect 19882 10906 19906 10908
rect 19962 10906 19968 10908
rect 19722 10854 19724 10906
rect 19904 10854 19906 10906
rect 19660 10852 19666 10854
rect 19722 10852 19746 10854
rect 19802 10852 19826 10854
rect 19882 10852 19906 10854
rect 19962 10852 19968 10854
rect 19660 10843 19968 10852
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 20272 10606 20300 11154
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20732 10606 20760 11086
rect 21180 11008 21232 11014
rect 21180 10950 21232 10956
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 10266 19932 10406
rect 20364 10266 20392 10542
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20916 10198 20944 10746
rect 21192 10606 21220 10950
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21376 10538 21404 12718
rect 21468 11082 21496 13126
rect 21560 12782 21588 13466
rect 21652 13138 21680 13824
rect 21732 13806 21784 13812
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21744 13394 21772 13670
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 21652 13110 21772 13138
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 21560 12306 21588 12718
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21652 12442 21680 12582
rect 21744 12442 21772 13110
rect 21836 12782 21864 13262
rect 21928 13258 21956 14436
rect 22020 14385 22048 15506
rect 22112 15366 22140 15642
rect 22480 15638 22508 15982
rect 22558 15943 22614 15952
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 22190 15464 22246 15473
rect 22190 15399 22192 15408
rect 22244 15399 22246 15408
rect 22192 15370 22244 15376
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 22112 14618 22140 15302
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 22100 14408 22152 14414
rect 22006 14376 22062 14385
rect 22100 14350 22152 14356
rect 22006 14311 22062 14320
rect 22112 13734 22140 14350
rect 22204 13870 22232 15098
rect 22296 13870 22324 15506
rect 22388 14278 22416 15506
rect 22480 14521 22508 15574
rect 22572 15162 22600 15846
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22756 14929 22784 16050
rect 22848 16046 22876 16351
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 22836 15904 22888 15910
rect 22836 15846 22888 15852
rect 22742 14920 22798 14929
rect 22742 14855 22798 14864
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22466 14512 22522 14521
rect 22466 14447 22522 14456
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22008 13728 22060 13734
rect 22008 13670 22060 13676
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22020 13530 22048 13670
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 22204 13326 22232 13806
rect 22572 13462 22600 14554
rect 22560 13456 22612 13462
rect 22560 13398 22612 13404
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 21916 13252 21968 13258
rect 21916 13194 21968 13200
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21560 11694 21588 12242
rect 21548 11688 21600 11694
rect 21548 11630 21600 11636
rect 21640 11688 21692 11694
rect 21744 11676 21772 12378
rect 21836 11694 21864 12718
rect 22204 12102 22232 13262
rect 22664 12850 22692 14758
rect 22848 14618 22876 15846
rect 22940 15706 22968 16759
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 23032 14890 23060 16934
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23020 14884 23072 14890
rect 23020 14826 23072 14832
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 23124 14550 23152 16730
rect 23216 15094 23244 19600
rect 23512 19068 23820 19077
rect 23512 19066 23518 19068
rect 23574 19066 23598 19068
rect 23654 19066 23678 19068
rect 23734 19066 23758 19068
rect 23814 19066 23820 19068
rect 23574 19014 23576 19066
rect 23756 19014 23758 19066
rect 23512 19012 23518 19014
rect 23574 19012 23598 19014
rect 23654 19012 23678 19014
rect 23734 19012 23758 19014
rect 23814 19012 23820 19014
rect 23512 19003 23820 19012
rect 23512 17980 23820 17989
rect 23512 17978 23518 17980
rect 23574 17978 23598 17980
rect 23654 17978 23678 17980
rect 23734 17978 23758 17980
rect 23814 17978 23820 17980
rect 23574 17926 23576 17978
rect 23756 17926 23758 17978
rect 23512 17924 23518 17926
rect 23574 17924 23598 17926
rect 23654 17924 23678 17926
rect 23734 17924 23758 17926
rect 23814 17924 23820 17926
rect 23512 17915 23820 17924
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 23308 16726 23336 17274
rect 23512 16892 23820 16901
rect 23512 16890 23518 16892
rect 23574 16890 23598 16892
rect 23654 16890 23678 16892
rect 23734 16890 23758 16892
rect 23814 16890 23820 16892
rect 23574 16838 23576 16890
rect 23756 16838 23758 16890
rect 23512 16836 23518 16838
rect 23574 16836 23598 16838
rect 23654 16836 23678 16838
rect 23734 16836 23758 16838
rect 23814 16836 23820 16838
rect 23512 16827 23820 16836
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23294 16280 23350 16289
rect 23294 16215 23296 16224
rect 23348 16215 23350 16224
rect 23296 16186 23348 16192
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23296 16040 23348 16046
rect 23296 15982 23348 15988
rect 23308 15706 23336 15982
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 23204 15088 23256 15094
rect 23204 15030 23256 15036
rect 23202 14648 23258 14657
rect 23202 14583 23258 14592
rect 23112 14544 23164 14550
rect 23112 14486 23164 14492
rect 23216 13530 23244 14583
rect 23308 14113 23336 15438
rect 23400 14958 23428 16118
rect 23584 16046 23612 16390
rect 23676 16250 23704 16594
rect 23756 16584 23808 16590
rect 23756 16526 23808 16532
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 23662 16008 23718 16017
rect 23768 15994 23796 16526
rect 23860 16017 23888 19600
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 23718 15966 23796 15994
rect 23662 15943 23718 15952
rect 23768 15892 23796 15966
rect 23846 16008 23902 16017
rect 23846 15943 23902 15952
rect 23768 15864 23888 15892
rect 23512 15804 23820 15813
rect 23512 15802 23518 15804
rect 23574 15802 23598 15804
rect 23654 15802 23678 15804
rect 23734 15802 23758 15804
rect 23814 15802 23820 15804
rect 23574 15750 23576 15802
rect 23756 15750 23758 15802
rect 23512 15748 23518 15750
rect 23574 15748 23598 15750
rect 23654 15748 23678 15750
rect 23734 15748 23758 15750
rect 23814 15748 23820 15750
rect 23512 15739 23820 15748
rect 23860 15688 23888 15864
rect 23768 15660 23888 15688
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23492 15026 23520 15302
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23768 14958 23796 15660
rect 23848 15496 23900 15502
rect 23846 15464 23848 15473
rect 23900 15464 23902 15473
rect 23846 15399 23902 15408
rect 23846 15328 23902 15337
rect 23846 15263 23902 15272
rect 23388 14952 23440 14958
rect 23388 14894 23440 14900
rect 23756 14952 23808 14958
rect 23756 14894 23808 14900
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23400 14498 23428 14758
rect 23512 14716 23820 14725
rect 23512 14714 23518 14716
rect 23574 14714 23598 14716
rect 23654 14714 23678 14716
rect 23734 14714 23758 14716
rect 23814 14714 23820 14716
rect 23574 14662 23576 14714
rect 23756 14662 23758 14714
rect 23512 14660 23518 14662
rect 23574 14660 23598 14662
rect 23654 14660 23678 14662
rect 23734 14660 23758 14662
rect 23814 14660 23820 14662
rect 23512 14651 23820 14660
rect 23400 14470 23520 14498
rect 23294 14104 23350 14113
rect 23294 14039 23350 14048
rect 23492 14006 23520 14470
rect 23860 14074 23888 15263
rect 23952 15162 23980 17206
rect 24214 17096 24270 17105
rect 24270 17054 24440 17082
rect 24214 17031 24270 17040
rect 24308 16516 24360 16522
rect 24308 16458 24360 16464
rect 24320 16182 24348 16458
rect 24308 16176 24360 16182
rect 24030 16144 24086 16153
rect 24308 16118 24360 16124
rect 24086 16088 24256 16096
rect 24030 16079 24032 16088
rect 24084 16068 24256 16088
rect 24032 16050 24084 16056
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 24136 15638 24164 15846
rect 24032 15632 24084 15638
rect 24032 15574 24084 15580
rect 24124 15632 24176 15638
rect 24124 15574 24176 15580
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 24044 14618 24072 15574
rect 24228 15570 24256 16068
rect 24320 16046 24348 16118
rect 24308 16040 24360 16046
rect 24308 15982 24360 15988
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 24228 15366 24256 15506
rect 24320 15473 24348 15982
rect 24306 15464 24362 15473
rect 24306 15399 24362 15408
rect 24216 15360 24268 15366
rect 24136 15320 24216 15348
rect 24136 14958 24164 15320
rect 24216 15302 24268 15308
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 24136 14482 24164 14554
rect 23940 14476 23992 14482
rect 24124 14476 24176 14482
rect 23992 14436 24072 14464
rect 23940 14418 23992 14424
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23480 14000 23532 14006
rect 23480 13942 23532 13948
rect 23768 13954 23796 14010
rect 23768 13926 23980 13954
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 23846 13832 23902 13841
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23308 13297 23336 13806
rect 23846 13767 23902 13776
rect 23512 13628 23820 13637
rect 23512 13626 23518 13628
rect 23574 13626 23598 13628
rect 23654 13626 23678 13628
rect 23734 13626 23758 13628
rect 23814 13626 23820 13628
rect 23574 13574 23576 13626
rect 23756 13574 23758 13626
rect 23512 13572 23518 13574
rect 23574 13572 23598 13574
rect 23654 13572 23678 13574
rect 23734 13572 23758 13574
rect 23814 13572 23820 13574
rect 23512 13563 23820 13572
rect 23664 13388 23716 13394
rect 23664 13330 23716 13336
rect 23294 13288 23350 13297
rect 23294 13223 23350 13232
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 23676 12753 23704 13330
rect 23860 12782 23888 13767
rect 23952 12782 23980 13926
rect 24044 12782 24072 14436
rect 24124 14418 24176 14424
rect 24228 14278 24256 15098
rect 24320 14618 24348 15399
rect 24412 14822 24440 17054
rect 24504 16538 24532 19600
rect 25148 19530 25176 19600
rect 25240 19530 25268 19638
rect 25148 19502 25268 19530
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24504 16510 24716 16538
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 24596 15570 24624 16390
rect 24584 15564 24636 15570
rect 24504 15524 24584 15552
rect 24504 14958 24532 15524
rect 24584 15506 24636 15512
rect 24688 15314 24716 16510
rect 24858 16416 24914 16425
rect 24858 16351 24914 16360
rect 24872 15570 24900 16351
rect 24964 15706 24992 17070
rect 25136 17060 25188 17066
rect 25136 17002 25188 17008
rect 25042 16280 25098 16289
rect 25042 16215 25098 16224
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24596 15286 24716 15314
rect 24596 15065 24624 15286
rect 24674 15192 24730 15201
rect 24674 15127 24730 15136
rect 24582 15056 24638 15065
rect 24582 14991 24638 15000
rect 24688 14958 24716 15127
rect 25056 15094 25084 16215
rect 25148 15094 25176 17002
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25044 15088 25096 15094
rect 25044 15030 25096 15036
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 25240 14958 25268 16050
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 24492 14952 24544 14958
rect 24492 14894 24544 14900
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24676 14952 24728 14958
rect 24768 14952 24820 14958
rect 24676 14894 24728 14900
rect 24766 14920 24768 14929
rect 25228 14952 25280 14958
rect 24820 14920 24822 14929
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24596 14618 24624 14894
rect 25228 14894 25280 14900
rect 24766 14855 24822 14864
rect 24952 14816 25004 14822
rect 24952 14758 25004 14764
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24584 14612 24636 14618
rect 24964 14600 24992 14758
rect 24584 14554 24636 14560
rect 24826 14572 24992 14600
rect 24400 14476 24452 14482
rect 24400 14418 24452 14424
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24412 13870 24440 14418
rect 24826 14414 24854 14572
rect 24952 14476 25004 14482
rect 25004 14436 25084 14464
rect 24952 14418 25004 14424
rect 24814 14408 24866 14414
rect 24490 14376 24546 14385
rect 24814 14350 24866 14356
rect 24490 14311 24546 14320
rect 24952 14340 25004 14346
rect 24504 13870 24532 14311
rect 24952 14282 25004 14288
rect 24584 14272 24636 14278
rect 24964 14249 24992 14282
rect 24584 14214 24636 14220
rect 24950 14240 25006 14249
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24216 13796 24268 13802
rect 24216 13738 24268 13744
rect 24228 13462 24256 13738
rect 24490 13696 24546 13705
rect 24490 13631 24546 13640
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 24504 13394 24532 13631
rect 24596 13569 24624 14214
rect 24950 14175 25006 14184
rect 24768 14000 24820 14006
rect 24674 13968 24730 13977
rect 24768 13942 24820 13948
rect 25056 13954 25084 14436
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 25148 14074 25176 14214
rect 25332 14074 25360 15370
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25228 14000 25280 14006
rect 25056 13948 25228 13954
rect 25056 13942 25280 13948
rect 24674 13903 24730 13912
rect 24582 13560 24638 13569
rect 24582 13495 24638 13504
rect 24584 13456 24636 13462
rect 24584 13398 24636 13404
rect 24492 13388 24544 13394
rect 24492 13330 24544 13336
rect 24490 13152 24546 13161
rect 24490 13087 24546 13096
rect 24504 12986 24532 13087
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 23848 12776 23900 12782
rect 23662 12744 23718 12753
rect 23848 12718 23900 12724
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 24308 12776 24360 12782
rect 24360 12736 24440 12764
rect 24308 12718 24360 12724
rect 23662 12679 23718 12688
rect 24412 12646 24440 12736
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22204 11694 22232 12038
rect 21692 11648 21772 11676
rect 21824 11688 21876 11694
rect 21640 11630 21692 11636
rect 21824 11630 21876 11636
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21560 11218 21588 11494
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21560 10606 21588 11018
rect 21652 11014 21680 11630
rect 21732 11280 21784 11286
rect 21836 11268 21864 11630
rect 21784 11240 21864 11268
rect 21732 11222 21784 11228
rect 22204 11218 22232 11630
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 21640 11008 21692 11014
rect 21640 10950 21692 10956
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 22100 10600 22152 10606
rect 22204 10588 22232 11154
rect 22152 10560 22232 10588
rect 22100 10542 22152 10548
rect 21364 10532 21416 10538
rect 21364 10474 21416 10480
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21284 10198 21312 10406
rect 20904 10192 20956 10198
rect 20904 10134 20956 10140
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 21928 10130 21956 10474
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 21364 10124 21416 10130
rect 21732 10124 21784 10130
rect 21364 10066 21416 10072
rect 21652 10084 21732 10112
rect 21376 9926 21404 10066
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 19660 9820 19968 9829
rect 19660 9818 19666 9820
rect 19722 9818 19746 9820
rect 19802 9818 19826 9820
rect 19882 9818 19906 9820
rect 19962 9818 19968 9820
rect 19722 9766 19724 9818
rect 19904 9766 19906 9818
rect 19660 9764 19666 9766
rect 19722 9764 19746 9766
rect 19802 9764 19826 9766
rect 19882 9764 19906 9766
rect 19962 9764 19968 9766
rect 19660 9755 19968 9764
rect 20180 9722 20208 9862
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 21362 9616 21418 9625
rect 21362 9551 21418 9560
rect 21376 9518 21404 9551
rect 21652 9518 21680 10084
rect 21732 10066 21784 10072
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 22112 9994 22140 10542
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 21928 9518 21956 9862
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21640 9512 21692 9518
rect 21640 9454 21692 9460
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18248 8634 18276 9454
rect 19338 9072 19394 9081
rect 19338 9007 19394 9016
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18340 8634 18368 8774
rect 18800 8634 18828 8910
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17972 7750 18000 8366
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18524 7954 18552 8298
rect 18788 8016 18840 8022
rect 18788 7958 18840 7964
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 17788 7546 17908 7562
rect 17776 7540 17908 7546
rect 17828 7534 17908 7540
rect 17776 7482 17828 7488
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17880 6798 17908 7534
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17880 5914 17908 6734
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 6322 18000 6598
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 16776 2746 16988 2774
rect 17420 2746 17540 2774
rect 16028 468 16080 474
rect 16304 468 16356 474
rect 16080 428 16160 456
rect 16028 410 16080 416
rect 16132 400 16160 428
rect 16304 410 16356 416
rect 16776 400 16804 2746
rect 17420 400 17448 2746
rect 18064 400 18092 6326
rect 18156 2774 18184 7686
rect 18800 7546 18828 7958
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18340 6390 18368 7142
rect 18432 7002 18460 7142
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 18328 6248 18380 6254
rect 18524 6236 18552 7142
rect 18616 6458 18644 7414
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18708 6866 18736 7278
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18800 6798 18828 7482
rect 18892 7342 18920 8434
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19064 7812 19116 7818
rect 19064 7754 19116 7760
rect 19076 7342 19104 7754
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 18972 7268 19024 7274
rect 18972 7210 19024 7216
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18892 6746 18920 6938
rect 18984 6848 19012 7210
rect 19168 7206 19196 8230
rect 19352 8022 19380 9007
rect 19444 8430 19472 9454
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 19660 8732 19968 8741
rect 19660 8730 19666 8732
rect 19722 8730 19746 8732
rect 19802 8730 19826 8732
rect 19882 8730 19906 8732
rect 19962 8730 19968 8732
rect 19722 8678 19724 8730
rect 19904 8678 19906 8730
rect 19660 8676 19666 8678
rect 19722 8676 19746 8678
rect 19802 8676 19826 8678
rect 19882 8676 19906 8678
rect 19962 8676 19968 8678
rect 19660 8667 19968 8676
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19444 7478 19472 8230
rect 19524 7812 19576 7818
rect 19524 7754 19576 7760
rect 19432 7472 19484 7478
rect 19432 7414 19484 7420
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 18984 6820 19104 6848
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18708 6322 18736 6598
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18380 6208 18552 6236
rect 18328 6190 18380 6196
rect 18800 5914 18828 6734
rect 18892 6718 19012 6746
rect 18880 6248 18932 6254
rect 18878 6216 18880 6225
rect 18932 6216 18934 6225
rect 18878 6151 18934 6160
rect 18984 5930 19012 6718
rect 19076 6458 19104 6820
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19168 6390 19196 7142
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19352 6458 19380 6802
rect 19536 6746 19564 7754
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19660 7644 19968 7653
rect 19660 7642 19666 7644
rect 19722 7642 19746 7644
rect 19802 7642 19826 7644
rect 19882 7642 19906 7644
rect 19962 7642 19968 7644
rect 19722 7590 19724 7642
rect 19904 7590 19906 7642
rect 19660 7588 19666 7590
rect 19722 7588 19746 7590
rect 19802 7588 19826 7590
rect 19882 7588 19906 7590
rect 19962 7588 19968 7590
rect 19660 7579 19968 7588
rect 19800 7472 19852 7478
rect 19800 7414 19852 7420
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19444 6718 19564 6746
rect 19628 6730 19656 7346
rect 19706 7304 19762 7313
rect 19706 7239 19762 7248
rect 19720 6934 19748 7239
rect 19812 7206 19840 7414
rect 19800 7200 19852 7206
rect 19800 7142 19852 7148
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19904 7002 19932 7142
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 19708 6928 19760 6934
rect 19708 6870 19760 6876
rect 19616 6724 19668 6730
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19156 6384 19208 6390
rect 19156 6326 19208 6332
rect 19168 6254 19196 6326
rect 19156 6248 19208 6254
rect 19444 6236 19472 6718
rect 19616 6666 19668 6672
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19536 6458 19564 6598
rect 19660 6556 19968 6565
rect 19660 6554 19666 6556
rect 19722 6554 19746 6556
rect 19802 6554 19826 6556
rect 19882 6554 19906 6556
rect 19962 6554 19968 6556
rect 19722 6502 19724 6554
rect 19904 6502 19906 6554
rect 19660 6500 19666 6502
rect 19722 6500 19746 6502
rect 19802 6500 19826 6502
rect 19882 6500 19906 6502
rect 19962 6500 19968 6502
rect 19660 6491 19968 6500
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19260 6225 19472 6236
rect 19156 6190 19208 6196
rect 19246 6216 19472 6225
rect 19302 6208 19472 6216
rect 19246 6151 19302 6160
rect 19248 6112 19300 6118
rect 19996 6100 20024 7686
rect 20088 6338 20116 9318
rect 20260 8900 20312 8906
rect 20260 8842 20312 8848
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20180 8401 20208 8774
rect 20272 8430 20300 8842
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20364 8566 20392 8774
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20260 8424 20312 8430
rect 20166 8392 20222 8401
rect 20260 8366 20312 8372
rect 20536 8424 20588 8430
rect 20732 8378 20760 9318
rect 21100 9178 21128 9386
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 20996 9104 21048 9110
rect 21048 9052 21128 9058
rect 20996 9046 21128 9052
rect 21008 9030 21128 9046
rect 21284 9042 21312 9318
rect 21560 9178 21588 9318
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 20812 8968 20864 8974
rect 20864 8928 20944 8956
rect 20812 8910 20864 8916
rect 20916 8566 20944 8928
rect 20904 8560 20956 8566
rect 20904 8502 20956 8508
rect 20588 8372 20852 8378
rect 20536 8366 20852 8372
rect 20548 8350 20852 8366
rect 20166 8327 20222 8336
rect 20260 8288 20312 8294
rect 20260 8230 20312 8236
rect 20272 7886 20300 8230
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20168 7336 20220 7342
rect 20166 7304 20168 7313
rect 20272 7324 20300 7822
rect 20220 7304 20300 7324
rect 20222 7296 20300 7304
rect 20166 7239 20222 7248
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20180 7002 20208 7142
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20088 6310 20208 6338
rect 20076 6180 20128 6186
rect 20076 6122 20128 6128
rect 19300 6072 20024 6100
rect 19248 6054 19300 6060
rect 20088 5953 20116 6122
rect 20074 5944 20130 5953
rect 18788 5908 18840 5914
rect 18984 5902 19472 5930
rect 18788 5850 18840 5856
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19062 5672 19118 5681
rect 19062 5607 19064 5616
rect 19116 5607 19118 5616
rect 19064 5578 19116 5584
rect 19168 5166 19196 5714
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19260 5370 19288 5578
rect 19352 5370 19380 5714
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18340 4282 18368 4422
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18156 2746 18368 2774
rect 8298 368 8354 377
rect 8298 303 8354 312
rect 8390 0 8446 400
rect 9034 0 9090 400
rect 9678 0 9734 400
rect 10322 0 10378 400
rect 10966 0 11022 400
rect 11610 0 11666 400
rect 12254 0 12310 400
rect 12898 0 12954 400
rect 13542 0 13598 400
rect 14186 0 14242 400
rect 14830 0 14886 400
rect 15474 0 15530 400
rect 16118 0 16174 400
rect 16762 0 16818 400
rect 17406 0 17462 400
rect 18050 0 18106 400
rect 18340 354 18368 2746
rect 18616 462 18736 490
rect 18616 354 18644 462
rect 18708 400 18736 462
rect 19352 400 19380 4558
rect 19444 2774 19472 5902
rect 20074 5879 20130 5888
rect 20076 5704 20128 5710
rect 19996 5664 20076 5692
rect 19660 5468 19968 5477
rect 19660 5466 19666 5468
rect 19722 5466 19746 5468
rect 19802 5466 19826 5468
rect 19882 5466 19906 5468
rect 19962 5466 19968 5468
rect 19722 5414 19724 5466
rect 19904 5414 19906 5466
rect 19660 5412 19666 5414
rect 19722 5412 19746 5414
rect 19802 5412 19826 5414
rect 19882 5412 19906 5414
rect 19962 5412 19968 5414
rect 19660 5403 19968 5412
rect 19996 5166 20024 5664
rect 20076 5646 20128 5652
rect 19708 5160 19760 5166
rect 19984 5160 20036 5166
rect 19760 5120 19984 5148
rect 19708 5102 19760 5108
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19536 4214 19564 4966
rect 19904 4826 19932 5120
rect 19984 5102 20036 5108
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 20088 4826 20116 4966
rect 19892 4820 19944 4826
rect 19892 4762 19944 4768
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 20180 4622 20208 6310
rect 20272 5234 20300 6394
rect 20364 6186 20392 7142
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20352 6180 20404 6186
rect 20352 6122 20404 6128
rect 20456 5914 20484 6802
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20548 5914 20576 6734
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20350 5808 20406 5817
rect 20548 5794 20576 5850
rect 20732 5846 20760 6598
rect 20824 6390 20852 8350
rect 21100 8276 21128 9030
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 21652 8906 21680 9454
rect 21744 9058 21772 9454
rect 22112 9450 22140 9930
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22204 9178 22232 9386
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22388 9110 22416 12582
rect 23512 12540 23820 12549
rect 23512 12538 23518 12540
rect 23574 12538 23598 12540
rect 23654 12538 23678 12540
rect 23734 12538 23758 12540
rect 23814 12538 23820 12540
rect 23574 12486 23576 12538
rect 23756 12486 23758 12538
rect 23512 12484 23518 12486
rect 23574 12484 23598 12486
rect 23654 12484 23678 12486
rect 23734 12484 23758 12486
rect 23814 12484 23820 12486
rect 23512 12475 23820 12484
rect 23294 11792 23350 11801
rect 23294 11727 23350 11736
rect 23308 11286 23336 11727
rect 24320 11694 24348 12582
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24308 11688 24360 11694
rect 24308 11630 24360 11636
rect 24032 11620 24084 11626
rect 24032 11562 24084 11568
rect 23512 11452 23820 11461
rect 23512 11450 23518 11452
rect 23574 11450 23598 11452
rect 23654 11450 23678 11452
rect 23734 11450 23758 11452
rect 23814 11450 23820 11452
rect 23574 11398 23576 11450
rect 23756 11398 23758 11450
rect 23512 11396 23518 11398
rect 23574 11396 23598 11398
rect 23654 11396 23678 11398
rect 23734 11396 23758 11398
rect 23814 11396 23820 11398
rect 23512 11387 23820 11396
rect 23296 11280 23348 11286
rect 23296 11222 23348 11228
rect 23848 11280 23900 11286
rect 24044 11268 24072 11562
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24216 11552 24268 11558
rect 24216 11494 24268 11500
rect 24136 11286 24164 11494
rect 24228 11354 24256 11494
rect 24412 11354 24440 12378
rect 24596 12306 24624 13398
rect 24688 12986 24716 13903
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24780 12764 24808 13942
rect 25056 13926 25268 13942
rect 24860 13864 24912 13870
rect 25424 13818 25452 19638
rect 31217 19068 31525 19077
rect 31217 19066 31223 19068
rect 31279 19066 31303 19068
rect 31359 19066 31383 19068
rect 31439 19066 31463 19068
rect 31519 19066 31525 19068
rect 31279 19014 31281 19066
rect 31461 19014 31463 19066
rect 31217 19012 31223 19014
rect 31279 19012 31303 19014
rect 31359 19012 31383 19014
rect 31439 19012 31463 19014
rect 31519 19012 31525 19014
rect 31217 19003 31525 19012
rect 27365 18524 27673 18533
rect 27365 18522 27371 18524
rect 27427 18522 27451 18524
rect 27507 18522 27531 18524
rect 27587 18522 27611 18524
rect 27667 18522 27673 18524
rect 27427 18470 27429 18522
rect 27609 18470 27611 18522
rect 27365 18468 27371 18470
rect 27427 18468 27451 18470
rect 27507 18468 27531 18470
rect 27587 18468 27611 18470
rect 27667 18468 27673 18470
rect 27365 18459 27673 18468
rect 31217 17980 31525 17989
rect 31217 17978 31223 17980
rect 31279 17978 31303 17980
rect 31359 17978 31383 17980
rect 31439 17978 31463 17980
rect 31519 17978 31525 17980
rect 31279 17926 31281 17978
rect 31461 17926 31463 17978
rect 31217 17924 31223 17926
rect 31279 17924 31303 17926
rect 31359 17924 31383 17926
rect 31439 17924 31463 17926
rect 31519 17924 31525 17926
rect 31217 17915 31525 17924
rect 27365 17436 27673 17445
rect 27365 17434 27371 17436
rect 27427 17434 27451 17436
rect 27507 17434 27531 17436
rect 27587 17434 27611 17436
rect 27667 17434 27673 17436
rect 27427 17382 27429 17434
rect 27609 17382 27611 17434
rect 27365 17380 27371 17382
rect 27427 17380 27451 17382
rect 27507 17380 27531 17382
rect 27587 17380 27611 17382
rect 27667 17380 27673 17382
rect 27365 17371 27673 17380
rect 31217 16892 31525 16901
rect 31217 16890 31223 16892
rect 31279 16890 31303 16892
rect 31359 16890 31383 16892
rect 31439 16890 31463 16892
rect 31519 16890 31525 16892
rect 31279 16838 31281 16890
rect 31461 16838 31463 16890
rect 31217 16836 31223 16838
rect 31279 16836 31303 16838
rect 31359 16836 31383 16838
rect 31439 16836 31463 16838
rect 31519 16836 31525 16838
rect 31217 16827 31525 16836
rect 27365 16348 27673 16357
rect 27365 16346 27371 16348
rect 27427 16346 27451 16348
rect 27507 16346 27531 16348
rect 27587 16346 27611 16348
rect 27667 16346 27673 16348
rect 27427 16294 27429 16346
rect 27609 16294 27611 16346
rect 27365 16292 27371 16294
rect 27427 16292 27451 16294
rect 27507 16292 27531 16294
rect 27587 16292 27611 16294
rect 27667 16292 27673 16294
rect 27365 16283 27673 16292
rect 26424 16040 26476 16046
rect 26424 15982 26476 15988
rect 25688 15632 25740 15638
rect 25688 15574 25740 15580
rect 25504 14816 25556 14822
rect 25556 14776 25636 14804
rect 25504 14758 25556 14764
rect 25502 14512 25558 14521
rect 25502 14447 25504 14456
rect 25556 14447 25558 14456
rect 25504 14418 25556 14424
rect 24860 13806 24912 13812
rect 24872 13394 24900 13806
rect 25240 13790 25452 13818
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24858 13152 24914 13161
rect 24858 13087 24914 13096
rect 24872 12918 24900 13087
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24952 12776 25004 12782
rect 24780 12736 24952 12764
rect 24952 12718 25004 12724
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24768 12300 24820 12306
rect 24768 12242 24820 12248
rect 24504 12102 24532 12242
rect 24676 12164 24728 12170
rect 24676 12106 24728 12112
rect 24492 12096 24544 12102
rect 24492 12038 24544 12044
rect 24688 11694 24716 12106
rect 24780 11898 24808 12242
rect 25240 12073 25268 13790
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 25516 13682 25544 14418
rect 25608 14074 25636 14776
rect 25700 14618 25728 15574
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 25872 14884 25924 14890
rect 25872 14826 25924 14832
rect 25780 14816 25832 14822
rect 25780 14758 25832 14764
rect 25792 14618 25820 14758
rect 25688 14612 25740 14618
rect 25688 14554 25740 14560
rect 25780 14612 25832 14618
rect 25780 14554 25832 14560
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25688 14408 25740 14414
rect 25688 14350 25740 14356
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25700 13977 25728 14350
rect 25686 13968 25742 13977
rect 25686 13903 25742 13912
rect 25596 13864 25648 13870
rect 25792 13852 25820 14418
rect 25884 13870 25912 14826
rect 26146 14240 26202 14249
rect 26146 14175 26202 14184
rect 25962 14104 26018 14113
rect 26160 14074 26188 14175
rect 25962 14039 26018 14048
rect 26148 14068 26200 14074
rect 25648 13824 25820 13852
rect 25596 13806 25648 13812
rect 25688 13728 25740 13734
rect 25424 13530 25452 13670
rect 25516 13654 25636 13682
rect 25688 13670 25740 13676
rect 25502 13560 25558 13569
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25412 13524 25464 13530
rect 25502 13495 25558 13504
rect 25412 13466 25464 13472
rect 25332 13433 25360 13466
rect 25318 13424 25374 13433
rect 25516 13394 25544 13495
rect 25318 13359 25374 13368
rect 25504 13388 25556 13394
rect 25504 13330 25556 13336
rect 25608 13002 25636 13654
rect 25700 13394 25728 13670
rect 25792 13462 25820 13824
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25780 13456 25832 13462
rect 25780 13398 25832 13404
rect 25688 13388 25740 13394
rect 25688 13330 25740 13336
rect 25608 12974 25820 13002
rect 25884 12986 25912 13806
rect 25976 13530 26004 14039
rect 26148 14010 26200 14016
rect 26344 13870 26372 15438
rect 26436 14074 26464 15982
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26620 13870 26648 15846
rect 31217 15804 31525 15813
rect 31217 15802 31223 15804
rect 31279 15802 31303 15804
rect 31359 15802 31383 15804
rect 31439 15802 31463 15804
rect 31519 15802 31525 15804
rect 31279 15750 31281 15802
rect 31461 15750 31463 15802
rect 31217 15748 31223 15750
rect 31279 15748 31303 15750
rect 31359 15748 31383 15750
rect 31439 15748 31463 15750
rect 31519 15748 31525 15750
rect 31217 15739 31525 15748
rect 31666 15736 31722 15745
rect 31666 15671 31722 15680
rect 27365 15260 27673 15269
rect 27365 15258 27371 15260
rect 27427 15258 27451 15260
rect 27507 15258 27531 15260
rect 27587 15258 27611 15260
rect 27667 15258 27673 15260
rect 27427 15206 27429 15258
rect 27609 15206 27611 15258
rect 27365 15204 27371 15206
rect 27427 15204 27451 15206
rect 27507 15204 27531 15206
rect 27587 15204 27611 15206
rect 27667 15204 27673 15206
rect 27365 15195 27673 15204
rect 28264 15156 28316 15162
rect 28264 15098 28316 15104
rect 28276 15065 28304 15098
rect 28262 15056 28318 15065
rect 28262 14991 28318 15000
rect 31680 14822 31708 15671
rect 28264 14816 28316 14822
rect 28264 14758 28316 14764
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 31668 14816 31720 14822
rect 31668 14758 31720 14764
rect 28276 14385 28304 14758
rect 28262 14376 28318 14385
rect 28262 14311 28318 14320
rect 27365 14172 27673 14181
rect 27365 14170 27371 14172
rect 27427 14170 27451 14172
rect 27507 14170 27531 14172
rect 27587 14170 27611 14172
rect 27667 14170 27673 14172
rect 27427 14118 27429 14170
rect 27609 14118 27611 14170
rect 27365 14116 27371 14118
rect 27427 14116 27451 14118
rect 27507 14116 27531 14118
rect 27587 14116 27611 14118
rect 27667 14116 27673 14118
rect 27365 14107 27673 14116
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26700 13728 26752 13734
rect 26700 13670 26752 13676
rect 25964 13524 26016 13530
rect 25964 13466 26016 13472
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 25594 12880 25650 12889
rect 25792 12850 25820 12974
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 25594 12815 25596 12824
rect 25648 12815 25650 12824
rect 25780 12844 25832 12850
rect 25596 12786 25648 12792
rect 25780 12786 25832 12792
rect 25596 12096 25648 12102
rect 25226 12064 25282 12073
rect 25596 12038 25648 12044
rect 25226 11999 25282 12008
rect 25608 11898 25636 12038
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25596 11892 25648 11898
rect 25596 11834 25648 11840
rect 24492 11688 24544 11694
rect 24490 11656 24492 11665
rect 24676 11688 24728 11694
rect 24544 11656 24546 11665
rect 24676 11630 24728 11636
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 25516 11642 25544 11834
rect 25976 11694 26004 13262
rect 26436 13190 26464 13466
rect 26712 13297 26740 13670
rect 26698 13288 26754 13297
rect 26698 13223 26754 13232
rect 26424 13184 26476 13190
rect 26424 13126 26476 13132
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 26332 12776 26384 12782
rect 26146 12744 26202 12753
rect 26056 12708 26108 12714
rect 26332 12718 26384 12724
rect 26146 12679 26202 12688
rect 26056 12650 26108 12656
rect 26068 12374 26096 12650
rect 26160 12374 26188 12679
rect 26056 12368 26108 12374
rect 26056 12310 26108 12316
rect 26148 12368 26200 12374
rect 26148 12310 26200 12316
rect 26344 12306 26372 12718
rect 26528 12374 26556 13126
rect 27365 13084 27673 13093
rect 27365 13082 27371 13084
rect 27427 13082 27451 13084
rect 27507 13082 27531 13084
rect 27587 13082 27611 13084
rect 27667 13082 27673 13084
rect 27427 13030 27429 13082
rect 27609 13030 27611 13082
rect 27365 13028 27371 13030
rect 27427 13028 27451 13030
rect 27507 13028 27531 13030
rect 27587 13028 27611 13030
rect 27667 13028 27673 13030
rect 27365 13019 27673 13028
rect 28276 13025 28304 13126
rect 28262 13016 28318 13025
rect 28262 12951 28318 12960
rect 28264 12436 28316 12442
rect 28264 12378 28316 12384
rect 26516 12368 26568 12374
rect 28276 12345 28304 12378
rect 26516 12310 26568 12316
rect 28262 12336 28318 12345
rect 26332 12300 26384 12306
rect 28262 12271 28318 12280
rect 26332 12242 26384 12248
rect 27365 11996 27673 12005
rect 27365 11994 27371 11996
rect 27427 11994 27451 11996
rect 27507 11994 27531 11996
rect 27587 11994 27611 11996
rect 27667 11994 27673 11996
rect 27427 11942 27429 11994
rect 27609 11942 27611 11994
rect 27365 11940 27371 11942
rect 27427 11940 27451 11942
rect 27507 11940 27531 11942
rect 27587 11940 27611 11942
rect 27667 11940 27673 11942
rect 27365 11931 27673 11940
rect 29656 11801 29684 14758
rect 31217 14716 31525 14725
rect 31217 14714 31223 14716
rect 31279 14714 31303 14716
rect 31359 14714 31383 14716
rect 31439 14714 31463 14716
rect 31519 14714 31525 14716
rect 31279 14662 31281 14714
rect 31461 14662 31463 14714
rect 31217 14660 31223 14662
rect 31279 14660 31303 14662
rect 31359 14660 31383 14662
rect 31439 14660 31463 14662
rect 31519 14660 31525 14662
rect 31217 14651 31525 14660
rect 31666 13696 31722 13705
rect 31217 13628 31525 13637
rect 31666 13631 31722 13640
rect 31217 13626 31223 13628
rect 31279 13626 31303 13628
rect 31359 13626 31383 13628
rect 31439 13626 31463 13628
rect 31519 13626 31525 13628
rect 31279 13574 31281 13626
rect 31461 13574 31463 13626
rect 31217 13572 31223 13574
rect 31279 13572 31303 13574
rect 31359 13572 31383 13574
rect 31439 13572 31463 13574
rect 31519 13572 31525 13574
rect 31217 13563 31525 13572
rect 31680 13530 31708 13631
rect 31668 13524 31720 13530
rect 31668 13466 31720 13472
rect 31217 12540 31525 12549
rect 31217 12538 31223 12540
rect 31279 12538 31303 12540
rect 31359 12538 31383 12540
rect 31439 12538 31463 12540
rect 31519 12538 31525 12540
rect 31279 12486 31281 12538
rect 31461 12486 31463 12538
rect 31217 12484 31223 12486
rect 31279 12484 31303 12486
rect 31359 12484 31383 12486
rect 31439 12484 31463 12486
rect 31519 12484 31525 12486
rect 31217 12475 31525 12484
rect 29642 11792 29698 11801
rect 29642 11727 29698 11736
rect 25964 11688 26016 11694
rect 25962 11656 25964 11665
rect 26016 11656 26018 11665
rect 24490 11591 24546 11600
rect 25056 11354 25084 11630
rect 25516 11626 25912 11642
rect 25516 11620 25924 11626
rect 25516 11614 25872 11620
rect 25962 11591 26018 11600
rect 28262 11656 28318 11665
rect 28262 11591 28318 11600
rect 25872 11562 25924 11568
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 25412 11552 25464 11558
rect 25412 11494 25464 11500
rect 24216 11348 24268 11354
rect 24216 11290 24268 11296
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 25044 11348 25096 11354
rect 25044 11290 25096 11296
rect 23900 11240 24072 11268
rect 24124 11280 24176 11286
rect 23848 11222 23900 11228
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23492 10606 23520 10950
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23584 10470 23612 11154
rect 23952 11082 23980 11240
rect 24124 11222 24176 11228
rect 24412 11234 24440 11290
rect 24412 11218 24532 11234
rect 24216 11212 24268 11218
rect 24412 11212 24544 11218
rect 24412 11206 24492 11212
rect 24216 11154 24268 11160
rect 24492 11154 24544 11160
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 24228 11098 24256 11154
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 24228 11070 24532 11098
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23512 10364 23820 10373
rect 23512 10362 23518 10364
rect 23574 10362 23598 10364
rect 23654 10362 23678 10364
rect 23734 10362 23758 10364
rect 23814 10362 23820 10364
rect 23574 10310 23576 10362
rect 23756 10310 23758 10362
rect 23512 10308 23518 10310
rect 23574 10308 23598 10310
rect 23654 10308 23678 10310
rect 23734 10308 23758 10310
rect 23814 10308 23820 10310
rect 23512 10299 23820 10308
rect 23388 10192 23440 10198
rect 23388 10134 23440 10140
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 22376 9104 22428 9110
rect 22374 9072 22376 9081
rect 22428 9072 22430 9081
rect 21744 9042 22232 9058
rect 21732 9036 22244 9042
rect 21784 9030 22192 9036
rect 21732 8978 21784 8984
rect 22374 9007 22430 9016
rect 22192 8978 22244 8984
rect 21640 8900 21692 8906
rect 21640 8842 21692 8848
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21192 8430 21220 8774
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21180 8288 21232 8294
rect 21100 8248 21180 8276
rect 21180 8230 21232 8236
rect 21468 8022 21496 8434
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21744 7954 21772 8978
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 22928 8968 22980 8974
rect 23308 8945 23336 9590
rect 22928 8910 22980 8916
rect 23294 8936 23350 8945
rect 21928 8786 21956 8910
rect 22006 8800 22062 8809
rect 21928 8758 22006 8786
rect 21824 8628 21876 8634
rect 21928 8616 21956 8758
rect 22006 8735 22062 8744
rect 21876 8588 21956 8616
rect 21824 8570 21876 8576
rect 22836 8560 22888 8566
rect 22834 8528 22836 8537
rect 22888 8528 22890 8537
rect 22834 8463 22890 8472
rect 21914 8392 21970 8401
rect 21914 8327 21916 8336
rect 21968 8327 21970 8336
rect 21916 8298 21968 8304
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 21008 7002 21036 7142
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20812 6384 20864 6390
rect 20812 6326 20864 6332
rect 20916 6254 20944 6598
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 20350 5743 20352 5752
rect 20404 5743 20406 5752
rect 20456 5766 20576 5794
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 20916 5778 20944 6190
rect 20812 5772 20864 5778
rect 20352 5714 20404 5720
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20456 4690 20484 5766
rect 20812 5714 20864 5720
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20720 5704 20772 5710
rect 20640 5652 20720 5658
rect 20640 5646 20772 5652
rect 20640 5630 20760 5646
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20548 5370 20576 5510
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20534 5264 20590 5273
rect 20534 5199 20590 5208
rect 20548 5030 20576 5199
rect 20640 5166 20668 5630
rect 20824 5370 20852 5714
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20916 5302 20944 5714
rect 20994 5536 21050 5545
rect 20994 5471 21050 5480
rect 20904 5296 20956 5302
rect 20904 5238 20956 5244
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 21008 4690 21036 5471
rect 21100 5098 21128 6938
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21088 5092 21140 5098
rect 21088 5034 21140 5040
rect 21192 4826 21220 6598
rect 21284 6322 21312 6802
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21272 6180 21324 6186
rect 21272 6122 21324 6128
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 19660 4380 19968 4389
rect 19660 4378 19666 4380
rect 19722 4378 19746 4380
rect 19802 4378 19826 4380
rect 19882 4378 19906 4380
rect 19962 4378 19968 4380
rect 19722 4326 19724 4378
rect 19904 4326 19906 4378
rect 19660 4324 19666 4326
rect 19722 4324 19746 4326
rect 19802 4324 19826 4326
rect 19882 4324 19906 4326
rect 19962 4324 19968 4326
rect 19660 4315 19968 4324
rect 19524 4208 19576 4214
rect 19524 4150 19576 4156
rect 20628 4208 20680 4214
rect 20628 4150 20680 4156
rect 19660 3292 19968 3301
rect 19660 3290 19666 3292
rect 19722 3290 19746 3292
rect 19802 3290 19826 3292
rect 19882 3290 19906 3292
rect 19962 3290 19968 3292
rect 19722 3238 19724 3290
rect 19904 3238 19906 3290
rect 19660 3236 19666 3238
rect 19722 3236 19746 3238
rect 19802 3236 19826 3238
rect 19882 3236 19906 3238
rect 19962 3236 19968 3238
rect 19660 3227 19968 3236
rect 19444 2746 20024 2774
rect 19660 2204 19968 2213
rect 19660 2202 19666 2204
rect 19722 2202 19746 2204
rect 19802 2202 19826 2204
rect 19882 2202 19906 2204
rect 19962 2202 19968 2204
rect 19722 2150 19724 2202
rect 19904 2150 19906 2202
rect 19660 2148 19666 2150
rect 19722 2148 19746 2150
rect 19802 2148 19826 2150
rect 19882 2148 19906 2150
rect 19962 2148 19968 2150
rect 19660 2139 19968 2148
rect 19660 1116 19968 1125
rect 19660 1114 19666 1116
rect 19722 1114 19746 1116
rect 19802 1114 19826 1116
rect 19882 1114 19906 1116
rect 19962 1114 19968 1116
rect 19722 1062 19724 1114
rect 19904 1062 19906 1114
rect 19660 1060 19666 1062
rect 19722 1060 19746 1062
rect 19802 1060 19826 1062
rect 19882 1060 19906 1062
rect 19962 1060 19968 1062
rect 19660 1051 19968 1060
rect 19996 400 20024 2746
rect 20640 400 20668 4150
rect 21284 400 21312 6122
rect 21376 5846 21404 7210
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21456 6112 21508 6118
rect 21456 6054 21508 6060
rect 21364 5840 21416 5846
rect 21364 5782 21416 5788
rect 21468 5778 21496 6054
rect 21560 5817 21588 7142
rect 21744 6458 21772 7686
rect 21928 7410 21956 7958
rect 22940 7954 22968 8910
rect 23294 8871 23350 8880
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 23032 8430 23060 8774
rect 23400 8566 23428 10134
rect 23848 9512 23900 9518
rect 23848 9454 23900 9460
rect 23512 9276 23820 9285
rect 23512 9274 23518 9276
rect 23574 9274 23598 9276
rect 23654 9274 23678 9276
rect 23734 9274 23758 9276
rect 23814 9274 23820 9276
rect 23574 9222 23576 9274
rect 23756 9222 23758 9274
rect 23512 9220 23518 9222
rect 23574 9220 23598 9222
rect 23654 9220 23678 9222
rect 23734 9220 23758 9222
rect 23814 9220 23820 9222
rect 23512 9211 23820 9220
rect 23860 9178 23888 9454
rect 23952 9382 23980 11018
rect 24032 11008 24084 11014
rect 24032 10950 24084 10956
rect 24044 10810 24072 10950
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 24228 10690 24256 11070
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24044 10662 24256 10690
rect 24044 10470 24072 10662
rect 24320 10606 24348 10950
rect 24504 10674 24532 11070
rect 24584 11008 24636 11014
rect 24584 10950 24636 10956
rect 24492 10668 24544 10674
rect 24492 10610 24544 10616
rect 24596 10606 24624 10950
rect 24688 10810 24716 11154
rect 25148 11150 25176 11494
rect 25424 11354 25452 11494
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 28276 11286 28304 11591
rect 31217 11452 31525 11461
rect 31217 11450 31223 11452
rect 31279 11450 31303 11452
rect 31359 11450 31383 11452
rect 31439 11450 31463 11452
rect 31519 11450 31525 11452
rect 31279 11398 31281 11450
rect 31461 11398 31463 11450
rect 31217 11396 31223 11398
rect 31279 11396 31303 11398
rect 31359 11396 31383 11398
rect 31439 11396 31463 11398
rect 31519 11396 31525 11398
rect 31217 11387 31525 11396
rect 28264 11280 28316 11286
rect 28264 11222 28316 11228
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 24860 11008 24912 11014
rect 24860 10950 24912 10956
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 24872 10810 24900 10950
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24308 10600 24360 10606
rect 24308 10542 24360 10548
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24044 10130 24072 10406
rect 24032 10124 24084 10130
rect 24032 10066 24084 10072
rect 24044 9625 24072 10066
rect 24228 9722 24256 10406
rect 24964 10198 24992 10950
rect 25240 10810 25268 11154
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 28262 10976 28318 10985
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25332 10606 25360 10950
rect 27365 10908 27673 10917
rect 28262 10911 28318 10920
rect 27365 10906 27371 10908
rect 27427 10906 27451 10908
rect 27507 10906 27531 10908
rect 27587 10906 27611 10908
rect 27667 10906 27673 10908
rect 27427 10854 27429 10906
rect 27609 10854 27611 10906
rect 27365 10852 27371 10854
rect 27427 10852 27451 10854
rect 27507 10852 27531 10854
rect 27587 10852 27611 10854
rect 27667 10852 27673 10854
rect 27365 10843 27673 10852
rect 28276 10742 28304 10911
rect 28264 10736 28316 10742
rect 28264 10678 28316 10684
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 24768 10124 24820 10130
rect 25044 10124 25096 10130
rect 24820 10084 24900 10112
rect 24768 10066 24820 10072
rect 24872 9994 24900 10084
rect 25044 10066 25096 10072
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24308 9920 24360 9926
rect 24308 9862 24360 9868
rect 24400 9920 24452 9926
rect 24400 9862 24452 9868
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24216 9716 24268 9722
rect 24216 9658 24268 9664
rect 24030 9616 24086 9625
rect 24086 9574 24164 9602
rect 24030 9551 24086 9560
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 23480 9104 23532 9110
rect 23480 9046 23532 9052
rect 23492 8566 23520 9046
rect 23848 8832 23900 8838
rect 23952 8809 23980 9114
rect 23848 8774 23900 8780
rect 23938 8800 23994 8809
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23480 8560 23532 8566
rect 23480 8502 23532 8508
rect 23020 8424 23072 8430
rect 23020 8366 23072 8372
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23032 8090 23060 8230
rect 23512 8188 23820 8197
rect 23512 8186 23518 8188
rect 23574 8186 23598 8188
rect 23654 8186 23678 8188
rect 23734 8186 23758 8188
rect 23814 8186 23820 8188
rect 23574 8134 23576 8186
rect 23756 8134 23758 8186
rect 23512 8132 23518 8134
rect 23574 8132 23598 8134
rect 23654 8132 23678 8134
rect 23734 8132 23758 8134
rect 23814 8132 23820 8134
rect 23512 8123 23820 8132
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 22928 7948 22980 7954
rect 22928 7890 22980 7896
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 21928 6866 21956 7346
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 21836 6458 21864 6802
rect 22006 6624 22062 6633
rect 22006 6559 22062 6568
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 21638 6352 21694 6361
rect 21928 6338 21956 6394
rect 21638 6287 21694 6296
rect 21836 6310 21956 6338
rect 21546 5808 21602 5817
rect 21456 5772 21508 5778
rect 21652 5778 21680 6287
rect 21732 6248 21784 6254
rect 21730 6216 21732 6225
rect 21784 6216 21786 6225
rect 21730 6151 21786 6160
rect 21836 5778 21864 6310
rect 22020 6254 22048 6559
rect 22112 6254 22140 7822
rect 23754 7712 23810 7721
rect 23754 7647 23810 7656
rect 23768 7478 23796 7647
rect 23388 7472 23440 7478
rect 23308 7432 23388 7460
rect 23112 7200 23164 7206
rect 23204 7200 23256 7206
rect 23112 7142 23164 7148
rect 23202 7168 23204 7177
rect 23256 7168 23258 7177
rect 23124 6916 23152 7142
rect 23202 7103 23258 7112
rect 23308 6984 23336 7432
rect 23388 7414 23440 7420
rect 23756 7472 23808 7478
rect 23756 7414 23808 7420
rect 23512 7100 23820 7109
rect 23512 7098 23518 7100
rect 23574 7098 23598 7100
rect 23654 7098 23678 7100
rect 23734 7098 23758 7100
rect 23814 7098 23820 7100
rect 23574 7046 23576 7098
rect 23756 7046 23758 7098
rect 23512 7044 23518 7046
rect 23574 7044 23598 7046
rect 23654 7044 23678 7046
rect 23734 7044 23758 7046
rect 23814 7044 23820 7046
rect 23512 7035 23820 7044
rect 23308 6956 23612 6984
rect 22650 6896 22706 6905
rect 22572 6854 22650 6882
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22204 6254 22232 6598
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22192 6248 22244 6254
rect 22284 6248 22336 6254
rect 22192 6190 22244 6196
rect 22282 6216 22284 6225
rect 22336 6216 22338 6225
rect 22282 6151 22338 6160
rect 22284 6112 22336 6118
rect 21914 6080 21970 6089
rect 22284 6054 22336 6060
rect 21914 6015 21970 6024
rect 21928 5914 21956 6015
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 21928 5778 21956 5850
rect 22006 5808 22062 5817
rect 21546 5743 21602 5752
rect 21640 5772 21692 5778
rect 21456 5714 21508 5720
rect 21640 5714 21692 5720
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21916 5772 21968 5778
rect 22006 5743 22062 5752
rect 21916 5714 21968 5720
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21376 4554 21404 5646
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21454 5400 21510 5409
rect 21454 5335 21456 5344
rect 21508 5335 21510 5344
rect 21456 5306 21508 5312
rect 21560 5166 21588 5578
rect 21916 5568 21968 5574
rect 21916 5510 21968 5516
rect 21928 5302 21956 5510
rect 22020 5370 22048 5743
rect 22190 5672 22246 5681
rect 22190 5607 22246 5616
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 21916 5296 21968 5302
rect 21916 5238 21968 5244
rect 22100 5296 22152 5302
rect 22100 5238 22152 5244
rect 22112 5166 22140 5238
rect 21548 5160 21600 5166
rect 21548 5102 21600 5108
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 21928 4826 21956 5102
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 21364 4548 21416 4554
rect 21364 4490 21416 4496
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21928 400 21956 4218
rect 18340 326 18644 354
rect 18694 0 18750 400
rect 19338 0 19394 400
rect 19982 0 20038 400
rect 20626 0 20682 400
rect 21270 0 21326 400
rect 21914 0 21970 400
rect 22204 354 22232 5607
rect 22296 5273 22324 6054
rect 22388 5642 22416 6734
rect 22466 5944 22522 5953
rect 22572 5914 22600 6854
rect 23124 6888 23244 6916
rect 22650 6831 22706 6840
rect 23216 6780 23244 6888
rect 23584 6866 23612 6956
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 23296 6792 23348 6798
rect 23110 6760 23166 6769
rect 23110 6695 23166 6704
rect 23216 6752 23296 6780
rect 23124 6662 23152 6695
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 22744 6656 22796 6662
rect 22744 6598 22796 6604
rect 23112 6656 23164 6662
rect 23112 6598 23164 6604
rect 22664 6225 22692 6598
rect 22650 6216 22706 6225
rect 22650 6151 22706 6160
rect 22466 5879 22522 5888
rect 22560 5908 22612 5914
rect 22480 5778 22508 5879
rect 22560 5850 22612 5856
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 22376 5636 22428 5642
rect 22376 5578 22428 5584
rect 22282 5264 22338 5273
rect 22282 5199 22338 5208
rect 22756 5030 22784 6598
rect 22928 6180 22980 6186
rect 22928 6122 22980 6128
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22848 4622 22876 6054
rect 22940 5642 22968 6122
rect 23032 5817 23060 6122
rect 23124 6089 23152 6598
rect 23216 6254 23244 6752
rect 23296 6734 23348 6740
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 23492 6361 23520 6598
rect 23676 6458 23704 6802
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23478 6352 23534 6361
rect 23768 6322 23796 6598
rect 23478 6287 23534 6296
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23204 6248 23256 6254
rect 23204 6190 23256 6196
rect 23388 6248 23440 6254
rect 23388 6190 23440 6196
rect 23296 6112 23348 6118
rect 23110 6080 23166 6089
rect 23296 6054 23348 6060
rect 23110 6015 23166 6024
rect 23308 5914 23336 6054
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 23018 5808 23074 5817
rect 23018 5743 23074 5752
rect 22928 5636 22980 5642
rect 22928 5578 22980 5584
rect 22940 5234 22968 5578
rect 23400 5234 23428 6190
rect 23860 6186 23888 8774
rect 23938 8735 23994 8744
rect 23952 7410 23980 8735
rect 24044 8634 24072 9318
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 24136 8430 24164 9574
rect 24320 9518 24348 9862
rect 24412 9722 24440 9862
rect 24688 9722 24716 9862
rect 24400 9716 24452 9722
rect 24400 9658 24452 9664
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 24308 9512 24360 9518
rect 24584 9512 24636 9518
rect 24308 9454 24360 9460
rect 24412 9472 24584 9500
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 24124 8424 24176 8430
rect 24412 8378 24440 9472
rect 24584 9454 24636 9460
rect 24768 9444 24820 9450
rect 24768 9386 24820 9392
rect 24584 8832 24636 8838
rect 24780 8820 24808 9386
rect 24872 9110 24900 9930
rect 25056 9178 25084 10066
rect 25148 9722 25176 10066
rect 25228 9920 25280 9926
rect 25228 9862 25280 9868
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 24860 9104 24912 9110
rect 24860 9046 24912 9052
rect 24636 8792 24808 8820
rect 24584 8774 24636 8780
rect 24596 8498 24624 8774
rect 25240 8634 25268 9862
rect 25332 9722 25360 10066
rect 25504 9920 25556 9926
rect 25504 9862 25556 9868
rect 25320 9716 25372 9722
rect 25320 9658 25372 9664
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 25332 9178 25360 9454
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25412 8900 25464 8906
rect 25412 8842 25464 8848
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 24124 8366 24176 8372
rect 23940 7404 23992 7410
rect 23940 7346 23992 7352
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23952 6202 23980 6938
rect 24044 6934 24072 8366
rect 24320 8350 24440 8378
rect 24584 8356 24636 8362
rect 24124 8288 24176 8294
rect 24124 8230 24176 8236
rect 24136 7342 24164 8230
rect 24214 7576 24270 7585
rect 24214 7511 24270 7520
rect 24228 7342 24256 7511
rect 24124 7336 24176 7342
rect 24124 7278 24176 7284
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 24032 6928 24084 6934
rect 24136 6905 24164 7142
rect 24032 6870 24084 6876
rect 24122 6896 24178 6905
rect 24228 6866 24256 7278
rect 24122 6831 24178 6840
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 24124 6792 24176 6798
rect 24124 6734 24176 6740
rect 23848 6180 23900 6186
rect 23952 6174 24072 6202
rect 23848 6122 23900 6128
rect 23512 6012 23820 6021
rect 23512 6010 23518 6012
rect 23574 6010 23598 6012
rect 23654 6010 23678 6012
rect 23734 6010 23758 6012
rect 23814 6010 23820 6012
rect 23574 5958 23576 6010
rect 23756 5958 23758 6010
rect 23512 5956 23518 5958
rect 23574 5956 23598 5958
rect 23654 5956 23678 5958
rect 23734 5956 23758 5958
rect 23814 5956 23820 5958
rect 23512 5947 23820 5956
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23512 4924 23820 4933
rect 23512 4922 23518 4924
rect 23574 4922 23598 4924
rect 23654 4922 23678 4924
rect 23734 4922 23758 4924
rect 23814 4922 23820 4924
rect 23574 4870 23576 4922
rect 23756 4870 23758 4922
rect 23512 4868 23518 4870
rect 23574 4868 23598 4870
rect 23654 4868 23678 4870
rect 23734 4868 23758 4870
rect 23814 4868 23820 4870
rect 23512 4859 23820 4868
rect 23860 4826 23888 6122
rect 24044 5545 24072 6174
rect 24136 5914 24164 6734
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24228 5642 24256 6802
rect 24320 6662 24348 8350
rect 24584 8298 24636 8304
rect 24596 7834 24624 8298
rect 25044 8288 25096 8294
rect 24674 8256 24730 8265
rect 25044 8230 25096 8236
rect 24674 8191 24730 8200
rect 24412 7806 24624 7834
rect 24412 6866 24440 7806
rect 24688 7698 24716 8191
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24504 7670 24716 7698
rect 24504 7546 24532 7670
rect 24492 7540 24544 7546
rect 24492 7482 24544 7488
rect 24584 7540 24636 7546
rect 24584 7482 24636 7488
rect 24492 7336 24544 7342
rect 24492 7278 24544 7284
rect 24504 7177 24532 7278
rect 24490 7168 24546 7177
rect 24490 7103 24546 7112
rect 24596 7002 24624 7482
rect 24584 6996 24636 7002
rect 24584 6938 24636 6944
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24308 6656 24360 6662
rect 24308 6598 24360 6604
rect 24504 6458 24532 6802
rect 24584 6656 24636 6662
rect 24780 6633 24808 7822
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 24584 6598 24636 6604
rect 24766 6624 24822 6633
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24216 5636 24268 5642
rect 24216 5578 24268 5584
rect 24030 5536 24086 5545
rect 24030 5471 24086 5480
rect 24596 5370 24624 6598
rect 24766 6559 24822 6568
rect 24872 5574 24900 7686
rect 25056 7342 25084 8230
rect 25240 7954 25268 8434
rect 25424 8430 25452 8842
rect 25516 8634 25544 9862
rect 25700 9722 25728 10542
rect 31668 10464 31720 10470
rect 31668 10406 31720 10412
rect 31217 10364 31525 10373
rect 31217 10362 31223 10364
rect 31279 10362 31303 10364
rect 31359 10362 31383 10364
rect 31439 10362 31463 10364
rect 31519 10362 31525 10364
rect 31279 10310 31281 10362
rect 31461 10310 31463 10362
rect 31217 10308 31223 10310
rect 31279 10308 31303 10310
rect 31359 10308 31383 10310
rect 31439 10308 31463 10310
rect 31519 10308 31525 10310
rect 31217 10299 31525 10308
rect 31680 10305 31708 10406
rect 31666 10296 31722 10305
rect 28264 10260 28316 10266
rect 31666 10231 31722 10240
rect 28264 10202 28316 10208
rect 26148 10192 26200 10198
rect 26148 10134 26200 10140
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 25964 9988 26016 9994
rect 25964 9930 26016 9936
rect 25688 9716 25740 9722
rect 25688 9658 25740 9664
rect 25872 9512 25924 9518
rect 25872 9454 25924 9460
rect 25884 9178 25912 9454
rect 25976 9178 26004 9930
rect 26068 9654 26096 9998
rect 26160 9654 26188 10134
rect 26240 9920 26292 9926
rect 26240 9862 26292 9868
rect 26056 9648 26108 9654
rect 26056 9590 26108 9596
rect 26148 9648 26200 9654
rect 26148 9590 26200 9596
rect 26252 9518 26280 9862
rect 27365 9820 27673 9829
rect 27365 9818 27371 9820
rect 27427 9818 27451 9820
rect 27507 9818 27531 9820
rect 27587 9818 27611 9820
rect 27667 9818 27673 9820
rect 27427 9766 27429 9818
rect 27609 9766 27611 9818
rect 27365 9764 27371 9766
rect 27427 9764 27451 9766
rect 27507 9764 27531 9766
rect 27587 9764 27611 9766
rect 27667 9764 27673 9766
rect 27365 9755 27673 9764
rect 28276 9625 28304 10202
rect 28262 9616 28318 9625
rect 28262 9551 28318 9560
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26976 9376 27028 9382
rect 26976 9318 27028 9324
rect 25872 9172 25924 9178
rect 25872 9114 25924 9120
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 26056 9036 26108 9042
rect 26056 8978 26108 8984
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25608 8537 25636 8774
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25594 8528 25650 8537
rect 25594 8463 25650 8472
rect 25412 8424 25464 8430
rect 25700 8378 25728 8570
rect 25412 8366 25464 8372
rect 25516 8350 25728 8378
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 25516 8022 25544 8350
rect 25596 8288 25648 8294
rect 25596 8230 25648 8236
rect 25608 8090 25636 8230
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 25504 8016 25556 8022
rect 25504 7958 25556 7964
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 25228 7948 25280 7954
rect 25228 7890 25280 7896
rect 25412 7948 25464 7954
rect 25412 7890 25464 7896
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 24964 6730 24992 7278
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 25056 6769 25084 7142
rect 25042 6760 25098 6769
rect 24952 6724 25004 6730
rect 25042 6695 25098 6704
rect 24952 6666 25004 6672
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 25148 5409 25176 7890
rect 25228 7472 25280 7478
rect 25228 7414 25280 7420
rect 25240 6934 25268 7414
rect 25424 7342 25452 7890
rect 25596 7880 25648 7886
rect 25884 7868 25912 8366
rect 25648 7840 25912 7868
rect 25596 7822 25648 7828
rect 25504 7812 25556 7818
rect 25504 7754 25556 7760
rect 25516 7426 25544 7754
rect 25688 7744 25740 7750
rect 25594 7712 25650 7721
rect 25688 7686 25740 7692
rect 25780 7744 25832 7750
rect 25780 7686 25832 7692
rect 25872 7744 25924 7750
rect 25872 7686 25924 7692
rect 25594 7647 25650 7656
rect 25608 7546 25636 7647
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25516 7398 25636 7426
rect 25412 7336 25464 7342
rect 25412 7278 25464 7284
rect 25504 7336 25556 7342
rect 25504 7278 25556 7284
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 25228 6928 25280 6934
rect 25228 6870 25280 6876
rect 25332 6254 25360 7142
rect 25516 7002 25544 7278
rect 25504 6996 25556 7002
rect 25504 6938 25556 6944
rect 25608 6905 25636 7398
rect 25594 6896 25650 6905
rect 25594 6831 25650 6840
rect 25320 6248 25372 6254
rect 25320 6190 25372 6196
rect 25134 5400 25190 5409
rect 24584 5364 24636 5370
rect 25134 5335 25190 5344
rect 24584 5306 24636 5312
rect 25700 5302 25728 7686
rect 25792 7546 25820 7686
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 25884 5710 25912 7686
rect 25976 7177 26004 8774
rect 26068 8566 26096 8978
rect 26252 8906 26280 9318
rect 26988 9178 27016 9318
rect 31217 9276 31525 9285
rect 31217 9274 31223 9276
rect 31279 9274 31303 9276
rect 31359 9274 31383 9276
rect 31439 9274 31463 9276
rect 31519 9274 31525 9276
rect 31279 9222 31281 9274
rect 31461 9222 31463 9274
rect 31217 9220 31223 9222
rect 31279 9220 31303 9222
rect 31359 9220 31383 9222
rect 31439 9220 31463 9222
rect 31519 9220 31525 9222
rect 31217 9211 31525 9220
rect 26976 9172 27028 9178
rect 26976 9114 27028 9120
rect 26240 8900 26292 8906
rect 26240 8842 26292 8848
rect 27365 8732 27673 8741
rect 27365 8730 27371 8732
rect 27427 8730 27451 8732
rect 27507 8730 27531 8732
rect 27587 8730 27611 8732
rect 27667 8730 27673 8732
rect 27427 8678 27429 8730
rect 27609 8678 27611 8730
rect 27365 8676 27371 8678
rect 27427 8676 27451 8678
rect 27507 8676 27531 8678
rect 27587 8676 27611 8678
rect 27667 8676 27673 8678
rect 27365 8667 27673 8676
rect 26056 8560 26108 8566
rect 26056 8502 26108 8508
rect 31666 8528 31722 8537
rect 31666 8463 31722 8472
rect 26332 8424 26384 8430
rect 26332 8366 26384 8372
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 25962 7168 26018 7177
rect 25962 7103 26018 7112
rect 26160 5778 26188 7686
rect 26344 7585 26372 8366
rect 31680 8265 31708 8463
rect 31666 8256 31722 8265
rect 31217 8188 31525 8197
rect 31666 8191 31722 8200
rect 31217 8186 31223 8188
rect 31279 8186 31303 8188
rect 31359 8186 31383 8188
rect 31439 8186 31463 8188
rect 31519 8186 31525 8188
rect 31279 8134 31281 8186
rect 31461 8134 31463 8186
rect 31217 8132 31223 8134
rect 31279 8132 31303 8134
rect 31359 8132 31383 8134
rect 31439 8132 31463 8134
rect 31519 8132 31525 8134
rect 31217 8123 31525 8132
rect 27365 7644 27673 7653
rect 27365 7642 27371 7644
rect 27427 7642 27451 7644
rect 27507 7642 27531 7644
rect 27587 7642 27611 7644
rect 27667 7642 27673 7644
rect 27427 7590 27429 7642
rect 27609 7590 27611 7642
rect 27365 7588 27371 7590
rect 27427 7588 27451 7590
rect 27507 7588 27531 7590
rect 27587 7588 27611 7590
rect 27667 7588 27673 7590
rect 26330 7576 26386 7585
rect 27365 7579 27673 7588
rect 26330 7511 26386 7520
rect 31666 7304 31722 7313
rect 31666 7239 31722 7248
rect 31217 7100 31525 7109
rect 31217 7098 31223 7100
rect 31279 7098 31303 7100
rect 31359 7098 31383 7100
rect 31439 7098 31463 7100
rect 31519 7098 31525 7100
rect 31279 7046 31281 7098
rect 31461 7046 31463 7098
rect 31217 7044 31223 7046
rect 31279 7044 31303 7046
rect 31359 7044 31383 7046
rect 31439 7044 31463 7046
rect 31519 7044 31525 7046
rect 31217 7035 31525 7044
rect 27365 6556 27673 6565
rect 27365 6554 27371 6556
rect 27427 6554 27451 6556
rect 27507 6554 27531 6556
rect 27587 6554 27611 6556
rect 27667 6554 27673 6556
rect 27427 6502 27429 6554
rect 27609 6502 27611 6554
rect 27365 6500 27371 6502
rect 27427 6500 27451 6502
rect 27507 6500 27531 6502
rect 27587 6500 27611 6502
rect 27667 6500 27673 6502
rect 27365 6491 27673 6500
rect 31217 6012 31525 6021
rect 31217 6010 31223 6012
rect 31279 6010 31303 6012
rect 31359 6010 31383 6012
rect 31439 6010 31463 6012
rect 31519 6010 31525 6012
rect 31279 5958 31281 6010
rect 31461 5958 31463 6010
rect 31217 5956 31223 5958
rect 31279 5956 31303 5958
rect 31359 5956 31383 5958
rect 31439 5956 31463 5958
rect 31519 5956 31525 5958
rect 31217 5947 31525 5956
rect 26148 5772 26200 5778
rect 26148 5714 26200 5720
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 27365 5468 27673 5477
rect 27365 5466 27371 5468
rect 27427 5466 27451 5468
rect 27507 5466 27531 5468
rect 27587 5466 27611 5468
rect 27667 5466 27673 5468
rect 27427 5414 27429 5466
rect 27609 5414 27611 5466
rect 27365 5412 27371 5414
rect 27427 5412 27451 5414
rect 27507 5412 27531 5414
rect 27587 5412 27611 5414
rect 27667 5412 27673 5414
rect 27365 5403 27673 5412
rect 25688 5296 25740 5302
rect 25688 5238 25740 5244
rect 31217 4924 31525 4933
rect 31217 4922 31223 4924
rect 31279 4922 31303 4924
rect 31359 4922 31383 4924
rect 31439 4922 31463 4924
rect 31519 4922 31525 4924
rect 31279 4870 31281 4922
rect 31461 4870 31463 4922
rect 31217 4868 31223 4870
rect 31279 4868 31303 4870
rect 31359 4868 31383 4870
rect 31439 4868 31463 4870
rect 31519 4868 31525 4870
rect 31217 4859 31525 4868
rect 31680 4865 31708 7239
rect 31666 4856 31722 4865
rect 23848 4820 23900 4826
rect 31666 4791 31722 4800
rect 23848 4762 23900 4768
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 27365 4380 27673 4389
rect 27365 4378 27371 4380
rect 27427 4378 27451 4380
rect 27507 4378 27531 4380
rect 27587 4378 27611 4380
rect 27667 4378 27673 4380
rect 27427 4326 27429 4378
rect 27609 4326 27611 4378
rect 27365 4324 27371 4326
rect 27427 4324 27451 4326
rect 27507 4324 27531 4326
rect 27587 4324 27611 4326
rect 27667 4324 27673 4326
rect 27365 4315 27673 4324
rect 23512 3836 23820 3845
rect 23512 3834 23518 3836
rect 23574 3834 23598 3836
rect 23654 3834 23678 3836
rect 23734 3834 23758 3836
rect 23814 3834 23820 3836
rect 23574 3782 23576 3834
rect 23756 3782 23758 3834
rect 23512 3780 23518 3782
rect 23574 3780 23598 3782
rect 23654 3780 23678 3782
rect 23734 3780 23758 3782
rect 23814 3780 23820 3782
rect 23512 3771 23820 3780
rect 31217 3836 31525 3845
rect 31217 3834 31223 3836
rect 31279 3834 31303 3836
rect 31359 3834 31383 3836
rect 31439 3834 31463 3836
rect 31519 3834 31525 3836
rect 31279 3782 31281 3834
rect 31461 3782 31463 3834
rect 31217 3780 31223 3782
rect 31279 3780 31303 3782
rect 31359 3780 31383 3782
rect 31439 3780 31463 3782
rect 31519 3780 31525 3782
rect 31217 3771 31525 3780
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 22480 462 22600 490
rect 22480 354 22508 462
rect 22572 400 22600 462
rect 23216 400 23244 3334
rect 27365 3292 27673 3301
rect 27365 3290 27371 3292
rect 27427 3290 27451 3292
rect 27507 3290 27531 3292
rect 27587 3290 27611 3292
rect 27667 3290 27673 3292
rect 27427 3238 27429 3290
rect 27609 3238 27611 3290
rect 27365 3236 27371 3238
rect 27427 3236 27451 3238
rect 27507 3236 27531 3238
rect 27587 3236 27611 3238
rect 27667 3236 27673 3238
rect 27365 3227 27673 3236
rect 23512 2748 23820 2757
rect 23512 2746 23518 2748
rect 23574 2746 23598 2748
rect 23654 2746 23678 2748
rect 23734 2746 23758 2748
rect 23814 2746 23820 2748
rect 23574 2694 23576 2746
rect 23756 2694 23758 2746
rect 23512 2692 23518 2694
rect 23574 2692 23598 2694
rect 23654 2692 23678 2694
rect 23734 2692 23758 2694
rect 23814 2692 23820 2694
rect 23512 2683 23820 2692
rect 31217 2748 31525 2757
rect 31217 2746 31223 2748
rect 31279 2746 31303 2748
rect 31359 2746 31383 2748
rect 31439 2746 31463 2748
rect 31519 2746 31525 2748
rect 31279 2694 31281 2746
rect 31461 2694 31463 2746
rect 31217 2692 31223 2694
rect 31279 2692 31303 2694
rect 31359 2692 31383 2694
rect 31439 2692 31463 2694
rect 31519 2692 31525 2694
rect 31217 2683 31525 2692
rect 27365 2204 27673 2213
rect 27365 2202 27371 2204
rect 27427 2202 27451 2204
rect 27507 2202 27531 2204
rect 27587 2202 27611 2204
rect 27667 2202 27673 2204
rect 27427 2150 27429 2202
rect 27609 2150 27611 2202
rect 27365 2148 27371 2150
rect 27427 2148 27451 2150
rect 27507 2148 27531 2150
rect 27587 2148 27611 2150
rect 27667 2148 27673 2150
rect 27365 2139 27673 2148
rect 23512 1660 23820 1669
rect 23512 1658 23518 1660
rect 23574 1658 23598 1660
rect 23654 1658 23678 1660
rect 23734 1658 23758 1660
rect 23814 1658 23820 1660
rect 23574 1606 23576 1658
rect 23756 1606 23758 1658
rect 23512 1604 23518 1606
rect 23574 1604 23598 1606
rect 23654 1604 23678 1606
rect 23734 1604 23758 1606
rect 23814 1604 23820 1606
rect 23512 1595 23820 1604
rect 31217 1660 31525 1669
rect 31217 1658 31223 1660
rect 31279 1658 31303 1660
rect 31359 1658 31383 1660
rect 31439 1658 31463 1660
rect 31519 1658 31525 1660
rect 31279 1606 31281 1658
rect 31461 1606 31463 1658
rect 31217 1604 31223 1606
rect 31279 1604 31303 1606
rect 31359 1604 31383 1606
rect 31439 1604 31463 1606
rect 31519 1604 31525 1606
rect 31217 1595 31525 1604
rect 27365 1116 27673 1125
rect 27365 1114 27371 1116
rect 27427 1114 27451 1116
rect 27507 1114 27531 1116
rect 27587 1114 27611 1116
rect 27667 1114 27673 1116
rect 27427 1062 27429 1114
rect 27609 1062 27611 1114
rect 27365 1060 27371 1062
rect 27427 1060 27451 1062
rect 27507 1060 27531 1062
rect 27587 1060 27611 1062
rect 27667 1060 27673 1062
rect 27365 1051 27673 1060
rect 23512 572 23820 581
rect 23512 570 23518 572
rect 23574 570 23598 572
rect 23654 570 23678 572
rect 23734 570 23758 572
rect 23814 570 23820 572
rect 23574 518 23576 570
rect 23756 518 23758 570
rect 23512 516 23518 518
rect 23574 516 23598 518
rect 23654 516 23678 518
rect 23734 516 23758 518
rect 23814 516 23820 518
rect 23512 507 23820 516
rect 31217 572 31525 581
rect 31217 570 31223 572
rect 31279 570 31303 572
rect 31359 570 31383 572
rect 31439 570 31463 572
rect 31519 570 31525 572
rect 31279 518 31281 570
rect 31461 518 31463 570
rect 31217 516 31223 518
rect 31279 516 31303 518
rect 31359 516 31383 518
rect 31439 516 31463 518
rect 31519 516 31525 518
rect 31217 507 31525 516
rect 22204 326 22508 354
rect 22558 0 22614 400
rect 23202 0 23258 400
<< via2 >>
rect 8108 19066 8164 19068
rect 8188 19066 8244 19068
rect 8268 19066 8324 19068
rect 8348 19066 8404 19068
rect 8108 19014 8154 19066
rect 8154 19014 8164 19066
rect 8188 19014 8218 19066
rect 8218 19014 8230 19066
rect 8230 19014 8244 19066
rect 8268 19014 8282 19066
rect 8282 19014 8294 19066
rect 8294 19014 8324 19066
rect 8348 19014 8358 19066
rect 8358 19014 8404 19066
rect 8108 19012 8164 19014
rect 8188 19012 8244 19014
rect 8268 19012 8324 19014
rect 8348 19012 8404 19014
rect 4256 18522 4312 18524
rect 4336 18522 4392 18524
rect 4416 18522 4472 18524
rect 4496 18522 4552 18524
rect 4256 18470 4302 18522
rect 4302 18470 4312 18522
rect 4336 18470 4366 18522
rect 4366 18470 4378 18522
rect 4378 18470 4392 18522
rect 4416 18470 4430 18522
rect 4430 18470 4442 18522
rect 4442 18470 4472 18522
rect 4496 18470 4506 18522
rect 4506 18470 4552 18522
rect 4256 18468 4312 18470
rect 4336 18468 4392 18470
rect 4416 18468 4472 18470
rect 4496 18468 4552 18470
rect 8108 17978 8164 17980
rect 8188 17978 8244 17980
rect 8268 17978 8324 17980
rect 8348 17978 8404 17980
rect 8108 17926 8154 17978
rect 8154 17926 8164 17978
rect 8188 17926 8218 17978
rect 8218 17926 8230 17978
rect 8230 17926 8244 17978
rect 8268 17926 8282 17978
rect 8282 17926 8294 17978
rect 8294 17926 8324 17978
rect 8348 17926 8358 17978
rect 8358 17926 8404 17978
rect 8108 17924 8164 17926
rect 8188 17924 8244 17926
rect 8268 17924 8324 17926
rect 8348 17924 8404 17926
rect 4256 17434 4312 17436
rect 4336 17434 4392 17436
rect 4416 17434 4472 17436
rect 4496 17434 4552 17436
rect 4256 17382 4302 17434
rect 4302 17382 4312 17434
rect 4336 17382 4366 17434
rect 4366 17382 4378 17434
rect 4378 17382 4392 17434
rect 4416 17382 4430 17434
rect 4430 17382 4442 17434
rect 4442 17382 4472 17434
rect 4496 17382 4506 17434
rect 4506 17382 4552 17434
rect 4256 17380 4312 17382
rect 4336 17380 4392 17382
rect 4416 17380 4472 17382
rect 4496 17380 4552 17382
rect 8108 16890 8164 16892
rect 8188 16890 8244 16892
rect 8268 16890 8324 16892
rect 8348 16890 8404 16892
rect 8108 16838 8154 16890
rect 8154 16838 8164 16890
rect 8188 16838 8218 16890
rect 8218 16838 8230 16890
rect 8230 16838 8244 16890
rect 8268 16838 8282 16890
rect 8282 16838 8294 16890
rect 8294 16838 8324 16890
rect 8348 16838 8358 16890
rect 8358 16838 8404 16890
rect 8108 16836 8164 16838
rect 8188 16836 8244 16838
rect 8268 16836 8324 16838
rect 8348 16836 8404 16838
rect 4256 16346 4312 16348
rect 4336 16346 4392 16348
rect 4416 16346 4472 16348
rect 4496 16346 4552 16348
rect 4256 16294 4302 16346
rect 4302 16294 4312 16346
rect 4336 16294 4366 16346
rect 4366 16294 4378 16346
rect 4378 16294 4392 16346
rect 4416 16294 4430 16346
rect 4430 16294 4442 16346
rect 4442 16294 4472 16346
rect 4496 16294 4506 16346
rect 4506 16294 4552 16346
rect 4256 16292 4312 16294
rect 4336 16292 4392 16294
rect 4416 16292 4472 16294
rect 4496 16292 4552 16294
rect 7378 15272 7434 15328
rect 4256 15258 4312 15260
rect 4336 15258 4392 15260
rect 4416 15258 4472 15260
rect 4496 15258 4552 15260
rect 4256 15206 4302 15258
rect 4302 15206 4312 15258
rect 4336 15206 4366 15258
rect 4366 15206 4378 15258
rect 4378 15206 4392 15258
rect 4416 15206 4430 15258
rect 4430 15206 4442 15258
rect 4442 15206 4472 15258
rect 4496 15206 4506 15258
rect 4506 15206 4552 15258
rect 4256 15204 4312 15206
rect 4336 15204 4392 15206
rect 4416 15204 4472 15206
rect 4496 15204 4552 15206
rect 4256 14170 4312 14172
rect 4336 14170 4392 14172
rect 4416 14170 4472 14172
rect 4496 14170 4552 14172
rect 4256 14118 4302 14170
rect 4302 14118 4312 14170
rect 4336 14118 4366 14170
rect 4366 14118 4378 14170
rect 4378 14118 4392 14170
rect 4416 14118 4430 14170
rect 4430 14118 4442 14170
rect 4442 14118 4472 14170
rect 4496 14118 4506 14170
rect 4506 14118 4552 14170
rect 4256 14116 4312 14118
rect 4336 14116 4392 14118
rect 4416 14116 4472 14118
rect 4496 14116 4552 14118
rect 7654 14456 7710 14512
rect 7838 15952 7894 16008
rect 7838 15136 7894 15192
rect 8482 16088 8538 16144
rect 8108 15802 8164 15804
rect 8188 15802 8244 15804
rect 8268 15802 8324 15804
rect 8348 15802 8404 15804
rect 8108 15750 8154 15802
rect 8154 15750 8164 15802
rect 8188 15750 8218 15802
rect 8218 15750 8230 15802
rect 8230 15750 8244 15802
rect 8268 15750 8282 15802
rect 8282 15750 8294 15802
rect 8294 15750 8324 15802
rect 8348 15750 8358 15802
rect 8358 15750 8404 15802
rect 8108 15748 8164 15750
rect 8188 15748 8244 15750
rect 8268 15748 8324 15750
rect 8348 15748 8404 15750
rect 8108 14714 8164 14716
rect 8188 14714 8244 14716
rect 8268 14714 8324 14716
rect 8348 14714 8404 14716
rect 8108 14662 8154 14714
rect 8154 14662 8164 14714
rect 8188 14662 8218 14714
rect 8218 14662 8230 14714
rect 8230 14662 8244 14714
rect 8268 14662 8282 14714
rect 8282 14662 8294 14714
rect 8294 14662 8324 14714
rect 8348 14662 8358 14714
rect 8358 14662 8404 14714
rect 8108 14660 8164 14662
rect 8188 14660 8244 14662
rect 8268 14660 8324 14662
rect 8348 14660 8404 14662
rect 4256 13082 4312 13084
rect 4336 13082 4392 13084
rect 4416 13082 4472 13084
rect 4496 13082 4552 13084
rect 4256 13030 4302 13082
rect 4302 13030 4312 13082
rect 4336 13030 4366 13082
rect 4366 13030 4378 13082
rect 4378 13030 4392 13082
rect 4416 13030 4430 13082
rect 4430 13030 4442 13082
rect 4442 13030 4472 13082
rect 4496 13030 4506 13082
rect 4506 13030 4552 13082
rect 4256 13028 4312 13030
rect 4336 13028 4392 13030
rect 4416 13028 4472 13030
rect 4496 13028 4552 13030
rect 7654 13404 7656 13424
rect 7656 13404 7708 13424
rect 7708 13404 7710 13424
rect 7654 13368 7710 13404
rect 8108 13626 8164 13628
rect 8188 13626 8244 13628
rect 8268 13626 8324 13628
rect 8348 13626 8404 13628
rect 8108 13574 8154 13626
rect 8154 13574 8164 13626
rect 8188 13574 8218 13626
rect 8218 13574 8230 13626
rect 8230 13574 8244 13626
rect 8268 13574 8282 13626
rect 8282 13574 8294 13626
rect 8294 13574 8324 13626
rect 8348 13574 8358 13626
rect 8358 13574 8404 13626
rect 8108 13572 8164 13574
rect 8188 13572 8244 13574
rect 8268 13572 8324 13574
rect 8348 13572 8404 13574
rect 9586 16224 9642 16280
rect 9126 15816 9182 15872
rect 9494 15564 9550 15600
rect 9494 15544 9496 15564
rect 9496 15544 9548 15564
rect 9548 15544 9550 15564
rect 10046 16532 10048 16552
rect 10048 16532 10100 16552
rect 10100 16532 10102 16552
rect 10046 16496 10102 16532
rect 10046 16360 10102 16416
rect 9678 15680 9734 15736
rect 8666 14864 8722 14920
rect 9310 15408 9366 15464
rect 9310 14900 9312 14920
rect 9312 14900 9364 14920
rect 9364 14900 9366 14920
rect 9310 14864 9366 14900
rect 7930 13232 7986 13288
rect 8108 12538 8164 12540
rect 8188 12538 8244 12540
rect 8268 12538 8324 12540
rect 8348 12538 8404 12540
rect 8108 12486 8154 12538
rect 8154 12486 8164 12538
rect 8188 12486 8218 12538
rect 8218 12486 8230 12538
rect 8230 12486 8244 12538
rect 8268 12486 8282 12538
rect 8282 12486 8294 12538
rect 8294 12486 8324 12538
rect 8348 12486 8358 12538
rect 8358 12486 8404 12538
rect 8108 12484 8164 12486
rect 8188 12484 8244 12486
rect 8268 12484 8324 12486
rect 8348 12484 8404 12486
rect 9310 13504 9366 13560
rect 9218 13232 9274 13288
rect 8942 12824 8998 12880
rect 4256 11994 4312 11996
rect 4336 11994 4392 11996
rect 4416 11994 4472 11996
rect 4496 11994 4552 11996
rect 4256 11942 4302 11994
rect 4302 11942 4312 11994
rect 4336 11942 4366 11994
rect 4366 11942 4378 11994
rect 4378 11942 4392 11994
rect 4416 11942 4430 11994
rect 4430 11942 4442 11994
rect 4442 11942 4472 11994
rect 4496 11942 4506 11994
rect 4506 11942 4552 11994
rect 4256 11940 4312 11942
rect 4336 11940 4392 11942
rect 4416 11940 4472 11942
rect 4496 11940 4552 11942
rect 10230 16632 10286 16688
rect 10966 16904 11022 16960
rect 10322 16496 10378 16552
rect 10138 15272 10194 15328
rect 10138 15136 10194 15192
rect 9862 15000 9918 15056
rect 9770 14864 9826 14920
rect 10138 15000 10194 15056
rect 9586 13640 9642 13696
rect 10414 15136 10470 15192
rect 10966 16652 11022 16688
rect 10966 16632 10968 16652
rect 10968 16632 11020 16652
rect 11020 16632 11022 16652
rect 11242 16360 11298 16416
rect 10966 15988 10968 16008
rect 10968 15988 11020 16008
rect 11020 15988 11022 16008
rect 10966 15952 11022 15988
rect 11150 15680 11206 15736
rect 11058 15580 11060 15600
rect 11060 15580 11112 15600
rect 11112 15580 11114 15600
rect 11058 15544 11114 15580
rect 10598 15272 10654 15328
rect 10414 14456 10470 14512
rect 10690 14728 10746 14784
rect 10046 12300 10102 12336
rect 10046 12280 10048 12300
rect 10048 12280 10100 12300
rect 10100 12280 10102 12300
rect 10966 15272 11022 15328
rect 11150 14864 11206 14920
rect 11334 15952 11390 16008
rect 11518 16224 11574 16280
rect 11334 14864 11390 14920
rect 10874 14456 10930 14512
rect 10966 13776 11022 13832
rect 12254 18672 12310 18728
rect 11961 18522 12017 18524
rect 12041 18522 12097 18524
rect 12121 18522 12177 18524
rect 12201 18522 12257 18524
rect 11961 18470 12007 18522
rect 12007 18470 12017 18522
rect 12041 18470 12071 18522
rect 12071 18470 12083 18522
rect 12083 18470 12097 18522
rect 12121 18470 12135 18522
rect 12135 18470 12147 18522
rect 12147 18470 12177 18522
rect 12201 18470 12211 18522
rect 12211 18470 12257 18522
rect 11961 18468 12017 18470
rect 12041 18468 12097 18470
rect 12121 18468 12177 18470
rect 12201 18468 12257 18470
rect 11961 17434 12017 17436
rect 12041 17434 12097 17436
rect 12121 17434 12177 17436
rect 12201 17434 12257 17436
rect 11961 17382 12007 17434
rect 12007 17382 12017 17434
rect 12041 17382 12071 17434
rect 12071 17382 12083 17434
rect 12083 17382 12097 17434
rect 12121 17382 12135 17434
rect 12135 17382 12147 17434
rect 12147 17382 12177 17434
rect 12201 17382 12211 17434
rect 12211 17382 12257 17434
rect 11961 17380 12017 17382
rect 12041 17380 12097 17382
rect 12121 17380 12177 17382
rect 12201 17380 12257 17382
rect 11961 16346 12017 16348
rect 12041 16346 12097 16348
rect 12121 16346 12177 16348
rect 12201 16346 12257 16348
rect 11961 16294 12007 16346
rect 12007 16294 12017 16346
rect 12041 16294 12071 16346
rect 12071 16294 12083 16346
rect 12083 16294 12097 16346
rect 12121 16294 12135 16346
rect 12135 16294 12147 16346
rect 12147 16294 12177 16346
rect 12201 16294 12211 16346
rect 12211 16294 12257 16346
rect 11961 16292 12017 16294
rect 12041 16292 12097 16294
rect 12121 16292 12177 16294
rect 12201 16292 12257 16294
rect 11978 15444 11980 15464
rect 11980 15444 12032 15464
rect 12032 15444 12034 15464
rect 11978 15408 12034 15444
rect 11961 15258 12017 15260
rect 12041 15258 12097 15260
rect 12121 15258 12177 15260
rect 12201 15258 12257 15260
rect 11961 15206 12007 15258
rect 12007 15206 12017 15258
rect 12041 15206 12071 15258
rect 12071 15206 12083 15258
rect 12083 15206 12097 15258
rect 12121 15206 12135 15258
rect 12135 15206 12147 15258
rect 12147 15206 12177 15258
rect 12201 15206 12211 15258
rect 12211 15206 12257 15258
rect 11961 15204 12017 15206
rect 12041 15204 12097 15206
rect 12121 15204 12177 15206
rect 12201 15204 12257 15206
rect 11961 14170 12017 14172
rect 12041 14170 12097 14172
rect 12121 14170 12177 14172
rect 12201 14170 12257 14172
rect 11961 14118 12007 14170
rect 12007 14118 12017 14170
rect 12041 14118 12071 14170
rect 12071 14118 12083 14170
rect 12083 14118 12097 14170
rect 12121 14118 12135 14170
rect 12135 14118 12147 14170
rect 12147 14118 12177 14170
rect 12201 14118 12211 14170
rect 12211 14118 12257 14170
rect 11961 14116 12017 14118
rect 12041 14116 12097 14118
rect 12121 14116 12177 14118
rect 12201 14116 12257 14118
rect 11334 12960 11390 13016
rect 8108 11450 8164 11452
rect 8188 11450 8244 11452
rect 8268 11450 8324 11452
rect 8348 11450 8404 11452
rect 8108 11398 8154 11450
rect 8154 11398 8164 11450
rect 8188 11398 8218 11450
rect 8218 11398 8230 11450
rect 8230 11398 8244 11450
rect 8268 11398 8282 11450
rect 8282 11398 8294 11450
rect 8294 11398 8324 11450
rect 8348 11398 8358 11450
rect 8358 11398 8404 11450
rect 8108 11396 8164 11398
rect 8188 11396 8244 11398
rect 8268 11396 8324 11398
rect 8348 11396 8404 11398
rect 9494 11192 9550 11248
rect 4256 10906 4312 10908
rect 4336 10906 4392 10908
rect 4416 10906 4472 10908
rect 4496 10906 4552 10908
rect 4256 10854 4302 10906
rect 4302 10854 4312 10906
rect 4336 10854 4366 10906
rect 4366 10854 4378 10906
rect 4378 10854 4392 10906
rect 4416 10854 4430 10906
rect 4430 10854 4442 10906
rect 4442 10854 4472 10906
rect 4496 10854 4506 10906
rect 4506 10854 4552 10906
rect 4256 10852 4312 10854
rect 4336 10852 4392 10854
rect 4416 10852 4472 10854
rect 4496 10852 4552 10854
rect 4256 9818 4312 9820
rect 4336 9818 4392 9820
rect 4416 9818 4472 9820
rect 4496 9818 4552 9820
rect 4256 9766 4302 9818
rect 4302 9766 4312 9818
rect 4336 9766 4366 9818
rect 4366 9766 4378 9818
rect 4378 9766 4392 9818
rect 4416 9766 4430 9818
rect 4430 9766 4442 9818
rect 4442 9766 4472 9818
rect 4496 9766 4506 9818
rect 4506 9766 4552 9818
rect 4256 9764 4312 9766
rect 4336 9764 4392 9766
rect 4416 9764 4472 9766
rect 4496 9764 4552 9766
rect 6458 9460 6460 9480
rect 6460 9460 6512 9480
rect 6512 9460 6514 9480
rect 6458 9424 6514 9460
rect 4256 8730 4312 8732
rect 4336 8730 4392 8732
rect 4416 8730 4472 8732
rect 4496 8730 4552 8732
rect 4256 8678 4302 8730
rect 4302 8678 4312 8730
rect 4336 8678 4366 8730
rect 4366 8678 4378 8730
rect 4378 8678 4392 8730
rect 4416 8678 4430 8730
rect 4430 8678 4442 8730
rect 4442 8678 4472 8730
rect 4496 8678 4506 8730
rect 4506 8678 4552 8730
rect 4256 8676 4312 8678
rect 4336 8676 4392 8678
rect 4416 8676 4472 8678
rect 4496 8676 4552 8678
rect 8108 10362 8164 10364
rect 8188 10362 8244 10364
rect 8268 10362 8324 10364
rect 8348 10362 8404 10364
rect 8108 10310 8154 10362
rect 8154 10310 8164 10362
rect 8188 10310 8218 10362
rect 8218 10310 8230 10362
rect 8230 10310 8244 10362
rect 8268 10310 8282 10362
rect 8282 10310 8294 10362
rect 8294 10310 8324 10362
rect 8348 10310 8358 10362
rect 8358 10310 8404 10362
rect 8108 10308 8164 10310
rect 8188 10308 8244 10310
rect 8268 10308 8324 10310
rect 8348 10308 8404 10310
rect 9126 10104 9182 10160
rect 8666 9596 8668 9616
rect 8668 9596 8720 9616
rect 8720 9596 8722 9616
rect 8666 9560 8722 9596
rect 8108 9274 8164 9276
rect 8188 9274 8244 9276
rect 8268 9274 8324 9276
rect 8348 9274 8404 9276
rect 8108 9222 8154 9274
rect 8154 9222 8164 9274
rect 8188 9222 8218 9274
rect 8218 9222 8230 9274
rect 8230 9222 8244 9274
rect 8268 9222 8282 9274
rect 8282 9222 8294 9274
rect 8294 9222 8324 9274
rect 8348 9222 8358 9274
rect 8358 9222 8404 9274
rect 8108 9220 8164 9222
rect 8188 9220 8244 9222
rect 8268 9220 8324 9222
rect 8348 9220 8404 9222
rect 6734 8372 6736 8392
rect 6736 8372 6788 8392
rect 6788 8372 6790 8392
rect 6734 8336 6790 8372
rect 4256 7642 4312 7644
rect 4336 7642 4392 7644
rect 4416 7642 4472 7644
rect 4496 7642 4552 7644
rect 4256 7590 4302 7642
rect 4302 7590 4312 7642
rect 4336 7590 4366 7642
rect 4366 7590 4378 7642
rect 4378 7590 4392 7642
rect 4416 7590 4430 7642
rect 4430 7590 4442 7642
rect 4442 7590 4472 7642
rect 4496 7590 4506 7642
rect 4506 7590 4552 7642
rect 4256 7588 4312 7590
rect 4336 7588 4392 7590
rect 4416 7588 4472 7590
rect 4496 7588 4552 7590
rect 7010 7384 7066 7440
rect 4256 6554 4312 6556
rect 4336 6554 4392 6556
rect 4416 6554 4472 6556
rect 4496 6554 4552 6556
rect 4256 6502 4302 6554
rect 4302 6502 4312 6554
rect 4336 6502 4366 6554
rect 4366 6502 4378 6554
rect 4378 6502 4392 6554
rect 4416 6502 4430 6554
rect 4430 6502 4442 6554
rect 4442 6502 4472 6554
rect 4496 6502 4506 6554
rect 4506 6502 4552 6554
rect 4256 6500 4312 6502
rect 4336 6500 4392 6502
rect 4416 6500 4472 6502
rect 4496 6500 4552 6502
rect 7654 6840 7710 6896
rect 8108 8186 8164 8188
rect 8188 8186 8244 8188
rect 8268 8186 8324 8188
rect 8348 8186 8404 8188
rect 8108 8134 8154 8186
rect 8154 8134 8164 8186
rect 8188 8134 8218 8186
rect 8218 8134 8230 8186
rect 8230 8134 8244 8186
rect 8268 8134 8282 8186
rect 8282 8134 8294 8186
rect 8294 8134 8324 8186
rect 8348 8134 8358 8186
rect 8358 8134 8404 8186
rect 8108 8132 8164 8134
rect 8188 8132 8244 8134
rect 8268 8132 8324 8134
rect 8348 8132 8404 8134
rect 8108 7098 8164 7100
rect 8188 7098 8244 7100
rect 8268 7098 8324 7100
rect 8348 7098 8404 7100
rect 8108 7046 8154 7098
rect 8154 7046 8164 7098
rect 8188 7046 8218 7098
rect 8218 7046 8230 7098
rect 8230 7046 8244 7098
rect 8268 7046 8282 7098
rect 8282 7046 8294 7098
rect 8294 7046 8324 7098
rect 8348 7046 8358 7098
rect 8358 7046 8404 7098
rect 8108 7044 8164 7046
rect 8188 7044 8244 7046
rect 8268 7044 8324 7046
rect 8348 7044 8404 7046
rect 9770 9444 9826 9480
rect 9770 9424 9772 9444
rect 9772 9424 9824 9444
rect 9824 9424 9826 9444
rect 8850 7928 8906 7984
rect 9770 8356 9826 8392
rect 9770 8336 9772 8356
rect 9772 8336 9824 8356
rect 9824 8336 9826 8356
rect 10230 10648 10286 10704
rect 11702 12960 11758 13016
rect 12162 13912 12218 13968
rect 12070 13812 12072 13832
rect 12072 13812 12124 13832
rect 12124 13812 12126 13832
rect 12070 13776 12126 13812
rect 11961 13082 12017 13084
rect 12041 13082 12097 13084
rect 12121 13082 12177 13084
rect 12201 13082 12257 13084
rect 11961 13030 12007 13082
rect 12007 13030 12017 13082
rect 12041 13030 12071 13082
rect 12071 13030 12083 13082
rect 12083 13030 12097 13082
rect 12121 13030 12135 13082
rect 12135 13030 12147 13082
rect 12147 13030 12177 13082
rect 12201 13030 12211 13082
rect 12211 13030 12257 13082
rect 11961 13028 12017 13030
rect 12041 13028 12097 13030
rect 12121 13028 12177 13030
rect 12201 13028 12257 13030
rect 12622 16632 12678 16688
rect 12990 15952 13046 16008
rect 12438 13504 12494 13560
rect 12622 15136 12678 15192
rect 11961 11994 12017 11996
rect 12041 11994 12097 11996
rect 12121 11994 12177 11996
rect 12201 11994 12257 11996
rect 11961 11942 12007 11994
rect 12007 11942 12017 11994
rect 12041 11942 12071 11994
rect 12071 11942 12083 11994
rect 12083 11942 12097 11994
rect 12121 11942 12135 11994
rect 12135 11942 12147 11994
rect 12147 11942 12177 11994
rect 12201 11942 12211 11994
rect 12211 11942 12257 11994
rect 11961 11940 12017 11942
rect 12041 11940 12097 11942
rect 12121 11940 12177 11942
rect 12201 11940 12257 11942
rect 12990 14864 13046 14920
rect 12898 13640 12954 13696
rect 14094 16088 14150 16144
rect 13542 15952 13598 16008
rect 13634 15816 13690 15872
rect 13082 12280 13138 12336
rect 15813 19066 15869 19068
rect 15893 19066 15949 19068
rect 15973 19066 16029 19068
rect 16053 19066 16109 19068
rect 15813 19014 15859 19066
rect 15859 19014 15869 19066
rect 15893 19014 15923 19066
rect 15923 19014 15935 19066
rect 15935 19014 15949 19066
rect 15973 19014 15987 19066
rect 15987 19014 15999 19066
rect 15999 19014 16029 19066
rect 16053 19014 16063 19066
rect 16063 19014 16109 19066
rect 15813 19012 15869 19014
rect 15893 19012 15949 19014
rect 15973 19012 16029 19014
rect 16053 19012 16109 19014
rect 15813 17978 15869 17980
rect 15893 17978 15949 17980
rect 15973 17978 16029 17980
rect 16053 17978 16109 17980
rect 15813 17926 15859 17978
rect 15859 17926 15869 17978
rect 15893 17926 15923 17978
rect 15923 17926 15935 17978
rect 15935 17926 15949 17978
rect 15973 17926 15987 17978
rect 15987 17926 15999 17978
rect 15999 17926 16029 17978
rect 16053 17926 16063 17978
rect 16063 17926 16109 17978
rect 15813 17924 15869 17926
rect 15893 17924 15949 17926
rect 15973 17924 16029 17926
rect 16053 17924 16109 17926
rect 15813 16890 15869 16892
rect 15893 16890 15949 16892
rect 15973 16890 16029 16892
rect 16053 16890 16109 16892
rect 15813 16838 15859 16890
rect 15859 16838 15869 16890
rect 15893 16838 15923 16890
rect 15923 16838 15935 16890
rect 15935 16838 15949 16890
rect 15973 16838 15987 16890
rect 15987 16838 15999 16890
rect 15999 16838 16029 16890
rect 16053 16838 16063 16890
rect 16063 16838 16109 16890
rect 15813 16836 15869 16838
rect 15893 16836 15949 16838
rect 15973 16836 16029 16838
rect 16053 16836 16109 16838
rect 15014 13912 15070 13968
rect 15813 15802 15869 15804
rect 15893 15802 15949 15804
rect 15973 15802 16029 15804
rect 16053 15802 16109 15804
rect 15813 15750 15859 15802
rect 15859 15750 15869 15802
rect 15893 15750 15923 15802
rect 15923 15750 15935 15802
rect 15935 15750 15949 15802
rect 15973 15750 15987 15802
rect 15987 15750 15999 15802
rect 15999 15750 16029 15802
rect 16053 15750 16063 15802
rect 16063 15750 16109 15802
rect 15813 15748 15869 15750
rect 15893 15748 15949 15750
rect 15973 15748 16029 15750
rect 16053 15748 16109 15750
rect 15813 14714 15869 14716
rect 15893 14714 15949 14716
rect 15973 14714 16029 14716
rect 16053 14714 16109 14716
rect 15813 14662 15859 14714
rect 15859 14662 15869 14714
rect 15893 14662 15923 14714
rect 15923 14662 15935 14714
rect 15935 14662 15949 14714
rect 15973 14662 15987 14714
rect 15987 14662 15999 14714
rect 15999 14662 16029 14714
rect 16053 14662 16063 14714
rect 16063 14662 16109 14714
rect 15813 14660 15869 14662
rect 15893 14660 15949 14662
rect 15973 14660 16029 14662
rect 16053 14660 16109 14662
rect 15813 13626 15869 13628
rect 15893 13626 15949 13628
rect 15973 13626 16029 13628
rect 16053 13626 16109 13628
rect 15813 13574 15859 13626
rect 15859 13574 15869 13626
rect 15893 13574 15923 13626
rect 15923 13574 15935 13626
rect 15935 13574 15949 13626
rect 15973 13574 15987 13626
rect 15987 13574 15999 13626
rect 15999 13574 16029 13626
rect 16053 13574 16063 13626
rect 16063 13574 16109 13626
rect 15813 13572 15869 13574
rect 15893 13572 15949 13574
rect 15973 13572 16029 13574
rect 16053 13572 16109 13574
rect 14922 11636 14924 11656
rect 14924 11636 14976 11656
rect 14976 11636 14978 11656
rect 14922 11600 14978 11636
rect 15198 11736 15254 11792
rect 11961 10906 12017 10908
rect 12041 10906 12097 10908
rect 12121 10906 12177 10908
rect 12201 10906 12257 10908
rect 11961 10854 12007 10906
rect 12007 10854 12017 10906
rect 12041 10854 12071 10906
rect 12071 10854 12083 10906
rect 12083 10854 12097 10906
rect 12121 10854 12135 10906
rect 12135 10854 12147 10906
rect 12147 10854 12177 10906
rect 12201 10854 12211 10906
rect 12211 10854 12257 10906
rect 11961 10852 12017 10854
rect 12041 10852 12097 10854
rect 12121 10852 12177 10854
rect 12201 10852 12257 10854
rect 13266 10920 13322 10976
rect 14830 11056 14886 11112
rect 15813 12538 15869 12540
rect 15893 12538 15949 12540
rect 15973 12538 16029 12540
rect 16053 12538 16109 12540
rect 15813 12486 15859 12538
rect 15859 12486 15869 12538
rect 15893 12486 15923 12538
rect 15923 12486 15935 12538
rect 15935 12486 15949 12538
rect 15973 12486 15987 12538
rect 15987 12486 15999 12538
rect 15999 12486 16029 12538
rect 16053 12486 16063 12538
rect 16063 12486 16109 12538
rect 15813 12484 15869 12486
rect 15893 12484 15949 12486
rect 15973 12484 16029 12486
rect 16053 12484 16109 12486
rect 15382 11872 15438 11928
rect 15658 11756 15714 11792
rect 15658 11736 15660 11756
rect 15660 11736 15712 11756
rect 15712 11736 15714 11756
rect 15842 11736 15898 11792
rect 11961 9818 12017 9820
rect 12041 9818 12097 9820
rect 12121 9818 12177 9820
rect 12201 9818 12257 9820
rect 11961 9766 12007 9818
rect 12007 9766 12017 9818
rect 12041 9766 12071 9818
rect 12071 9766 12083 9818
rect 12083 9766 12097 9818
rect 12121 9766 12135 9818
rect 12135 9766 12147 9818
rect 12147 9766 12177 9818
rect 12201 9766 12211 9818
rect 12211 9766 12257 9818
rect 11961 9764 12017 9766
rect 12041 9764 12097 9766
rect 12121 9764 12177 9766
rect 12201 9764 12257 9766
rect 11334 9152 11390 9208
rect 9218 7284 9220 7304
rect 9220 7284 9272 7304
rect 9272 7284 9274 7304
rect 9218 7248 9274 7284
rect 9034 6180 9090 6216
rect 9034 6160 9036 6180
rect 9036 6160 9088 6180
rect 9088 6160 9090 6180
rect 8108 6010 8164 6012
rect 8188 6010 8244 6012
rect 8268 6010 8324 6012
rect 8348 6010 8404 6012
rect 8108 5958 8154 6010
rect 8154 5958 8164 6010
rect 8188 5958 8218 6010
rect 8218 5958 8230 6010
rect 8230 5958 8244 6010
rect 8268 5958 8282 6010
rect 8282 5958 8294 6010
rect 8294 5958 8324 6010
rect 8348 5958 8358 6010
rect 8358 5958 8404 6010
rect 8108 5956 8164 5958
rect 8188 5956 8244 5958
rect 8268 5956 8324 5958
rect 8348 5956 8404 5958
rect 4256 5466 4312 5468
rect 4336 5466 4392 5468
rect 4416 5466 4472 5468
rect 4496 5466 4552 5468
rect 4256 5414 4302 5466
rect 4302 5414 4312 5466
rect 4336 5414 4366 5466
rect 4366 5414 4378 5466
rect 4378 5414 4392 5466
rect 4416 5414 4430 5466
rect 4430 5414 4442 5466
rect 4442 5414 4472 5466
rect 4496 5414 4506 5466
rect 4506 5414 4552 5466
rect 4256 5412 4312 5414
rect 4336 5412 4392 5414
rect 4416 5412 4472 5414
rect 4496 5412 4552 5414
rect 8108 4922 8164 4924
rect 8188 4922 8244 4924
rect 8268 4922 8324 4924
rect 8348 4922 8404 4924
rect 8108 4870 8154 4922
rect 8154 4870 8164 4922
rect 8188 4870 8218 4922
rect 8218 4870 8230 4922
rect 8230 4870 8244 4922
rect 8268 4870 8282 4922
rect 8282 4870 8294 4922
rect 8294 4870 8324 4922
rect 8348 4870 8358 4922
rect 8358 4870 8404 4922
rect 8108 4868 8164 4870
rect 8188 4868 8244 4870
rect 8268 4868 8324 4870
rect 8348 4868 8404 4870
rect 4256 4378 4312 4380
rect 4336 4378 4392 4380
rect 4416 4378 4472 4380
rect 4496 4378 4552 4380
rect 4256 4326 4302 4378
rect 4302 4326 4312 4378
rect 4336 4326 4366 4378
rect 4366 4326 4378 4378
rect 4378 4326 4392 4378
rect 4416 4326 4430 4378
rect 4430 4326 4442 4378
rect 4442 4326 4472 4378
rect 4496 4326 4506 4378
rect 4506 4326 4552 4378
rect 4256 4324 4312 4326
rect 4336 4324 4392 4326
rect 4416 4324 4472 4326
rect 4496 4324 4552 4326
rect 8108 3834 8164 3836
rect 8188 3834 8244 3836
rect 8268 3834 8324 3836
rect 8348 3834 8404 3836
rect 8108 3782 8154 3834
rect 8154 3782 8164 3834
rect 8188 3782 8218 3834
rect 8218 3782 8230 3834
rect 8230 3782 8244 3834
rect 8268 3782 8282 3834
rect 8282 3782 8294 3834
rect 8294 3782 8324 3834
rect 8348 3782 8358 3834
rect 8358 3782 8404 3834
rect 8108 3780 8164 3782
rect 8188 3780 8244 3782
rect 8268 3780 8324 3782
rect 8348 3780 8404 3782
rect 4256 3290 4312 3292
rect 4336 3290 4392 3292
rect 4416 3290 4472 3292
rect 4496 3290 4552 3292
rect 4256 3238 4302 3290
rect 4302 3238 4312 3290
rect 4336 3238 4366 3290
rect 4366 3238 4378 3290
rect 4378 3238 4392 3290
rect 4416 3238 4430 3290
rect 4430 3238 4442 3290
rect 4442 3238 4472 3290
rect 4496 3238 4506 3290
rect 4506 3238 4552 3290
rect 4256 3236 4312 3238
rect 4336 3236 4392 3238
rect 4416 3236 4472 3238
rect 4496 3236 4552 3238
rect 8108 2746 8164 2748
rect 8188 2746 8244 2748
rect 8268 2746 8324 2748
rect 8348 2746 8404 2748
rect 8108 2694 8154 2746
rect 8154 2694 8164 2746
rect 8188 2694 8218 2746
rect 8218 2694 8230 2746
rect 8230 2694 8244 2746
rect 8268 2694 8282 2746
rect 8282 2694 8294 2746
rect 8294 2694 8324 2746
rect 8348 2694 8358 2746
rect 8358 2694 8404 2746
rect 8108 2692 8164 2694
rect 8188 2692 8244 2694
rect 8268 2692 8324 2694
rect 8348 2692 8404 2694
rect 4256 2202 4312 2204
rect 4336 2202 4392 2204
rect 4416 2202 4472 2204
rect 4496 2202 4552 2204
rect 4256 2150 4302 2202
rect 4302 2150 4312 2202
rect 4336 2150 4366 2202
rect 4366 2150 4378 2202
rect 4378 2150 4392 2202
rect 4416 2150 4430 2202
rect 4430 2150 4442 2202
rect 4442 2150 4472 2202
rect 4496 2150 4506 2202
rect 4506 2150 4552 2202
rect 4256 2148 4312 2150
rect 4336 2148 4392 2150
rect 4416 2148 4472 2150
rect 4496 2148 4552 2150
rect 8108 1658 8164 1660
rect 8188 1658 8244 1660
rect 8268 1658 8324 1660
rect 8348 1658 8404 1660
rect 8108 1606 8154 1658
rect 8154 1606 8164 1658
rect 8188 1606 8218 1658
rect 8218 1606 8230 1658
rect 8230 1606 8244 1658
rect 8268 1606 8282 1658
rect 8282 1606 8294 1658
rect 8294 1606 8324 1658
rect 8348 1606 8358 1658
rect 8358 1606 8404 1658
rect 8108 1604 8164 1606
rect 8188 1604 8244 1606
rect 8268 1604 8324 1606
rect 8348 1604 8404 1606
rect 4256 1114 4312 1116
rect 4336 1114 4392 1116
rect 4416 1114 4472 1116
rect 4496 1114 4552 1116
rect 4256 1062 4302 1114
rect 4302 1062 4312 1114
rect 4336 1062 4366 1114
rect 4366 1062 4378 1114
rect 4378 1062 4392 1114
rect 4416 1062 4430 1114
rect 4430 1062 4442 1114
rect 4442 1062 4472 1114
rect 4496 1062 4506 1114
rect 4506 1062 4552 1114
rect 4256 1060 4312 1062
rect 4336 1060 4392 1062
rect 4416 1060 4472 1062
rect 4496 1060 4552 1062
rect 9586 7248 9642 7304
rect 11961 8730 12017 8732
rect 12041 8730 12097 8732
rect 12121 8730 12177 8732
rect 12201 8730 12257 8732
rect 11961 8678 12007 8730
rect 12007 8678 12017 8730
rect 12041 8678 12071 8730
rect 12071 8678 12083 8730
rect 12083 8678 12097 8730
rect 12121 8678 12135 8730
rect 12135 8678 12147 8730
rect 12147 8678 12177 8730
rect 12201 8678 12211 8730
rect 12211 8678 12257 8730
rect 11961 8676 12017 8678
rect 12041 8676 12097 8678
rect 12121 8676 12177 8678
rect 12201 8676 12257 8678
rect 12714 9036 12770 9072
rect 12714 9016 12716 9036
rect 12716 9016 12768 9036
rect 12768 9016 12770 9036
rect 10138 7384 10194 7440
rect 10322 6840 10378 6896
rect 9770 6160 9826 6216
rect 9310 4664 9366 4720
rect 10690 4684 10746 4720
rect 10690 4664 10692 4684
rect 10692 4664 10744 4684
rect 10744 4664 10746 4684
rect 8108 570 8164 572
rect 8188 570 8244 572
rect 8268 570 8324 572
rect 8348 570 8404 572
rect 8108 518 8154 570
rect 8154 518 8164 570
rect 8188 518 8218 570
rect 8218 518 8230 570
rect 8230 518 8244 570
rect 8268 518 8282 570
rect 8282 518 8294 570
rect 8294 518 8324 570
rect 8348 518 8358 570
rect 8358 518 8404 570
rect 8108 516 8164 518
rect 8188 516 8244 518
rect 8268 516 8324 518
rect 8348 516 8404 518
rect 13450 9152 13506 9208
rect 15813 11450 15869 11452
rect 15893 11450 15949 11452
rect 15973 11450 16029 11452
rect 16053 11450 16109 11452
rect 15813 11398 15859 11450
rect 15859 11398 15869 11450
rect 15893 11398 15923 11450
rect 15923 11398 15935 11450
rect 15935 11398 15949 11450
rect 15973 11398 15987 11450
rect 15987 11398 15999 11450
rect 15999 11398 16029 11450
rect 16053 11398 16063 11450
rect 16063 11398 16109 11450
rect 15813 11396 15869 11398
rect 15893 11396 15949 11398
rect 15973 11396 16029 11398
rect 16053 11396 16109 11398
rect 16118 11212 16174 11248
rect 16118 11192 16120 11212
rect 16120 11192 16172 11212
rect 16172 11192 16174 11212
rect 15658 10376 15714 10432
rect 15813 10362 15869 10364
rect 15893 10362 15949 10364
rect 15973 10362 16029 10364
rect 16053 10362 16109 10364
rect 15813 10310 15859 10362
rect 15859 10310 15869 10362
rect 15893 10310 15923 10362
rect 15923 10310 15935 10362
rect 15935 10310 15949 10362
rect 15973 10310 15987 10362
rect 15987 10310 15999 10362
rect 15999 10310 16029 10362
rect 16053 10310 16063 10362
rect 16063 10310 16109 10362
rect 15813 10308 15869 10310
rect 15893 10308 15949 10310
rect 15973 10308 16029 10310
rect 16053 10308 16109 10310
rect 15474 9968 15530 10024
rect 11961 7642 12017 7644
rect 12041 7642 12097 7644
rect 12121 7642 12177 7644
rect 12201 7642 12257 7644
rect 11961 7590 12007 7642
rect 12007 7590 12017 7642
rect 12041 7590 12071 7642
rect 12071 7590 12083 7642
rect 12083 7590 12097 7642
rect 12121 7590 12135 7642
rect 12135 7590 12147 7642
rect 12147 7590 12177 7642
rect 12201 7590 12211 7642
rect 12211 7590 12257 7642
rect 11961 7588 12017 7590
rect 12041 7588 12097 7590
rect 12121 7588 12177 7590
rect 12201 7588 12257 7590
rect 11518 6976 11574 7032
rect 11961 6554 12017 6556
rect 12041 6554 12097 6556
rect 12121 6554 12177 6556
rect 12201 6554 12257 6556
rect 11961 6502 12007 6554
rect 12007 6502 12017 6554
rect 12041 6502 12071 6554
rect 12071 6502 12083 6554
rect 12083 6502 12097 6554
rect 12121 6502 12135 6554
rect 12135 6502 12147 6554
rect 12147 6502 12177 6554
rect 12201 6502 12211 6554
rect 12211 6502 12257 6554
rect 11961 6500 12017 6502
rect 12041 6500 12097 6502
rect 12121 6500 12177 6502
rect 12201 6500 12257 6502
rect 11961 5466 12017 5468
rect 12041 5466 12097 5468
rect 12121 5466 12177 5468
rect 12201 5466 12257 5468
rect 11961 5414 12007 5466
rect 12007 5414 12017 5466
rect 12041 5414 12071 5466
rect 12071 5414 12083 5466
rect 12083 5414 12097 5466
rect 12121 5414 12135 5466
rect 12135 5414 12147 5466
rect 12147 5414 12177 5466
rect 12201 5414 12211 5466
rect 12211 5414 12257 5466
rect 11961 5412 12017 5414
rect 12041 5412 12097 5414
rect 12121 5412 12177 5414
rect 12201 5412 12257 5414
rect 11961 4378 12017 4380
rect 12041 4378 12097 4380
rect 12121 4378 12177 4380
rect 12201 4378 12257 4380
rect 11961 4326 12007 4378
rect 12007 4326 12017 4378
rect 12041 4326 12071 4378
rect 12071 4326 12083 4378
rect 12083 4326 12097 4378
rect 12121 4326 12135 4378
rect 12135 4326 12147 4378
rect 12147 4326 12177 4378
rect 12201 4326 12211 4378
rect 12211 4326 12257 4378
rect 11961 4324 12017 4326
rect 12041 4324 12097 4326
rect 12121 4324 12177 4326
rect 12201 4324 12257 4326
rect 11961 3290 12017 3292
rect 12041 3290 12097 3292
rect 12121 3290 12177 3292
rect 12201 3290 12257 3292
rect 11961 3238 12007 3290
rect 12007 3238 12017 3290
rect 12041 3238 12071 3290
rect 12071 3238 12083 3290
rect 12083 3238 12097 3290
rect 12121 3238 12135 3290
rect 12135 3238 12147 3290
rect 12147 3238 12177 3290
rect 12201 3238 12211 3290
rect 12211 3238 12257 3290
rect 11961 3236 12017 3238
rect 12041 3236 12097 3238
rect 12121 3236 12177 3238
rect 12201 3236 12257 3238
rect 11961 2202 12017 2204
rect 12041 2202 12097 2204
rect 12121 2202 12177 2204
rect 12201 2202 12257 2204
rect 11961 2150 12007 2202
rect 12007 2150 12017 2202
rect 12041 2150 12071 2202
rect 12071 2150 12083 2202
rect 12083 2150 12097 2202
rect 12121 2150 12135 2202
rect 12135 2150 12147 2202
rect 12147 2150 12177 2202
rect 12201 2150 12211 2202
rect 12211 2150 12257 2202
rect 11961 2148 12017 2150
rect 12041 2148 12097 2150
rect 12121 2148 12177 2150
rect 12201 2148 12257 2150
rect 11961 1114 12017 1116
rect 12041 1114 12097 1116
rect 12121 1114 12177 1116
rect 12201 1114 12257 1116
rect 11961 1062 12007 1114
rect 12007 1062 12017 1114
rect 12041 1062 12071 1114
rect 12071 1062 12083 1114
rect 12083 1062 12097 1114
rect 12121 1062 12135 1114
rect 12135 1062 12147 1114
rect 12147 1062 12177 1114
rect 12201 1062 12211 1114
rect 12211 1062 12257 1114
rect 11961 1060 12017 1062
rect 12041 1060 12097 1062
rect 12121 1060 12177 1062
rect 12201 1060 12257 1062
rect 14554 5480 14610 5536
rect 15566 9580 15622 9616
rect 15566 9560 15568 9580
rect 15568 9560 15620 9580
rect 15620 9560 15622 9580
rect 15934 10104 15990 10160
rect 15842 10004 15844 10024
rect 15844 10004 15896 10024
rect 15896 10004 15898 10024
rect 15842 9968 15898 10004
rect 16486 11056 16542 11112
rect 17130 11872 17186 11928
rect 18602 15036 18604 15056
rect 18604 15036 18656 15056
rect 18656 15036 18658 15056
rect 18602 15000 18658 15036
rect 18510 12280 18566 12336
rect 15813 9274 15869 9276
rect 15893 9274 15949 9276
rect 15973 9274 16029 9276
rect 16053 9274 16109 9276
rect 15813 9222 15859 9274
rect 15859 9222 15869 9274
rect 15893 9222 15923 9274
rect 15923 9222 15935 9274
rect 15935 9222 15949 9274
rect 15973 9222 15987 9274
rect 15987 9222 15999 9274
rect 15999 9222 16029 9274
rect 16053 9222 16063 9274
rect 16063 9222 16109 9274
rect 15813 9220 15869 9222
rect 15893 9220 15949 9222
rect 15973 9220 16029 9222
rect 16053 9220 16109 9222
rect 18234 11736 18290 11792
rect 15198 8336 15254 8392
rect 15813 8186 15869 8188
rect 15893 8186 15949 8188
rect 15973 8186 16029 8188
rect 16053 8186 16109 8188
rect 15813 8134 15859 8186
rect 15859 8134 15869 8186
rect 15893 8134 15923 8186
rect 15923 8134 15935 8186
rect 15935 8134 15949 8186
rect 15973 8134 15987 8186
rect 15987 8134 15999 8186
rect 15999 8134 16029 8186
rect 16053 8134 16063 8186
rect 16063 8134 16109 8186
rect 15813 8132 15869 8134
rect 15893 8132 15949 8134
rect 15973 8132 16029 8134
rect 16053 8132 16109 8134
rect 14830 7148 14832 7168
rect 14832 7148 14884 7168
rect 14884 7148 14886 7168
rect 14830 7112 14886 7148
rect 15474 7112 15530 7168
rect 15382 6840 15438 6896
rect 15106 5480 15162 5536
rect 15014 5344 15070 5400
rect 14922 4936 14978 4992
rect 15813 7098 15869 7100
rect 15893 7098 15949 7100
rect 15973 7098 16029 7100
rect 16053 7098 16109 7100
rect 15813 7046 15859 7098
rect 15859 7046 15869 7098
rect 15893 7046 15923 7098
rect 15923 7046 15935 7098
rect 15935 7046 15949 7098
rect 15973 7046 15987 7098
rect 15987 7046 15999 7098
rect 15999 7046 16029 7098
rect 16053 7046 16063 7098
rect 16063 7046 16109 7098
rect 15813 7044 15869 7046
rect 15893 7044 15949 7046
rect 15973 7044 16029 7046
rect 16053 7044 16109 7046
rect 15813 6010 15869 6012
rect 15893 6010 15949 6012
rect 15973 6010 16029 6012
rect 16053 6010 16109 6012
rect 15813 5958 15859 6010
rect 15859 5958 15869 6010
rect 15893 5958 15923 6010
rect 15923 5958 15935 6010
rect 15935 5958 15949 6010
rect 15973 5958 15987 6010
rect 15987 5958 15999 6010
rect 15999 5958 16029 6010
rect 16053 5958 16063 6010
rect 16063 5958 16109 6010
rect 15813 5956 15869 5958
rect 15893 5956 15949 5958
rect 15973 5956 16029 5958
rect 16053 5956 16109 5958
rect 15813 4922 15869 4924
rect 15893 4922 15949 4924
rect 15973 4922 16029 4924
rect 16053 4922 16109 4924
rect 15813 4870 15859 4922
rect 15859 4870 15869 4922
rect 15893 4870 15923 4922
rect 15923 4870 15935 4922
rect 15935 4870 15949 4922
rect 15973 4870 15987 4922
rect 15987 4870 15999 4922
rect 15999 4870 16029 4922
rect 16053 4870 16063 4922
rect 16063 4870 16109 4922
rect 15813 4868 15869 4870
rect 15893 4868 15949 4870
rect 15973 4868 16029 4870
rect 16053 4868 16109 4870
rect 15813 3834 15869 3836
rect 15893 3834 15949 3836
rect 15973 3834 16029 3836
rect 16053 3834 16109 3836
rect 15813 3782 15859 3834
rect 15859 3782 15869 3834
rect 15893 3782 15923 3834
rect 15923 3782 15935 3834
rect 15935 3782 15949 3834
rect 15973 3782 15987 3834
rect 15987 3782 15999 3834
rect 15999 3782 16029 3834
rect 16053 3782 16063 3834
rect 16063 3782 16109 3834
rect 15813 3780 15869 3782
rect 15893 3780 15949 3782
rect 15973 3780 16029 3782
rect 16053 3780 16109 3782
rect 15813 2746 15869 2748
rect 15893 2746 15949 2748
rect 15973 2746 16029 2748
rect 16053 2746 16109 2748
rect 15813 2694 15859 2746
rect 15859 2694 15869 2746
rect 15893 2694 15923 2746
rect 15923 2694 15935 2746
rect 15935 2694 15949 2746
rect 15973 2694 15987 2746
rect 15987 2694 15999 2746
rect 15999 2694 16029 2746
rect 16053 2694 16063 2746
rect 16063 2694 16109 2746
rect 15813 2692 15869 2694
rect 15893 2692 15949 2694
rect 15973 2692 16029 2694
rect 16053 2692 16109 2694
rect 15813 1658 15869 1660
rect 15893 1658 15949 1660
rect 15973 1658 16029 1660
rect 16053 1658 16109 1660
rect 15813 1606 15859 1658
rect 15859 1606 15869 1658
rect 15893 1606 15923 1658
rect 15923 1606 15935 1658
rect 15935 1606 15949 1658
rect 15973 1606 15987 1658
rect 15987 1606 15999 1658
rect 15999 1606 16029 1658
rect 16053 1606 16063 1658
rect 16063 1606 16109 1658
rect 15813 1604 15869 1606
rect 15893 1604 15949 1606
rect 15973 1604 16029 1606
rect 16053 1604 16109 1606
rect 15813 570 15869 572
rect 15893 570 15949 572
rect 15973 570 16029 572
rect 16053 570 16109 572
rect 15813 518 15859 570
rect 15859 518 15869 570
rect 15893 518 15923 570
rect 15923 518 15935 570
rect 15935 518 15949 570
rect 15973 518 15987 570
rect 15987 518 15999 570
rect 15999 518 16029 570
rect 16053 518 16063 570
rect 16063 518 16109 570
rect 15813 516 15869 518
rect 15893 516 15949 518
rect 15973 516 16029 518
rect 16053 516 16109 518
rect 17958 9596 17960 9616
rect 17960 9596 18012 9616
rect 18012 9596 18014 9616
rect 17958 9560 18014 9596
rect 17774 9052 17776 9072
rect 17776 9052 17828 9072
rect 17828 9052 17830 9072
rect 17774 9016 17830 9052
rect 19666 18522 19722 18524
rect 19746 18522 19802 18524
rect 19826 18522 19882 18524
rect 19906 18522 19962 18524
rect 19666 18470 19712 18522
rect 19712 18470 19722 18522
rect 19746 18470 19776 18522
rect 19776 18470 19788 18522
rect 19788 18470 19802 18522
rect 19826 18470 19840 18522
rect 19840 18470 19852 18522
rect 19852 18470 19882 18522
rect 19906 18470 19916 18522
rect 19916 18470 19962 18522
rect 19666 18468 19722 18470
rect 19746 18468 19802 18470
rect 19826 18468 19882 18470
rect 19906 18468 19962 18470
rect 19666 17434 19722 17436
rect 19746 17434 19802 17436
rect 19826 17434 19882 17436
rect 19906 17434 19962 17436
rect 19666 17382 19712 17434
rect 19712 17382 19722 17434
rect 19746 17382 19776 17434
rect 19776 17382 19788 17434
rect 19788 17382 19802 17434
rect 19826 17382 19840 17434
rect 19840 17382 19852 17434
rect 19852 17382 19882 17434
rect 19906 17382 19916 17434
rect 19916 17382 19962 17434
rect 19666 17380 19722 17382
rect 19746 17380 19802 17382
rect 19826 17380 19882 17382
rect 19906 17380 19962 17382
rect 19338 17040 19394 17096
rect 20350 16904 20406 16960
rect 20350 16768 20406 16824
rect 19666 16346 19722 16348
rect 19746 16346 19802 16348
rect 19826 16346 19882 16348
rect 19906 16346 19962 16348
rect 19666 16294 19712 16346
rect 19712 16294 19722 16346
rect 19746 16294 19776 16346
rect 19776 16294 19788 16346
rect 19788 16294 19802 16346
rect 19826 16294 19840 16346
rect 19840 16294 19852 16346
rect 19852 16294 19882 16346
rect 19906 16294 19916 16346
rect 19916 16294 19962 16346
rect 19666 16292 19722 16294
rect 19746 16292 19802 16294
rect 19826 16292 19882 16294
rect 19906 16292 19962 16294
rect 19666 15258 19722 15260
rect 19746 15258 19802 15260
rect 19826 15258 19882 15260
rect 19906 15258 19962 15260
rect 19666 15206 19712 15258
rect 19712 15206 19722 15258
rect 19746 15206 19776 15258
rect 19776 15206 19788 15258
rect 19788 15206 19802 15258
rect 19826 15206 19840 15258
rect 19840 15206 19852 15258
rect 19852 15206 19882 15258
rect 19906 15206 19916 15258
rect 19916 15206 19962 15258
rect 19666 15204 19722 15206
rect 19746 15204 19802 15206
rect 19826 15204 19882 15206
rect 19906 15204 19962 15206
rect 19666 14170 19722 14172
rect 19746 14170 19802 14172
rect 19826 14170 19882 14172
rect 19906 14170 19962 14172
rect 19666 14118 19712 14170
rect 19712 14118 19722 14170
rect 19746 14118 19776 14170
rect 19776 14118 19788 14170
rect 19788 14118 19802 14170
rect 19826 14118 19840 14170
rect 19840 14118 19852 14170
rect 19852 14118 19882 14170
rect 19906 14118 19916 14170
rect 19916 14118 19962 14170
rect 19666 14116 19722 14118
rect 19746 14116 19802 14118
rect 19826 14116 19882 14118
rect 19906 14116 19962 14118
rect 19062 13640 19118 13696
rect 19666 13082 19722 13084
rect 19746 13082 19802 13084
rect 19826 13082 19882 13084
rect 19906 13082 19962 13084
rect 19666 13030 19712 13082
rect 19712 13030 19722 13082
rect 19746 13030 19776 13082
rect 19776 13030 19788 13082
rect 19788 13030 19802 13082
rect 19826 13030 19840 13082
rect 19840 13030 19852 13082
rect 19852 13030 19882 13082
rect 19906 13030 19916 13082
rect 19916 13030 19962 13082
rect 19666 13028 19722 13030
rect 19746 13028 19802 13030
rect 19826 13028 19882 13030
rect 19906 13028 19962 13030
rect 20442 16224 20498 16280
rect 21546 17040 21602 17096
rect 21178 16496 21234 16552
rect 20442 13776 20498 13832
rect 21454 16496 21510 16552
rect 20902 15272 20958 15328
rect 21362 15816 21418 15872
rect 21178 13096 21234 13152
rect 21730 16904 21786 16960
rect 21454 15136 21510 15192
rect 21638 15816 21694 15872
rect 21546 14592 21602 14648
rect 22006 16904 22062 16960
rect 22282 16224 22338 16280
rect 21822 15680 21878 15736
rect 22374 16108 22430 16144
rect 22374 16088 22376 16108
rect 22376 16088 22428 16108
rect 22428 16088 22430 16108
rect 22834 16904 22890 16960
rect 22926 16768 22982 16824
rect 22834 16360 22890 16416
rect 21914 15564 21970 15600
rect 21914 15544 21916 15564
rect 21916 15544 21968 15564
rect 21968 15544 21970 15564
rect 21638 13912 21694 13968
rect 19338 11736 19394 11792
rect 19430 11600 19486 11656
rect 19666 11994 19722 11996
rect 19746 11994 19802 11996
rect 19826 11994 19882 11996
rect 19906 11994 19962 11996
rect 19666 11942 19712 11994
rect 19712 11942 19722 11994
rect 19746 11942 19776 11994
rect 19776 11942 19788 11994
rect 19788 11942 19802 11994
rect 19826 11942 19840 11994
rect 19840 11942 19852 11994
rect 19852 11942 19882 11994
rect 19906 11942 19916 11994
rect 19916 11942 19962 11994
rect 19666 11940 19722 11942
rect 19746 11940 19802 11942
rect 19826 11940 19882 11942
rect 19906 11940 19962 11942
rect 20350 12008 20406 12064
rect 19666 10906 19722 10908
rect 19746 10906 19802 10908
rect 19826 10906 19882 10908
rect 19906 10906 19962 10908
rect 19666 10854 19712 10906
rect 19712 10854 19722 10906
rect 19746 10854 19776 10906
rect 19776 10854 19788 10906
rect 19788 10854 19802 10906
rect 19826 10854 19840 10906
rect 19840 10854 19852 10906
rect 19852 10854 19882 10906
rect 19906 10854 19916 10906
rect 19916 10854 19962 10906
rect 19666 10852 19722 10854
rect 19746 10852 19802 10854
rect 19826 10852 19882 10854
rect 19906 10852 19962 10854
rect 22558 15952 22614 16008
rect 22190 15428 22246 15464
rect 22190 15408 22192 15428
rect 22192 15408 22244 15428
rect 22244 15408 22246 15428
rect 22006 14320 22062 14376
rect 22742 14864 22798 14920
rect 22466 14456 22522 14512
rect 23518 19066 23574 19068
rect 23598 19066 23654 19068
rect 23678 19066 23734 19068
rect 23758 19066 23814 19068
rect 23518 19014 23564 19066
rect 23564 19014 23574 19066
rect 23598 19014 23628 19066
rect 23628 19014 23640 19066
rect 23640 19014 23654 19066
rect 23678 19014 23692 19066
rect 23692 19014 23704 19066
rect 23704 19014 23734 19066
rect 23758 19014 23768 19066
rect 23768 19014 23814 19066
rect 23518 19012 23574 19014
rect 23598 19012 23654 19014
rect 23678 19012 23734 19014
rect 23758 19012 23814 19014
rect 23518 17978 23574 17980
rect 23598 17978 23654 17980
rect 23678 17978 23734 17980
rect 23758 17978 23814 17980
rect 23518 17926 23564 17978
rect 23564 17926 23574 17978
rect 23598 17926 23628 17978
rect 23628 17926 23640 17978
rect 23640 17926 23654 17978
rect 23678 17926 23692 17978
rect 23692 17926 23704 17978
rect 23704 17926 23734 17978
rect 23758 17926 23768 17978
rect 23768 17926 23814 17978
rect 23518 17924 23574 17926
rect 23598 17924 23654 17926
rect 23678 17924 23734 17926
rect 23758 17924 23814 17926
rect 23518 16890 23574 16892
rect 23598 16890 23654 16892
rect 23678 16890 23734 16892
rect 23758 16890 23814 16892
rect 23518 16838 23564 16890
rect 23564 16838 23574 16890
rect 23598 16838 23628 16890
rect 23628 16838 23640 16890
rect 23640 16838 23654 16890
rect 23678 16838 23692 16890
rect 23692 16838 23704 16890
rect 23704 16838 23734 16890
rect 23758 16838 23768 16890
rect 23768 16838 23814 16890
rect 23518 16836 23574 16838
rect 23598 16836 23654 16838
rect 23678 16836 23734 16838
rect 23758 16836 23814 16838
rect 23294 16244 23350 16280
rect 23294 16224 23296 16244
rect 23296 16224 23348 16244
rect 23348 16224 23350 16244
rect 23202 14592 23258 14648
rect 23662 15952 23718 16008
rect 23846 15952 23902 16008
rect 23518 15802 23574 15804
rect 23598 15802 23654 15804
rect 23678 15802 23734 15804
rect 23758 15802 23814 15804
rect 23518 15750 23564 15802
rect 23564 15750 23574 15802
rect 23598 15750 23628 15802
rect 23628 15750 23640 15802
rect 23640 15750 23654 15802
rect 23678 15750 23692 15802
rect 23692 15750 23704 15802
rect 23704 15750 23734 15802
rect 23758 15750 23768 15802
rect 23768 15750 23814 15802
rect 23518 15748 23574 15750
rect 23598 15748 23654 15750
rect 23678 15748 23734 15750
rect 23758 15748 23814 15750
rect 23846 15444 23848 15464
rect 23848 15444 23900 15464
rect 23900 15444 23902 15464
rect 23846 15408 23902 15444
rect 23846 15272 23902 15328
rect 23518 14714 23574 14716
rect 23598 14714 23654 14716
rect 23678 14714 23734 14716
rect 23758 14714 23814 14716
rect 23518 14662 23564 14714
rect 23564 14662 23574 14714
rect 23598 14662 23628 14714
rect 23628 14662 23640 14714
rect 23640 14662 23654 14714
rect 23678 14662 23692 14714
rect 23692 14662 23704 14714
rect 23704 14662 23734 14714
rect 23758 14662 23768 14714
rect 23768 14662 23814 14714
rect 23518 14660 23574 14662
rect 23598 14660 23654 14662
rect 23678 14660 23734 14662
rect 23758 14660 23814 14662
rect 23294 14048 23350 14104
rect 24214 17040 24270 17096
rect 24030 16108 24086 16144
rect 24030 16088 24032 16108
rect 24032 16088 24084 16108
rect 24084 16088 24086 16108
rect 24306 15408 24362 15464
rect 23846 13776 23902 13832
rect 23518 13626 23574 13628
rect 23598 13626 23654 13628
rect 23678 13626 23734 13628
rect 23758 13626 23814 13628
rect 23518 13574 23564 13626
rect 23564 13574 23574 13626
rect 23598 13574 23628 13626
rect 23628 13574 23640 13626
rect 23640 13574 23654 13626
rect 23678 13574 23692 13626
rect 23692 13574 23704 13626
rect 23704 13574 23734 13626
rect 23758 13574 23768 13626
rect 23768 13574 23814 13626
rect 23518 13572 23574 13574
rect 23598 13572 23654 13574
rect 23678 13572 23734 13574
rect 23758 13572 23814 13574
rect 23294 13232 23350 13288
rect 24858 16360 24914 16416
rect 25042 16224 25098 16280
rect 24674 15136 24730 15192
rect 24582 15000 24638 15056
rect 24766 14900 24768 14920
rect 24768 14900 24820 14920
rect 24820 14900 24822 14920
rect 24766 14864 24822 14900
rect 24490 14320 24546 14376
rect 24490 13640 24546 13696
rect 24950 14184 25006 14240
rect 24674 13912 24730 13968
rect 24582 13504 24638 13560
rect 24490 13096 24546 13152
rect 23662 12688 23718 12744
rect 19666 9818 19722 9820
rect 19746 9818 19802 9820
rect 19826 9818 19882 9820
rect 19906 9818 19962 9820
rect 19666 9766 19712 9818
rect 19712 9766 19722 9818
rect 19746 9766 19776 9818
rect 19776 9766 19788 9818
rect 19788 9766 19802 9818
rect 19826 9766 19840 9818
rect 19840 9766 19852 9818
rect 19852 9766 19882 9818
rect 19906 9766 19916 9818
rect 19916 9766 19962 9818
rect 19666 9764 19722 9766
rect 19746 9764 19802 9766
rect 19826 9764 19882 9766
rect 19906 9764 19962 9766
rect 21362 9560 21418 9616
rect 19338 9016 19394 9072
rect 19666 8730 19722 8732
rect 19746 8730 19802 8732
rect 19826 8730 19882 8732
rect 19906 8730 19962 8732
rect 19666 8678 19712 8730
rect 19712 8678 19722 8730
rect 19746 8678 19776 8730
rect 19776 8678 19788 8730
rect 19788 8678 19802 8730
rect 19826 8678 19840 8730
rect 19840 8678 19852 8730
rect 19852 8678 19882 8730
rect 19906 8678 19916 8730
rect 19916 8678 19962 8730
rect 19666 8676 19722 8678
rect 19746 8676 19802 8678
rect 19826 8676 19882 8678
rect 19906 8676 19962 8678
rect 18878 6196 18880 6216
rect 18880 6196 18932 6216
rect 18932 6196 18934 6216
rect 18878 6160 18934 6196
rect 19666 7642 19722 7644
rect 19746 7642 19802 7644
rect 19826 7642 19882 7644
rect 19906 7642 19962 7644
rect 19666 7590 19712 7642
rect 19712 7590 19722 7642
rect 19746 7590 19776 7642
rect 19776 7590 19788 7642
rect 19788 7590 19802 7642
rect 19826 7590 19840 7642
rect 19840 7590 19852 7642
rect 19852 7590 19882 7642
rect 19906 7590 19916 7642
rect 19916 7590 19962 7642
rect 19666 7588 19722 7590
rect 19746 7588 19802 7590
rect 19826 7588 19882 7590
rect 19906 7588 19962 7590
rect 19706 7248 19762 7304
rect 19666 6554 19722 6556
rect 19746 6554 19802 6556
rect 19826 6554 19882 6556
rect 19906 6554 19962 6556
rect 19666 6502 19712 6554
rect 19712 6502 19722 6554
rect 19746 6502 19776 6554
rect 19776 6502 19788 6554
rect 19788 6502 19802 6554
rect 19826 6502 19840 6554
rect 19840 6502 19852 6554
rect 19852 6502 19882 6554
rect 19906 6502 19916 6554
rect 19916 6502 19962 6554
rect 19666 6500 19722 6502
rect 19746 6500 19802 6502
rect 19826 6500 19882 6502
rect 19906 6500 19962 6502
rect 19246 6160 19302 6216
rect 20166 8336 20222 8392
rect 20166 7284 20168 7304
rect 20168 7284 20220 7304
rect 20220 7284 20222 7304
rect 20166 7248 20222 7284
rect 19062 5636 19118 5672
rect 19062 5616 19064 5636
rect 19064 5616 19116 5636
rect 19116 5616 19118 5636
rect 8298 312 8354 368
rect 20074 5888 20130 5944
rect 19666 5466 19722 5468
rect 19746 5466 19802 5468
rect 19826 5466 19882 5468
rect 19906 5466 19962 5468
rect 19666 5414 19712 5466
rect 19712 5414 19722 5466
rect 19746 5414 19776 5466
rect 19776 5414 19788 5466
rect 19788 5414 19802 5466
rect 19826 5414 19840 5466
rect 19840 5414 19852 5466
rect 19852 5414 19882 5466
rect 19906 5414 19916 5466
rect 19916 5414 19962 5466
rect 19666 5412 19722 5414
rect 19746 5412 19802 5414
rect 19826 5412 19882 5414
rect 19906 5412 19962 5414
rect 20350 5772 20406 5808
rect 23518 12538 23574 12540
rect 23598 12538 23654 12540
rect 23678 12538 23734 12540
rect 23758 12538 23814 12540
rect 23518 12486 23564 12538
rect 23564 12486 23574 12538
rect 23598 12486 23628 12538
rect 23628 12486 23640 12538
rect 23640 12486 23654 12538
rect 23678 12486 23692 12538
rect 23692 12486 23704 12538
rect 23704 12486 23734 12538
rect 23758 12486 23768 12538
rect 23768 12486 23814 12538
rect 23518 12484 23574 12486
rect 23598 12484 23654 12486
rect 23678 12484 23734 12486
rect 23758 12484 23814 12486
rect 23294 11736 23350 11792
rect 23518 11450 23574 11452
rect 23598 11450 23654 11452
rect 23678 11450 23734 11452
rect 23758 11450 23814 11452
rect 23518 11398 23564 11450
rect 23564 11398 23574 11450
rect 23598 11398 23628 11450
rect 23628 11398 23640 11450
rect 23640 11398 23654 11450
rect 23678 11398 23692 11450
rect 23692 11398 23704 11450
rect 23704 11398 23734 11450
rect 23758 11398 23768 11450
rect 23768 11398 23814 11450
rect 23518 11396 23574 11398
rect 23598 11396 23654 11398
rect 23678 11396 23734 11398
rect 23758 11396 23814 11398
rect 31223 19066 31279 19068
rect 31303 19066 31359 19068
rect 31383 19066 31439 19068
rect 31463 19066 31519 19068
rect 31223 19014 31269 19066
rect 31269 19014 31279 19066
rect 31303 19014 31333 19066
rect 31333 19014 31345 19066
rect 31345 19014 31359 19066
rect 31383 19014 31397 19066
rect 31397 19014 31409 19066
rect 31409 19014 31439 19066
rect 31463 19014 31473 19066
rect 31473 19014 31519 19066
rect 31223 19012 31279 19014
rect 31303 19012 31359 19014
rect 31383 19012 31439 19014
rect 31463 19012 31519 19014
rect 27371 18522 27427 18524
rect 27451 18522 27507 18524
rect 27531 18522 27587 18524
rect 27611 18522 27667 18524
rect 27371 18470 27417 18522
rect 27417 18470 27427 18522
rect 27451 18470 27481 18522
rect 27481 18470 27493 18522
rect 27493 18470 27507 18522
rect 27531 18470 27545 18522
rect 27545 18470 27557 18522
rect 27557 18470 27587 18522
rect 27611 18470 27621 18522
rect 27621 18470 27667 18522
rect 27371 18468 27427 18470
rect 27451 18468 27507 18470
rect 27531 18468 27587 18470
rect 27611 18468 27667 18470
rect 31223 17978 31279 17980
rect 31303 17978 31359 17980
rect 31383 17978 31439 17980
rect 31463 17978 31519 17980
rect 31223 17926 31269 17978
rect 31269 17926 31279 17978
rect 31303 17926 31333 17978
rect 31333 17926 31345 17978
rect 31345 17926 31359 17978
rect 31383 17926 31397 17978
rect 31397 17926 31409 17978
rect 31409 17926 31439 17978
rect 31463 17926 31473 17978
rect 31473 17926 31519 17978
rect 31223 17924 31279 17926
rect 31303 17924 31359 17926
rect 31383 17924 31439 17926
rect 31463 17924 31519 17926
rect 27371 17434 27427 17436
rect 27451 17434 27507 17436
rect 27531 17434 27587 17436
rect 27611 17434 27667 17436
rect 27371 17382 27417 17434
rect 27417 17382 27427 17434
rect 27451 17382 27481 17434
rect 27481 17382 27493 17434
rect 27493 17382 27507 17434
rect 27531 17382 27545 17434
rect 27545 17382 27557 17434
rect 27557 17382 27587 17434
rect 27611 17382 27621 17434
rect 27621 17382 27667 17434
rect 27371 17380 27427 17382
rect 27451 17380 27507 17382
rect 27531 17380 27587 17382
rect 27611 17380 27667 17382
rect 31223 16890 31279 16892
rect 31303 16890 31359 16892
rect 31383 16890 31439 16892
rect 31463 16890 31519 16892
rect 31223 16838 31269 16890
rect 31269 16838 31279 16890
rect 31303 16838 31333 16890
rect 31333 16838 31345 16890
rect 31345 16838 31359 16890
rect 31383 16838 31397 16890
rect 31397 16838 31409 16890
rect 31409 16838 31439 16890
rect 31463 16838 31473 16890
rect 31473 16838 31519 16890
rect 31223 16836 31279 16838
rect 31303 16836 31359 16838
rect 31383 16836 31439 16838
rect 31463 16836 31519 16838
rect 27371 16346 27427 16348
rect 27451 16346 27507 16348
rect 27531 16346 27587 16348
rect 27611 16346 27667 16348
rect 27371 16294 27417 16346
rect 27417 16294 27427 16346
rect 27451 16294 27481 16346
rect 27481 16294 27493 16346
rect 27493 16294 27507 16346
rect 27531 16294 27545 16346
rect 27545 16294 27557 16346
rect 27557 16294 27587 16346
rect 27611 16294 27621 16346
rect 27621 16294 27667 16346
rect 27371 16292 27427 16294
rect 27451 16292 27507 16294
rect 27531 16292 27587 16294
rect 27611 16292 27667 16294
rect 25502 14476 25558 14512
rect 25502 14456 25504 14476
rect 25504 14456 25556 14476
rect 25556 14456 25558 14476
rect 24858 13096 24914 13152
rect 25686 13912 25742 13968
rect 26146 14184 26202 14240
rect 25962 14048 26018 14104
rect 25502 13504 25558 13560
rect 25318 13368 25374 13424
rect 31223 15802 31279 15804
rect 31303 15802 31359 15804
rect 31383 15802 31439 15804
rect 31463 15802 31519 15804
rect 31223 15750 31269 15802
rect 31269 15750 31279 15802
rect 31303 15750 31333 15802
rect 31333 15750 31345 15802
rect 31345 15750 31359 15802
rect 31383 15750 31397 15802
rect 31397 15750 31409 15802
rect 31409 15750 31439 15802
rect 31463 15750 31473 15802
rect 31473 15750 31519 15802
rect 31223 15748 31279 15750
rect 31303 15748 31359 15750
rect 31383 15748 31439 15750
rect 31463 15748 31519 15750
rect 31666 15680 31722 15736
rect 27371 15258 27427 15260
rect 27451 15258 27507 15260
rect 27531 15258 27587 15260
rect 27611 15258 27667 15260
rect 27371 15206 27417 15258
rect 27417 15206 27427 15258
rect 27451 15206 27481 15258
rect 27481 15206 27493 15258
rect 27493 15206 27507 15258
rect 27531 15206 27545 15258
rect 27545 15206 27557 15258
rect 27557 15206 27587 15258
rect 27611 15206 27621 15258
rect 27621 15206 27667 15258
rect 27371 15204 27427 15206
rect 27451 15204 27507 15206
rect 27531 15204 27587 15206
rect 27611 15204 27667 15206
rect 28262 15000 28318 15056
rect 28262 14320 28318 14376
rect 27371 14170 27427 14172
rect 27451 14170 27507 14172
rect 27531 14170 27587 14172
rect 27611 14170 27667 14172
rect 27371 14118 27417 14170
rect 27417 14118 27427 14170
rect 27451 14118 27481 14170
rect 27481 14118 27493 14170
rect 27493 14118 27507 14170
rect 27531 14118 27545 14170
rect 27545 14118 27557 14170
rect 27557 14118 27587 14170
rect 27611 14118 27621 14170
rect 27621 14118 27667 14170
rect 27371 14116 27427 14118
rect 27451 14116 27507 14118
rect 27531 14116 27587 14118
rect 27611 14116 27667 14118
rect 25594 12844 25650 12880
rect 25594 12824 25596 12844
rect 25596 12824 25648 12844
rect 25648 12824 25650 12844
rect 25226 12008 25282 12064
rect 24490 11636 24492 11656
rect 24492 11636 24544 11656
rect 24544 11636 24546 11656
rect 24490 11600 24546 11636
rect 26698 13232 26754 13288
rect 26146 12688 26202 12744
rect 27371 13082 27427 13084
rect 27451 13082 27507 13084
rect 27531 13082 27587 13084
rect 27611 13082 27667 13084
rect 27371 13030 27417 13082
rect 27417 13030 27427 13082
rect 27451 13030 27481 13082
rect 27481 13030 27493 13082
rect 27493 13030 27507 13082
rect 27531 13030 27545 13082
rect 27545 13030 27557 13082
rect 27557 13030 27587 13082
rect 27611 13030 27621 13082
rect 27621 13030 27667 13082
rect 27371 13028 27427 13030
rect 27451 13028 27507 13030
rect 27531 13028 27587 13030
rect 27611 13028 27667 13030
rect 28262 12960 28318 13016
rect 28262 12280 28318 12336
rect 27371 11994 27427 11996
rect 27451 11994 27507 11996
rect 27531 11994 27587 11996
rect 27611 11994 27667 11996
rect 27371 11942 27417 11994
rect 27417 11942 27427 11994
rect 27451 11942 27481 11994
rect 27481 11942 27493 11994
rect 27493 11942 27507 11994
rect 27531 11942 27545 11994
rect 27545 11942 27557 11994
rect 27557 11942 27587 11994
rect 27611 11942 27621 11994
rect 27621 11942 27667 11994
rect 27371 11940 27427 11942
rect 27451 11940 27507 11942
rect 27531 11940 27587 11942
rect 27611 11940 27667 11942
rect 31223 14714 31279 14716
rect 31303 14714 31359 14716
rect 31383 14714 31439 14716
rect 31463 14714 31519 14716
rect 31223 14662 31269 14714
rect 31269 14662 31279 14714
rect 31303 14662 31333 14714
rect 31333 14662 31345 14714
rect 31345 14662 31359 14714
rect 31383 14662 31397 14714
rect 31397 14662 31409 14714
rect 31409 14662 31439 14714
rect 31463 14662 31473 14714
rect 31473 14662 31519 14714
rect 31223 14660 31279 14662
rect 31303 14660 31359 14662
rect 31383 14660 31439 14662
rect 31463 14660 31519 14662
rect 31666 13640 31722 13696
rect 31223 13626 31279 13628
rect 31303 13626 31359 13628
rect 31383 13626 31439 13628
rect 31463 13626 31519 13628
rect 31223 13574 31269 13626
rect 31269 13574 31279 13626
rect 31303 13574 31333 13626
rect 31333 13574 31345 13626
rect 31345 13574 31359 13626
rect 31383 13574 31397 13626
rect 31397 13574 31409 13626
rect 31409 13574 31439 13626
rect 31463 13574 31473 13626
rect 31473 13574 31519 13626
rect 31223 13572 31279 13574
rect 31303 13572 31359 13574
rect 31383 13572 31439 13574
rect 31463 13572 31519 13574
rect 31223 12538 31279 12540
rect 31303 12538 31359 12540
rect 31383 12538 31439 12540
rect 31463 12538 31519 12540
rect 31223 12486 31269 12538
rect 31269 12486 31279 12538
rect 31303 12486 31333 12538
rect 31333 12486 31345 12538
rect 31345 12486 31359 12538
rect 31383 12486 31397 12538
rect 31397 12486 31409 12538
rect 31409 12486 31439 12538
rect 31463 12486 31473 12538
rect 31473 12486 31519 12538
rect 31223 12484 31279 12486
rect 31303 12484 31359 12486
rect 31383 12484 31439 12486
rect 31463 12484 31519 12486
rect 29642 11736 29698 11792
rect 25962 11636 25964 11656
rect 25964 11636 26016 11656
rect 26016 11636 26018 11656
rect 25962 11600 26018 11636
rect 28262 11600 28318 11656
rect 23518 10362 23574 10364
rect 23598 10362 23654 10364
rect 23678 10362 23734 10364
rect 23758 10362 23814 10364
rect 23518 10310 23564 10362
rect 23564 10310 23574 10362
rect 23598 10310 23628 10362
rect 23628 10310 23640 10362
rect 23640 10310 23654 10362
rect 23678 10310 23692 10362
rect 23692 10310 23704 10362
rect 23704 10310 23734 10362
rect 23758 10310 23768 10362
rect 23768 10310 23814 10362
rect 23518 10308 23574 10310
rect 23598 10308 23654 10310
rect 23678 10308 23734 10310
rect 23758 10308 23814 10310
rect 22374 9052 22376 9072
rect 22376 9052 22428 9072
rect 22428 9052 22430 9072
rect 22374 9016 22430 9052
rect 22006 8744 22062 8800
rect 22834 8508 22836 8528
rect 22836 8508 22888 8528
rect 22888 8508 22890 8528
rect 22834 8472 22890 8508
rect 21914 8356 21970 8392
rect 21914 8336 21916 8356
rect 21916 8336 21968 8356
rect 21968 8336 21970 8356
rect 20350 5752 20352 5772
rect 20352 5752 20404 5772
rect 20404 5752 20406 5772
rect 20534 5208 20590 5264
rect 20994 5480 21050 5536
rect 19666 4378 19722 4380
rect 19746 4378 19802 4380
rect 19826 4378 19882 4380
rect 19906 4378 19962 4380
rect 19666 4326 19712 4378
rect 19712 4326 19722 4378
rect 19746 4326 19776 4378
rect 19776 4326 19788 4378
rect 19788 4326 19802 4378
rect 19826 4326 19840 4378
rect 19840 4326 19852 4378
rect 19852 4326 19882 4378
rect 19906 4326 19916 4378
rect 19916 4326 19962 4378
rect 19666 4324 19722 4326
rect 19746 4324 19802 4326
rect 19826 4324 19882 4326
rect 19906 4324 19962 4326
rect 19666 3290 19722 3292
rect 19746 3290 19802 3292
rect 19826 3290 19882 3292
rect 19906 3290 19962 3292
rect 19666 3238 19712 3290
rect 19712 3238 19722 3290
rect 19746 3238 19776 3290
rect 19776 3238 19788 3290
rect 19788 3238 19802 3290
rect 19826 3238 19840 3290
rect 19840 3238 19852 3290
rect 19852 3238 19882 3290
rect 19906 3238 19916 3290
rect 19916 3238 19962 3290
rect 19666 3236 19722 3238
rect 19746 3236 19802 3238
rect 19826 3236 19882 3238
rect 19906 3236 19962 3238
rect 19666 2202 19722 2204
rect 19746 2202 19802 2204
rect 19826 2202 19882 2204
rect 19906 2202 19962 2204
rect 19666 2150 19712 2202
rect 19712 2150 19722 2202
rect 19746 2150 19776 2202
rect 19776 2150 19788 2202
rect 19788 2150 19802 2202
rect 19826 2150 19840 2202
rect 19840 2150 19852 2202
rect 19852 2150 19882 2202
rect 19906 2150 19916 2202
rect 19916 2150 19962 2202
rect 19666 2148 19722 2150
rect 19746 2148 19802 2150
rect 19826 2148 19882 2150
rect 19906 2148 19962 2150
rect 19666 1114 19722 1116
rect 19746 1114 19802 1116
rect 19826 1114 19882 1116
rect 19906 1114 19962 1116
rect 19666 1062 19712 1114
rect 19712 1062 19722 1114
rect 19746 1062 19776 1114
rect 19776 1062 19788 1114
rect 19788 1062 19802 1114
rect 19826 1062 19840 1114
rect 19840 1062 19852 1114
rect 19852 1062 19882 1114
rect 19906 1062 19916 1114
rect 19916 1062 19962 1114
rect 19666 1060 19722 1062
rect 19746 1060 19802 1062
rect 19826 1060 19882 1062
rect 19906 1060 19962 1062
rect 23294 8880 23350 8936
rect 23518 9274 23574 9276
rect 23598 9274 23654 9276
rect 23678 9274 23734 9276
rect 23758 9274 23814 9276
rect 23518 9222 23564 9274
rect 23564 9222 23574 9274
rect 23598 9222 23628 9274
rect 23628 9222 23640 9274
rect 23640 9222 23654 9274
rect 23678 9222 23692 9274
rect 23692 9222 23704 9274
rect 23704 9222 23734 9274
rect 23758 9222 23768 9274
rect 23768 9222 23814 9274
rect 23518 9220 23574 9222
rect 23598 9220 23654 9222
rect 23678 9220 23734 9222
rect 23758 9220 23814 9222
rect 31223 11450 31279 11452
rect 31303 11450 31359 11452
rect 31383 11450 31439 11452
rect 31463 11450 31519 11452
rect 31223 11398 31269 11450
rect 31269 11398 31279 11450
rect 31303 11398 31333 11450
rect 31333 11398 31345 11450
rect 31345 11398 31359 11450
rect 31383 11398 31397 11450
rect 31397 11398 31409 11450
rect 31409 11398 31439 11450
rect 31463 11398 31473 11450
rect 31473 11398 31519 11450
rect 31223 11396 31279 11398
rect 31303 11396 31359 11398
rect 31383 11396 31439 11398
rect 31463 11396 31519 11398
rect 28262 10920 28318 10976
rect 27371 10906 27427 10908
rect 27451 10906 27507 10908
rect 27531 10906 27587 10908
rect 27611 10906 27667 10908
rect 27371 10854 27417 10906
rect 27417 10854 27427 10906
rect 27451 10854 27481 10906
rect 27481 10854 27493 10906
rect 27493 10854 27507 10906
rect 27531 10854 27545 10906
rect 27545 10854 27557 10906
rect 27557 10854 27587 10906
rect 27611 10854 27621 10906
rect 27621 10854 27667 10906
rect 27371 10852 27427 10854
rect 27451 10852 27507 10854
rect 27531 10852 27587 10854
rect 27611 10852 27667 10854
rect 24030 9560 24086 9616
rect 23518 8186 23574 8188
rect 23598 8186 23654 8188
rect 23678 8186 23734 8188
rect 23758 8186 23814 8188
rect 23518 8134 23564 8186
rect 23564 8134 23574 8186
rect 23598 8134 23628 8186
rect 23628 8134 23640 8186
rect 23640 8134 23654 8186
rect 23678 8134 23692 8186
rect 23692 8134 23704 8186
rect 23704 8134 23734 8186
rect 23758 8134 23768 8186
rect 23768 8134 23814 8186
rect 23518 8132 23574 8134
rect 23598 8132 23654 8134
rect 23678 8132 23734 8134
rect 23758 8132 23814 8134
rect 22006 6568 22062 6624
rect 21638 6296 21694 6352
rect 21546 5752 21602 5808
rect 21730 6196 21732 6216
rect 21732 6196 21784 6216
rect 21784 6196 21786 6216
rect 21730 6160 21786 6196
rect 23754 7656 23810 7712
rect 23202 7148 23204 7168
rect 23204 7148 23256 7168
rect 23256 7148 23258 7168
rect 23202 7112 23258 7148
rect 23518 7098 23574 7100
rect 23598 7098 23654 7100
rect 23678 7098 23734 7100
rect 23758 7098 23814 7100
rect 23518 7046 23564 7098
rect 23564 7046 23574 7098
rect 23598 7046 23628 7098
rect 23628 7046 23640 7098
rect 23640 7046 23654 7098
rect 23678 7046 23692 7098
rect 23692 7046 23704 7098
rect 23704 7046 23734 7098
rect 23758 7046 23768 7098
rect 23768 7046 23814 7098
rect 23518 7044 23574 7046
rect 23598 7044 23654 7046
rect 23678 7044 23734 7046
rect 23758 7044 23814 7046
rect 22282 6196 22284 6216
rect 22284 6196 22336 6216
rect 22336 6196 22338 6216
rect 22282 6160 22338 6196
rect 21914 6024 21970 6080
rect 22006 5752 22062 5808
rect 21454 5364 21510 5400
rect 21454 5344 21456 5364
rect 21456 5344 21508 5364
rect 21508 5344 21510 5364
rect 22190 5616 22246 5672
rect 22466 5888 22522 5944
rect 22650 6840 22706 6896
rect 23110 6704 23166 6760
rect 22650 6160 22706 6216
rect 22282 5208 22338 5264
rect 23478 6296 23534 6352
rect 23110 6024 23166 6080
rect 23018 5752 23074 5808
rect 23938 8744 23994 8800
rect 24214 7520 24270 7576
rect 24122 6840 24178 6896
rect 23518 6010 23574 6012
rect 23598 6010 23654 6012
rect 23678 6010 23734 6012
rect 23758 6010 23814 6012
rect 23518 5958 23564 6010
rect 23564 5958 23574 6010
rect 23598 5958 23628 6010
rect 23628 5958 23640 6010
rect 23640 5958 23654 6010
rect 23678 5958 23692 6010
rect 23692 5958 23704 6010
rect 23704 5958 23734 6010
rect 23758 5958 23768 6010
rect 23768 5958 23814 6010
rect 23518 5956 23574 5958
rect 23598 5956 23654 5958
rect 23678 5956 23734 5958
rect 23758 5956 23814 5958
rect 23518 4922 23574 4924
rect 23598 4922 23654 4924
rect 23678 4922 23734 4924
rect 23758 4922 23814 4924
rect 23518 4870 23564 4922
rect 23564 4870 23574 4922
rect 23598 4870 23628 4922
rect 23628 4870 23640 4922
rect 23640 4870 23654 4922
rect 23678 4870 23692 4922
rect 23692 4870 23704 4922
rect 23704 4870 23734 4922
rect 23758 4870 23768 4922
rect 23768 4870 23814 4922
rect 23518 4868 23574 4870
rect 23598 4868 23654 4870
rect 23678 4868 23734 4870
rect 23758 4868 23814 4870
rect 24674 8200 24730 8256
rect 24490 7112 24546 7168
rect 24030 5480 24086 5536
rect 24766 6568 24822 6624
rect 31223 10362 31279 10364
rect 31303 10362 31359 10364
rect 31383 10362 31439 10364
rect 31463 10362 31519 10364
rect 31223 10310 31269 10362
rect 31269 10310 31279 10362
rect 31303 10310 31333 10362
rect 31333 10310 31345 10362
rect 31345 10310 31359 10362
rect 31383 10310 31397 10362
rect 31397 10310 31409 10362
rect 31409 10310 31439 10362
rect 31463 10310 31473 10362
rect 31473 10310 31519 10362
rect 31223 10308 31279 10310
rect 31303 10308 31359 10310
rect 31383 10308 31439 10310
rect 31463 10308 31519 10310
rect 31666 10240 31722 10296
rect 27371 9818 27427 9820
rect 27451 9818 27507 9820
rect 27531 9818 27587 9820
rect 27611 9818 27667 9820
rect 27371 9766 27417 9818
rect 27417 9766 27427 9818
rect 27451 9766 27481 9818
rect 27481 9766 27493 9818
rect 27493 9766 27507 9818
rect 27531 9766 27545 9818
rect 27545 9766 27557 9818
rect 27557 9766 27587 9818
rect 27611 9766 27621 9818
rect 27621 9766 27667 9818
rect 27371 9764 27427 9766
rect 27451 9764 27507 9766
rect 27531 9764 27587 9766
rect 27611 9764 27667 9766
rect 28262 9560 28318 9616
rect 25594 8472 25650 8528
rect 25042 6704 25098 6760
rect 25594 7656 25650 7712
rect 25594 6840 25650 6896
rect 25134 5344 25190 5400
rect 31223 9274 31279 9276
rect 31303 9274 31359 9276
rect 31383 9274 31439 9276
rect 31463 9274 31519 9276
rect 31223 9222 31269 9274
rect 31269 9222 31279 9274
rect 31303 9222 31333 9274
rect 31333 9222 31345 9274
rect 31345 9222 31359 9274
rect 31383 9222 31397 9274
rect 31397 9222 31409 9274
rect 31409 9222 31439 9274
rect 31463 9222 31473 9274
rect 31473 9222 31519 9274
rect 31223 9220 31279 9222
rect 31303 9220 31359 9222
rect 31383 9220 31439 9222
rect 31463 9220 31519 9222
rect 27371 8730 27427 8732
rect 27451 8730 27507 8732
rect 27531 8730 27587 8732
rect 27611 8730 27667 8732
rect 27371 8678 27417 8730
rect 27417 8678 27427 8730
rect 27451 8678 27481 8730
rect 27481 8678 27493 8730
rect 27493 8678 27507 8730
rect 27531 8678 27545 8730
rect 27545 8678 27557 8730
rect 27557 8678 27587 8730
rect 27611 8678 27621 8730
rect 27621 8678 27667 8730
rect 27371 8676 27427 8678
rect 27451 8676 27507 8678
rect 27531 8676 27587 8678
rect 27611 8676 27667 8678
rect 31666 8472 31722 8528
rect 25962 7112 26018 7168
rect 31666 8200 31722 8256
rect 31223 8186 31279 8188
rect 31303 8186 31359 8188
rect 31383 8186 31439 8188
rect 31463 8186 31519 8188
rect 31223 8134 31269 8186
rect 31269 8134 31279 8186
rect 31303 8134 31333 8186
rect 31333 8134 31345 8186
rect 31345 8134 31359 8186
rect 31383 8134 31397 8186
rect 31397 8134 31409 8186
rect 31409 8134 31439 8186
rect 31463 8134 31473 8186
rect 31473 8134 31519 8186
rect 31223 8132 31279 8134
rect 31303 8132 31359 8134
rect 31383 8132 31439 8134
rect 31463 8132 31519 8134
rect 27371 7642 27427 7644
rect 27451 7642 27507 7644
rect 27531 7642 27587 7644
rect 27611 7642 27667 7644
rect 27371 7590 27417 7642
rect 27417 7590 27427 7642
rect 27451 7590 27481 7642
rect 27481 7590 27493 7642
rect 27493 7590 27507 7642
rect 27531 7590 27545 7642
rect 27545 7590 27557 7642
rect 27557 7590 27587 7642
rect 27611 7590 27621 7642
rect 27621 7590 27667 7642
rect 27371 7588 27427 7590
rect 27451 7588 27507 7590
rect 27531 7588 27587 7590
rect 27611 7588 27667 7590
rect 26330 7520 26386 7576
rect 31666 7248 31722 7304
rect 31223 7098 31279 7100
rect 31303 7098 31359 7100
rect 31383 7098 31439 7100
rect 31463 7098 31519 7100
rect 31223 7046 31269 7098
rect 31269 7046 31279 7098
rect 31303 7046 31333 7098
rect 31333 7046 31345 7098
rect 31345 7046 31359 7098
rect 31383 7046 31397 7098
rect 31397 7046 31409 7098
rect 31409 7046 31439 7098
rect 31463 7046 31473 7098
rect 31473 7046 31519 7098
rect 31223 7044 31279 7046
rect 31303 7044 31359 7046
rect 31383 7044 31439 7046
rect 31463 7044 31519 7046
rect 27371 6554 27427 6556
rect 27451 6554 27507 6556
rect 27531 6554 27587 6556
rect 27611 6554 27667 6556
rect 27371 6502 27417 6554
rect 27417 6502 27427 6554
rect 27451 6502 27481 6554
rect 27481 6502 27493 6554
rect 27493 6502 27507 6554
rect 27531 6502 27545 6554
rect 27545 6502 27557 6554
rect 27557 6502 27587 6554
rect 27611 6502 27621 6554
rect 27621 6502 27667 6554
rect 27371 6500 27427 6502
rect 27451 6500 27507 6502
rect 27531 6500 27587 6502
rect 27611 6500 27667 6502
rect 31223 6010 31279 6012
rect 31303 6010 31359 6012
rect 31383 6010 31439 6012
rect 31463 6010 31519 6012
rect 31223 5958 31269 6010
rect 31269 5958 31279 6010
rect 31303 5958 31333 6010
rect 31333 5958 31345 6010
rect 31345 5958 31359 6010
rect 31383 5958 31397 6010
rect 31397 5958 31409 6010
rect 31409 5958 31439 6010
rect 31463 5958 31473 6010
rect 31473 5958 31519 6010
rect 31223 5956 31279 5958
rect 31303 5956 31359 5958
rect 31383 5956 31439 5958
rect 31463 5956 31519 5958
rect 27371 5466 27427 5468
rect 27451 5466 27507 5468
rect 27531 5466 27587 5468
rect 27611 5466 27667 5468
rect 27371 5414 27417 5466
rect 27417 5414 27427 5466
rect 27451 5414 27481 5466
rect 27481 5414 27493 5466
rect 27493 5414 27507 5466
rect 27531 5414 27545 5466
rect 27545 5414 27557 5466
rect 27557 5414 27587 5466
rect 27611 5414 27621 5466
rect 27621 5414 27667 5466
rect 27371 5412 27427 5414
rect 27451 5412 27507 5414
rect 27531 5412 27587 5414
rect 27611 5412 27667 5414
rect 31223 4922 31279 4924
rect 31303 4922 31359 4924
rect 31383 4922 31439 4924
rect 31463 4922 31519 4924
rect 31223 4870 31269 4922
rect 31269 4870 31279 4922
rect 31303 4870 31333 4922
rect 31333 4870 31345 4922
rect 31345 4870 31359 4922
rect 31383 4870 31397 4922
rect 31397 4870 31409 4922
rect 31409 4870 31439 4922
rect 31463 4870 31473 4922
rect 31473 4870 31519 4922
rect 31223 4868 31279 4870
rect 31303 4868 31359 4870
rect 31383 4868 31439 4870
rect 31463 4868 31519 4870
rect 31666 4800 31722 4856
rect 27371 4378 27427 4380
rect 27451 4378 27507 4380
rect 27531 4378 27587 4380
rect 27611 4378 27667 4380
rect 27371 4326 27417 4378
rect 27417 4326 27427 4378
rect 27451 4326 27481 4378
rect 27481 4326 27493 4378
rect 27493 4326 27507 4378
rect 27531 4326 27545 4378
rect 27545 4326 27557 4378
rect 27557 4326 27587 4378
rect 27611 4326 27621 4378
rect 27621 4326 27667 4378
rect 27371 4324 27427 4326
rect 27451 4324 27507 4326
rect 27531 4324 27587 4326
rect 27611 4324 27667 4326
rect 23518 3834 23574 3836
rect 23598 3834 23654 3836
rect 23678 3834 23734 3836
rect 23758 3834 23814 3836
rect 23518 3782 23564 3834
rect 23564 3782 23574 3834
rect 23598 3782 23628 3834
rect 23628 3782 23640 3834
rect 23640 3782 23654 3834
rect 23678 3782 23692 3834
rect 23692 3782 23704 3834
rect 23704 3782 23734 3834
rect 23758 3782 23768 3834
rect 23768 3782 23814 3834
rect 23518 3780 23574 3782
rect 23598 3780 23654 3782
rect 23678 3780 23734 3782
rect 23758 3780 23814 3782
rect 31223 3834 31279 3836
rect 31303 3834 31359 3836
rect 31383 3834 31439 3836
rect 31463 3834 31519 3836
rect 31223 3782 31269 3834
rect 31269 3782 31279 3834
rect 31303 3782 31333 3834
rect 31333 3782 31345 3834
rect 31345 3782 31359 3834
rect 31383 3782 31397 3834
rect 31397 3782 31409 3834
rect 31409 3782 31439 3834
rect 31463 3782 31473 3834
rect 31473 3782 31519 3834
rect 31223 3780 31279 3782
rect 31303 3780 31359 3782
rect 31383 3780 31439 3782
rect 31463 3780 31519 3782
rect 27371 3290 27427 3292
rect 27451 3290 27507 3292
rect 27531 3290 27587 3292
rect 27611 3290 27667 3292
rect 27371 3238 27417 3290
rect 27417 3238 27427 3290
rect 27451 3238 27481 3290
rect 27481 3238 27493 3290
rect 27493 3238 27507 3290
rect 27531 3238 27545 3290
rect 27545 3238 27557 3290
rect 27557 3238 27587 3290
rect 27611 3238 27621 3290
rect 27621 3238 27667 3290
rect 27371 3236 27427 3238
rect 27451 3236 27507 3238
rect 27531 3236 27587 3238
rect 27611 3236 27667 3238
rect 23518 2746 23574 2748
rect 23598 2746 23654 2748
rect 23678 2746 23734 2748
rect 23758 2746 23814 2748
rect 23518 2694 23564 2746
rect 23564 2694 23574 2746
rect 23598 2694 23628 2746
rect 23628 2694 23640 2746
rect 23640 2694 23654 2746
rect 23678 2694 23692 2746
rect 23692 2694 23704 2746
rect 23704 2694 23734 2746
rect 23758 2694 23768 2746
rect 23768 2694 23814 2746
rect 23518 2692 23574 2694
rect 23598 2692 23654 2694
rect 23678 2692 23734 2694
rect 23758 2692 23814 2694
rect 31223 2746 31279 2748
rect 31303 2746 31359 2748
rect 31383 2746 31439 2748
rect 31463 2746 31519 2748
rect 31223 2694 31269 2746
rect 31269 2694 31279 2746
rect 31303 2694 31333 2746
rect 31333 2694 31345 2746
rect 31345 2694 31359 2746
rect 31383 2694 31397 2746
rect 31397 2694 31409 2746
rect 31409 2694 31439 2746
rect 31463 2694 31473 2746
rect 31473 2694 31519 2746
rect 31223 2692 31279 2694
rect 31303 2692 31359 2694
rect 31383 2692 31439 2694
rect 31463 2692 31519 2694
rect 27371 2202 27427 2204
rect 27451 2202 27507 2204
rect 27531 2202 27587 2204
rect 27611 2202 27667 2204
rect 27371 2150 27417 2202
rect 27417 2150 27427 2202
rect 27451 2150 27481 2202
rect 27481 2150 27493 2202
rect 27493 2150 27507 2202
rect 27531 2150 27545 2202
rect 27545 2150 27557 2202
rect 27557 2150 27587 2202
rect 27611 2150 27621 2202
rect 27621 2150 27667 2202
rect 27371 2148 27427 2150
rect 27451 2148 27507 2150
rect 27531 2148 27587 2150
rect 27611 2148 27667 2150
rect 23518 1658 23574 1660
rect 23598 1658 23654 1660
rect 23678 1658 23734 1660
rect 23758 1658 23814 1660
rect 23518 1606 23564 1658
rect 23564 1606 23574 1658
rect 23598 1606 23628 1658
rect 23628 1606 23640 1658
rect 23640 1606 23654 1658
rect 23678 1606 23692 1658
rect 23692 1606 23704 1658
rect 23704 1606 23734 1658
rect 23758 1606 23768 1658
rect 23768 1606 23814 1658
rect 23518 1604 23574 1606
rect 23598 1604 23654 1606
rect 23678 1604 23734 1606
rect 23758 1604 23814 1606
rect 31223 1658 31279 1660
rect 31303 1658 31359 1660
rect 31383 1658 31439 1660
rect 31463 1658 31519 1660
rect 31223 1606 31269 1658
rect 31269 1606 31279 1658
rect 31303 1606 31333 1658
rect 31333 1606 31345 1658
rect 31345 1606 31359 1658
rect 31383 1606 31397 1658
rect 31397 1606 31409 1658
rect 31409 1606 31439 1658
rect 31463 1606 31473 1658
rect 31473 1606 31519 1658
rect 31223 1604 31279 1606
rect 31303 1604 31359 1606
rect 31383 1604 31439 1606
rect 31463 1604 31519 1606
rect 27371 1114 27427 1116
rect 27451 1114 27507 1116
rect 27531 1114 27587 1116
rect 27611 1114 27667 1116
rect 27371 1062 27417 1114
rect 27417 1062 27427 1114
rect 27451 1062 27481 1114
rect 27481 1062 27493 1114
rect 27493 1062 27507 1114
rect 27531 1062 27545 1114
rect 27545 1062 27557 1114
rect 27557 1062 27587 1114
rect 27611 1062 27621 1114
rect 27621 1062 27667 1114
rect 27371 1060 27427 1062
rect 27451 1060 27507 1062
rect 27531 1060 27587 1062
rect 27611 1060 27667 1062
rect 23518 570 23574 572
rect 23598 570 23654 572
rect 23678 570 23734 572
rect 23758 570 23814 572
rect 23518 518 23564 570
rect 23564 518 23574 570
rect 23598 518 23628 570
rect 23628 518 23640 570
rect 23640 518 23654 570
rect 23678 518 23692 570
rect 23692 518 23704 570
rect 23704 518 23734 570
rect 23758 518 23768 570
rect 23768 518 23814 570
rect 23518 516 23574 518
rect 23598 516 23654 518
rect 23678 516 23734 518
rect 23758 516 23814 518
rect 31223 570 31279 572
rect 31303 570 31359 572
rect 31383 570 31439 572
rect 31463 570 31519 572
rect 31223 518 31269 570
rect 31269 518 31279 570
rect 31303 518 31333 570
rect 31333 518 31345 570
rect 31345 518 31359 570
rect 31383 518 31397 570
rect 31397 518 31409 570
rect 31409 518 31439 570
rect 31463 518 31473 570
rect 31473 518 31519 570
rect 31223 516 31279 518
rect 31303 516 31359 518
rect 31383 516 31439 518
rect 31463 516 31519 518
<< metal3 >>
rect 8098 19072 8414 19073
rect 8098 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8414 19072
rect 8098 19007 8414 19008
rect 15803 19072 16119 19073
rect 15803 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16119 19072
rect 15803 19007 16119 19008
rect 23508 19072 23824 19073
rect 23508 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23824 19072
rect 23508 19007 23824 19008
rect 31213 19072 31529 19073
rect 31213 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31529 19072
rect 31213 19007 31529 19008
rect 11646 18668 11652 18732
rect 11716 18730 11722 18732
rect 12249 18730 12315 18733
rect 11716 18728 12315 18730
rect 11716 18672 12254 18728
rect 12310 18672 12315 18728
rect 11716 18670 12315 18672
rect 11716 18668 11722 18670
rect 12249 18667 12315 18670
rect 4246 18528 4562 18529
rect 4246 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4562 18528
rect 4246 18463 4562 18464
rect 11951 18528 12267 18529
rect 11951 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12267 18528
rect 11951 18463 12267 18464
rect 19656 18528 19972 18529
rect 19656 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19972 18528
rect 19656 18463 19972 18464
rect 27361 18528 27677 18529
rect 27361 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27677 18528
rect 27361 18463 27677 18464
rect 8098 17984 8414 17985
rect 8098 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8414 17984
rect 8098 17919 8414 17920
rect 15803 17984 16119 17985
rect 15803 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16119 17984
rect 15803 17919 16119 17920
rect 23508 17984 23824 17985
rect 23508 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23824 17984
rect 23508 17919 23824 17920
rect 31213 17984 31529 17985
rect 31213 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31529 17984
rect 31213 17919 31529 17920
rect 4246 17440 4562 17441
rect 4246 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4562 17440
rect 4246 17375 4562 17376
rect 11951 17440 12267 17441
rect 11951 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12267 17440
rect 11951 17375 12267 17376
rect 19656 17440 19972 17441
rect 19656 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19972 17440
rect 19656 17375 19972 17376
rect 27361 17440 27677 17441
rect 27361 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27677 17440
rect 27361 17375 27677 17376
rect 19333 17100 19399 17101
rect 19333 17096 19380 17100
rect 19444 17098 19450 17100
rect 21541 17098 21607 17101
rect 24209 17098 24275 17101
rect 19333 17040 19338 17096
rect 19333 17036 19380 17040
rect 19444 17038 19490 17098
rect 21541 17096 24275 17098
rect 21541 17040 21546 17096
rect 21602 17040 24214 17096
rect 24270 17040 24275 17096
rect 21541 17038 24275 17040
rect 19444 17036 19450 17038
rect 19333 17035 19399 17036
rect 21541 17035 21607 17038
rect 24209 17035 24275 17038
rect 10961 16962 11027 16965
rect 11278 16962 11284 16964
rect 10961 16960 11284 16962
rect 10961 16904 10966 16960
rect 11022 16904 11284 16960
rect 10961 16902 11284 16904
rect 10961 16899 11027 16902
rect 11278 16900 11284 16902
rect 11348 16900 11354 16964
rect 20345 16962 20411 16965
rect 21725 16962 21791 16965
rect 20345 16960 21791 16962
rect 20345 16904 20350 16960
rect 20406 16904 21730 16960
rect 21786 16904 21791 16960
rect 20345 16902 21791 16904
rect 20345 16899 20411 16902
rect 21725 16899 21791 16902
rect 22001 16962 22067 16965
rect 22829 16962 22895 16965
rect 22001 16960 22895 16962
rect 22001 16904 22006 16960
rect 22062 16904 22834 16960
rect 22890 16904 22895 16960
rect 22001 16902 22895 16904
rect 22001 16899 22067 16902
rect 22829 16899 22895 16902
rect 8098 16896 8414 16897
rect 8098 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8414 16896
rect 8098 16831 8414 16832
rect 15803 16896 16119 16897
rect 15803 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16119 16896
rect 15803 16831 16119 16832
rect 23508 16896 23824 16897
rect 23508 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23824 16896
rect 23508 16831 23824 16832
rect 31213 16896 31529 16897
rect 31213 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31529 16896
rect 31213 16831 31529 16832
rect 10358 16764 10364 16828
rect 10428 16826 10434 16828
rect 20345 16826 20411 16829
rect 22921 16826 22987 16829
rect 10428 16766 11024 16826
rect 10428 16764 10434 16766
rect 10964 16693 11024 16766
rect 20345 16824 22987 16826
rect 20345 16768 20350 16824
rect 20406 16768 22926 16824
rect 22982 16768 22987 16824
rect 20345 16766 22987 16768
rect 20345 16763 20411 16766
rect 22921 16763 22987 16766
rect 10225 16690 10291 16693
rect 10961 16690 11027 16693
rect 12617 16690 12683 16693
rect 10225 16688 10794 16690
rect 10225 16632 10230 16688
rect 10286 16632 10794 16688
rect 10225 16630 10794 16632
rect 10225 16627 10291 16630
rect 10041 16556 10107 16557
rect 9990 16554 9996 16556
rect 9950 16494 9996 16554
rect 10060 16552 10107 16556
rect 10102 16496 10107 16552
rect 9990 16492 9996 16494
rect 10060 16492 10107 16496
rect 10041 16491 10107 16492
rect 10317 16554 10383 16557
rect 10734 16556 10794 16630
rect 10961 16688 12683 16690
rect 10961 16632 10966 16688
rect 11022 16632 12622 16688
rect 12678 16632 12683 16688
rect 10961 16630 12683 16632
rect 10961 16627 11027 16630
rect 12617 16627 12683 16630
rect 10542 16554 10548 16556
rect 10317 16552 10548 16554
rect 10317 16496 10322 16552
rect 10378 16496 10548 16552
rect 10317 16494 10548 16496
rect 10317 16491 10383 16494
rect 10542 16492 10548 16494
rect 10612 16492 10618 16556
rect 10726 16492 10732 16556
rect 10796 16492 10802 16556
rect 21173 16554 21239 16557
rect 21449 16554 21515 16557
rect 21173 16552 21515 16554
rect 21173 16496 21178 16552
rect 21234 16496 21454 16552
rect 21510 16496 21515 16552
rect 21173 16494 21515 16496
rect 21173 16491 21239 16494
rect 21449 16491 21515 16494
rect 10041 16418 10107 16421
rect 11237 16418 11303 16421
rect 10041 16416 11303 16418
rect 10041 16360 10046 16416
rect 10102 16360 11242 16416
rect 11298 16360 11303 16416
rect 10041 16358 11303 16360
rect 10041 16355 10107 16358
rect 11237 16355 11303 16358
rect 22829 16418 22895 16421
rect 24853 16418 24919 16421
rect 22829 16416 24919 16418
rect 22829 16360 22834 16416
rect 22890 16360 24858 16416
rect 24914 16360 24919 16416
rect 22829 16358 24919 16360
rect 22829 16355 22895 16358
rect 24853 16355 24919 16358
rect 4246 16352 4562 16353
rect 4246 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4562 16352
rect 4246 16287 4562 16288
rect 11951 16352 12267 16353
rect 11951 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12267 16352
rect 11951 16287 12267 16288
rect 19656 16352 19972 16353
rect 19656 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19972 16352
rect 19656 16287 19972 16288
rect 27361 16352 27677 16353
rect 27361 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27677 16352
rect 27361 16287 27677 16288
rect 9581 16282 9647 16285
rect 11513 16282 11579 16285
rect 9581 16280 11579 16282
rect 9581 16224 9586 16280
rect 9642 16224 11518 16280
rect 11574 16224 11579 16280
rect 9581 16222 11579 16224
rect 9581 16219 9647 16222
rect 11513 16219 11579 16222
rect 20437 16282 20503 16285
rect 22277 16282 22343 16285
rect 20437 16280 22343 16282
rect 20437 16224 20442 16280
rect 20498 16224 22282 16280
rect 22338 16224 22343 16280
rect 20437 16222 22343 16224
rect 20437 16219 20503 16222
rect 22277 16219 22343 16222
rect 23289 16282 23355 16285
rect 25037 16282 25103 16285
rect 23289 16280 25103 16282
rect 23289 16224 23294 16280
rect 23350 16224 25042 16280
rect 25098 16224 25103 16280
rect 23289 16222 25103 16224
rect 23289 16219 23355 16222
rect 25037 16219 25103 16222
rect 8477 16146 8543 16149
rect 14089 16146 14155 16149
rect 8477 16144 14155 16146
rect 8477 16088 8482 16144
rect 8538 16088 14094 16144
rect 14150 16088 14155 16144
rect 8477 16086 14155 16088
rect 8477 16083 8543 16086
rect 14089 16083 14155 16086
rect 22369 16146 22435 16149
rect 24025 16146 24091 16149
rect 22369 16144 24091 16146
rect 22369 16088 22374 16144
rect 22430 16088 24030 16144
rect 24086 16088 24091 16144
rect 22369 16086 24091 16088
rect 22369 16083 22435 16086
rect 24025 16083 24091 16086
rect 7833 16010 7899 16013
rect 10961 16010 11027 16013
rect 7833 16008 11027 16010
rect 7833 15952 7838 16008
rect 7894 15952 10966 16008
rect 11022 15952 11027 16008
rect 7833 15950 11027 15952
rect 7833 15947 7899 15950
rect 10961 15947 11027 15950
rect 11329 16010 11395 16013
rect 12985 16010 13051 16013
rect 11329 16008 13051 16010
rect 11329 15952 11334 16008
rect 11390 15952 12990 16008
rect 13046 15952 13051 16008
rect 11329 15950 13051 15952
rect 11329 15947 11395 15950
rect 12985 15947 13051 15950
rect 13302 15948 13308 16012
rect 13372 16010 13378 16012
rect 13537 16010 13603 16013
rect 13372 16008 13603 16010
rect 13372 15952 13542 16008
rect 13598 15952 13603 16008
rect 13372 15950 13603 15952
rect 13372 15948 13378 15950
rect 13537 15947 13603 15950
rect 22318 15948 22324 16012
rect 22388 16010 22394 16012
rect 22553 16010 22619 16013
rect 23657 16010 23723 16013
rect 22388 16008 22619 16010
rect 22388 15952 22558 16008
rect 22614 15952 22619 16008
rect 22388 15950 22619 15952
rect 22388 15948 22394 15950
rect 22553 15947 22619 15950
rect 22694 16008 23723 16010
rect 22694 15952 23662 16008
rect 23718 15952 23723 16008
rect 22694 15950 23723 15952
rect 9121 15874 9187 15877
rect 13629 15874 13695 15877
rect 9121 15872 13695 15874
rect 9121 15816 9126 15872
rect 9182 15816 13634 15872
rect 13690 15816 13695 15872
rect 9121 15814 13695 15816
rect 9121 15811 9187 15814
rect 13629 15811 13695 15814
rect 21357 15874 21423 15877
rect 21633 15874 21699 15877
rect 22694 15874 22754 15950
rect 23657 15947 23723 15950
rect 23841 16010 23907 16013
rect 23974 16010 23980 16012
rect 23841 16008 23980 16010
rect 23841 15952 23846 16008
rect 23902 15952 23980 16008
rect 23841 15950 23980 15952
rect 23841 15947 23907 15950
rect 23974 15948 23980 15950
rect 24044 15948 24050 16012
rect 21357 15872 22754 15874
rect 21357 15816 21362 15872
rect 21418 15816 21638 15872
rect 21694 15816 22754 15872
rect 21357 15814 22754 15816
rect 21357 15811 21423 15814
rect 21633 15811 21699 15814
rect 8098 15808 8414 15809
rect 8098 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8414 15808
rect 8098 15743 8414 15744
rect 15803 15808 16119 15809
rect 15803 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16119 15808
rect 15803 15743 16119 15744
rect 23508 15808 23824 15809
rect 23508 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23824 15808
rect 23508 15743 23824 15744
rect 31213 15808 31529 15809
rect 31213 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31529 15808
rect 31213 15743 31529 15744
rect 9673 15738 9739 15741
rect 11145 15740 11211 15741
rect 9806 15738 9812 15740
rect 9673 15736 9812 15738
rect 9673 15680 9678 15736
rect 9734 15680 9812 15736
rect 9673 15678 9812 15680
rect 9673 15675 9739 15678
rect 9806 15676 9812 15678
rect 9876 15676 9882 15740
rect 11094 15738 11100 15740
rect 11054 15678 11100 15738
rect 11164 15736 11211 15740
rect 11206 15680 11211 15736
rect 11094 15676 11100 15678
rect 11164 15676 11211 15680
rect 11145 15675 11211 15676
rect 21817 15738 21883 15741
rect 21950 15738 21956 15740
rect 21817 15736 21956 15738
rect 21817 15680 21822 15736
rect 21878 15680 21956 15736
rect 21817 15678 21956 15680
rect 21817 15675 21883 15678
rect 21950 15676 21956 15678
rect 22020 15676 22026 15740
rect 31600 15736 32000 15768
rect 31600 15680 31666 15736
rect 31722 15680 32000 15736
rect 31600 15648 32000 15680
rect 9489 15602 9555 15605
rect 11053 15602 11119 15605
rect 9489 15600 11119 15602
rect 9489 15544 9494 15600
rect 9550 15544 11058 15600
rect 11114 15544 11119 15600
rect 9489 15542 11119 15544
rect 9489 15539 9555 15542
rect 11053 15539 11119 15542
rect 21909 15602 21975 15605
rect 24894 15602 24900 15604
rect 21909 15600 24900 15602
rect 21909 15544 21914 15600
rect 21970 15544 24900 15600
rect 21909 15542 24900 15544
rect 21909 15539 21975 15542
rect 24894 15540 24900 15542
rect 24964 15540 24970 15604
rect 9305 15466 9371 15469
rect 11973 15466 12039 15469
rect 9305 15464 12039 15466
rect 9305 15408 9310 15464
rect 9366 15408 11978 15464
rect 12034 15408 12039 15464
rect 9305 15406 12039 15408
rect 9305 15403 9371 15406
rect 11973 15403 12039 15406
rect 22185 15466 22251 15469
rect 23238 15466 23244 15468
rect 22185 15464 23244 15466
rect 22185 15408 22190 15464
rect 22246 15408 23244 15464
rect 22185 15406 23244 15408
rect 22185 15403 22251 15406
rect 23238 15404 23244 15406
rect 23308 15404 23314 15468
rect 23841 15466 23907 15469
rect 24301 15466 24367 15469
rect 23841 15464 24367 15466
rect 23841 15408 23846 15464
rect 23902 15408 24306 15464
rect 24362 15408 24367 15464
rect 23841 15406 24367 15408
rect 23841 15403 23907 15406
rect 24301 15403 24367 15406
rect 7373 15330 7439 15333
rect 10133 15330 10199 15333
rect 7373 15328 10199 15330
rect 7373 15272 7378 15328
rect 7434 15272 10138 15328
rect 10194 15272 10199 15328
rect 7373 15270 10199 15272
rect 7373 15267 7439 15270
rect 10133 15267 10199 15270
rect 10358 15268 10364 15332
rect 10428 15330 10434 15332
rect 10593 15330 10659 15333
rect 10428 15328 10659 15330
rect 10428 15272 10598 15328
rect 10654 15272 10659 15328
rect 10428 15270 10659 15272
rect 10428 15268 10434 15270
rect 10593 15267 10659 15270
rect 10726 15268 10732 15332
rect 10796 15330 10802 15332
rect 10961 15330 11027 15333
rect 10796 15328 11027 15330
rect 10796 15272 10966 15328
rect 11022 15272 11027 15328
rect 10796 15270 11027 15272
rect 10796 15268 10802 15270
rect 10961 15267 11027 15270
rect 20897 15330 20963 15333
rect 23841 15330 23907 15333
rect 20897 15328 23907 15330
rect 20897 15272 20902 15328
rect 20958 15272 23846 15328
rect 23902 15272 23907 15328
rect 20897 15270 23907 15272
rect 20897 15267 20963 15270
rect 23841 15267 23907 15270
rect 4246 15264 4562 15265
rect 4246 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4562 15264
rect 4246 15199 4562 15200
rect 11951 15264 12267 15265
rect 11951 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12267 15264
rect 11951 15199 12267 15200
rect 19656 15264 19972 15265
rect 19656 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19972 15264
rect 19656 15199 19972 15200
rect 27361 15264 27677 15265
rect 27361 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27677 15264
rect 27361 15199 27677 15200
rect 7833 15194 7899 15197
rect 9990 15194 9996 15196
rect 7833 15192 9996 15194
rect 7833 15136 7838 15192
rect 7894 15136 9996 15192
rect 7833 15134 9996 15136
rect 7833 15131 7899 15134
rect 9990 15132 9996 15134
rect 10060 15132 10066 15196
rect 10133 15194 10199 15197
rect 10409 15194 10475 15197
rect 10133 15192 10475 15194
rect 10133 15136 10138 15192
rect 10194 15136 10414 15192
rect 10470 15136 10475 15192
rect 10133 15134 10475 15136
rect 10133 15131 10199 15134
rect 10409 15131 10475 15134
rect 12617 15192 12683 15197
rect 12617 15136 12622 15192
rect 12678 15136 12683 15192
rect 12617 15131 12683 15136
rect 21449 15194 21515 15197
rect 24669 15194 24735 15197
rect 21449 15192 24735 15194
rect 21449 15136 21454 15192
rect 21510 15136 24674 15192
rect 24730 15136 24735 15192
rect 21449 15134 24735 15136
rect 21449 15131 21515 15134
rect 24669 15131 24735 15134
rect 9857 15060 9923 15061
rect 9806 14996 9812 15060
rect 9876 15058 9923 15060
rect 10133 15058 10199 15061
rect 12620 15058 12680 15131
rect 9876 15056 9968 15058
rect 9918 15000 9968 15056
rect 9876 14998 9968 15000
rect 10133 15056 12680 15058
rect 10133 15000 10138 15056
rect 10194 15000 12680 15056
rect 10133 14998 12680 15000
rect 18597 15058 18663 15061
rect 24577 15058 24643 15061
rect 18597 15056 24643 15058
rect 18597 15000 18602 15056
rect 18658 15000 24582 15056
rect 24638 15000 24643 15056
rect 18597 14998 24643 15000
rect 9876 14996 9923 14998
rect 9857 14995 9923 14996
rect 10133 14995 10199 14998
rect 18597 14995 18663 14998
rect 24577 14995 24643 14998
rect 28257 15058 28323 15061
rect 31600 15058 32000 15088
rect 28257 15056 32000 15058
rect 28257 15000 28262 15056
rect 28318 15000 32000 15056
rect 28257 14998 32000 15000
rect 28257 14995 28323 14998
rect 31600 14968 32000 14998
rect 8661 14922 8727 14925
rect 9305 14922 9371 14925
rect 8661 14920 9371 14922
rect 8661 14864 8666 14920
rect 8722 14864 9310 14920
rect 9366 14864 9371 14920
rect 8661 14862 9371 14864
rect 8661 14859 8727 14862
rect 9305 14859 9371 14862
rect 9765 14922 9831 14925
rect 11145 14922 11211 14925
rect 9765 14920 11211 14922
rect 9765 14864 9770 14920
rect 9826 14864 11150 14920
rect 11206 14864 11211 14920
rect 9765 14862 11211 14864
rect 9765 14859 9831 14862
rect 11145 14859 11211 14862
rect 11329 14922 11395 14925
rect 12985 14922 13051 14925
rect 11329 14920 13051 14922
rect 11329 14864 11334 14920
rect 11390 14864 12990 14920
rect 13046 14864 13051 14920
rect 11329 14862 13051 14864
rect 11329 14859 11395 14862
rect 12985 14859 13051 14862
rect 22737 14922 22803 14925
rect 24761 14922 24827 14925
rect 22737 14920 24827 14922
rect 22737 14864 22742 14920
rect 22798 14864 24766 14920
rect 24822 14864 24827 14920
rect 22737 14862 24827 14864
rect 22737 14859 22803 14862
rect 24761 14859 24827 14862
rect 10542 14724 10548 14788
rect 10612 14786 10618 14788
rect 10685 14786 10751 14789
rect 10612 14784 10751 14786
rect 10612 14728 10690 14784
rect 10746 14728 10751 14784
rect 10612 14726 10751 14728
rect 10612 14724 10618 14726
rect 10685 14723 10751 14726
rect 8098 14720 8414 14721
rect 8098 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8414 14720
rect 8098 14655 8414 14656
rect 15803 14720 16119 14721
rect 15803 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16119 14720
rect 15803 14655 16119 14656
rect 23508 14720 23824 14721
rect 23508 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23824 14720
rect 23508 14655 23824 14656
rect 31213 14720 31529 14721
rect 31213 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31529 14720
rect 31213 14655 31529 14656
rect 21541 14650 21607 14653
rect 23197 14650 23263 14653
rect 21541 14648 23263 14650
rect 21541 14592 21546 14648
rect 21602 14592 23202 14648
rect 23258 14592 23263 14648
rect 21541 14590 23263 14592
rect 21541 14587 21607 14590
rect 23197 14587 23263 14590
rect 7649 14514 7715 14517
rect 10409 14514 10475 14517
rect 10869 14514 10935 14517
rect 7649 14512 10935 14514
rect 7649 14456 7654 14512
rect 7710 14456 10414 14512
rect 10470 14456 10874 14512
rect 10930 14456 10935 14512
rect 7649 14454 10935 14456
rect 7649 14451 7715 14454
rect 10409 14451 10475 14454
rect 10869 14451 10935 14454
rect 22461 14514 22527 14517
rect 25497 14514 25563 14517
rect 22461 14512 25563 14514
rect 22461 14456 22466 14512
rect 22522 14456 25502 14512
rect 25558 14456 25563 14512
rect 22461 14454 25563 14456
rect 22461 14451 22527 14454
rect 25497 14451 25563 14454
rect 22001 14378 22067 14381
rect 24485 14378 24551 14381
rect 22001 14376 24551 14378
rect 22001 14320 22006 14376
rect 22062 14320 24490 14376
rect 24546 14320 24551 14376
rect 22001 14318 24551 14320
rect 22001 14315 22067 14318
rect 24485 14315 24551 14318
rect 28257 14378 28323 14381
rect 31600 14378 32000 14408
rect 28257 14376 32000 14378
rect 28257 14320 28262 14376
rect 28318 14320 32000 14376
rect 28257 14318 32000 14320
rect 28257 14315 28323 14318
rect 31600 14288 32000 14318
rect 24945 14242 25011 14245
rect 26141 14242 26207 14245
rect 24945 14240 26207 14242
rect 24945 14184 24950 14240
rect 25006 14184 26146 14240
rect 26202 14184 26207 14240
rect 24945 14182 26207 14184
rect 24945 14179 25011 14182
rect 26141 14179 26207 14182
rect 4246 14176 4562 14177
rect 4246 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4562 14176
rect 4246 14111 4562 14112
rect 11951 14176 12267 14177
rect 11951 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12267 14176
rect 11951 14111 12267 14112
rect 19656 14176 19972 14177
rect 19656 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19972 14176
rect 19656 14111 19972 14112
rect 27361 14176 27677 14177
rect 27361 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27677 14176
rect 27361 14111 27677 14112
rect 23289 14106 23355 14109
rect 25957 14106 26023 14109
rect 23289 14104 26023 14106
rect 23289 14048 23294 14104
rect 23350 14048 25962 14104
rect 26018 14048 26023 14104
rect 23289 14046 26023 14048
rect 23289 14043 23355 14046
rect 25957 14043 26023 14046
rect 12157 13970 12223 13973
rect 15009 13970 15075 13973
rect 12157 13968 15075 13970
rect 12157 13912 12162 13968
rect 12218 13912 15014 13968
rect 15070 13912 15075 13968
rect 12157 13910 15075 13912
rect 12157 13907 12223 13910
rect 15009 13907 15075 13910
rect 21633 13970 21699 13973
rect 24669 13970 24735 13973
rect 25681 13970 25747 13973
rect 21633 13968 24735 13970
rect 21633 13912 21638 13968
rect 21694 13912 24674 13968
rect 24730 13912 24735 13968
rect 21633 13910 24735 13912
rect 21633 13907 21699 13910
rect 24669 13907 24735 13910
rect 24810 13968 25747 13970
rect 24810 13912 25686 13968
rect 25742 13912 25747 13968
rect 24810 13910 25747 13912
rect 10961 13834 11027 13837
rect 12065 13834 12131 13837
rect 10961 13832 12131 13834
rect 10961 13776 10966 13832
rect 11022 13776 12070 13832
rect 12126 13776 12131 13832
rect 10961 13774 12131 13776
rect 10961 13771 11027 13774
rect 12065 13771 12131 13774
rect 20437 13834 20503 13837
rect 23841 13834 23907 13837
rect 20437 13832 23907 13834
rect 20437 13776 20442 13832
rect 20498 13776 23846 13832
rect 23902 13776 23907 13832
rect 20437 13774 23907 13776
rect 20437 13771 20503 13774
rect 23841 13771 23907 13774
rect 9581 13698 9647 13701
rect 12893 13698 12959 13701
rect 9581 13696 12959 13698
rect 9581 13640 9586 13696
rect 9642 13640 12898 13696
rect 12954 13640 12959 13696
rect 9581 13638 12959 13640
rect 9581 13635 9647 13638
rect 12893 13635 12959 13638
rect 19057 13698 19123 13701
rect 22318 13698 22324 13700
rect 19057 13696 22324 13698
rect 19057 13640 19062 13696
rect 19118 13640 22324 13696
rect 19057 13638 22324 13640
rect 19057 13635 19123 13638
rect 22318 13636 22324 13638
rect 22388 13636 22394 13700
rect 24485 13698 24551 13701
rect 24810 13698 24870 13910
rect 25681 13907 25747 13910
rect 24485 13696 24870 13698
rect 24485 13640 24490 13696
rect 24546 13640 24870 13696
rect 24485 13638 24870 13640
rect 31600 13696 32000 13728
rect 31600 13640 31666 13696
rect 31722 13640 32000 13696
rect 24485 13635 24551 13638
rect 8098 13632 8414 13633
rect 8098 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8414 13632
rect 8098 13567 8414 13568
rect 15803 13632 16119 13633
rect 15803 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16119 13632
rect 15803 13567 16119 13568
rect 23508 13632 23824 13633
rect 23508 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23824 13632
rect 23508 13567 23824 13568
rect 31213 13632 31529 13633
rect 31213 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31529 13632
rect 31600 13608 32000 13640
rect 31213 13567 31529 13568
rect 9305 13562 9371 13565
rect 12433 13562 12499 13565
rect 9305 13560 12499 13562
rect 9305 13504 9310 13560
rect 9366 13504 12438 13560
rect 12494 13504 12499 13560
rect 9305 13502 12499 13504
rect 9305 13499 9371 13502
rect 12433 13499 12499 13502
rect 24577 13562 24643 13565
rect 25497 13562 25563 13565
rect 24577 13560 25563 13562
rect 24577 13504 24582 13560
rect 24638 13504 25502 13560
rect 25558 13504 25563 13560
rect 24577 13502 25563 13504
rect 24577 13499 24643 13502
rect 25497 13499 25563 13502
rect 7649 13426 7715 13429
rect 11094 13426 11100 13428
rect 7649 13424 11100 13426
rect 7649 13368 7654 13424
rect 7710 13368 11100 13424
rect 7649 13366 11100 13368
rect 7649 13363 7715 13366
rect 11094 13364 11100 13366
rect 11164 13364 11170 13428
rect 21950 13364 21956 13428
rect 22020 13426 22026 13428
rect 25313 13426 25379 13429
rect 22020 13424 25379 13426
rect 22020 13368 25318 13424
rect 25374 13368 25379 13424
rect 22020 13366 25379 13368
rect 22020 13364 22026 13366
rect 25313 13363 25379 13366
rect 7925 13290 7991 13293
rect 9213 13290 9279 13293
rect 7925 13288 9279 13290
rect 7925 13232 7930 13288
rect 7986 13232 9218 13288
rect 9274 13232 9279 13288
rect 7925 13230 9279 13232
rect 7925 13227 7991 13230
rect 9213 13227 9279 13230
rect 23289 13290 23355 13293
rect 26693 13290 26759 13293
rect 23289 13288 26759 13290
rect 23289 13232 23294 13288
rect 23350 13232 26698 13288
rect 26754 13232 26759 13288
rect 23289 13230 26759 13232
rect 23289 13227 23355 13230
rect 26693 13227 26759 13230
rect 21173 13154 21239 13157
rect 24485 13154 24551 13157
rect 21173 13152 24551 13154
rect 21173 13096 21178 13152
rect 21234 13096 24490 13152
rect 24546 13096 24551 13152
rect 21173 13094 24551 13096
rect 21173 13091 21239 13094
rect 24485 13091 24551 13094
rect 24853 13156 24919 13157
rect 24853 13152 24900 13156
rect 24964 13154 24970 13156
rect 24853 13096 24858 13152
rect 24853 13092 24900 13096
rect 24964 13094 25010 13154
rect 24964 13092 24970 13094
rect 24853 13091 24919 13092
rect 4246 13088 4562 13089
rect 0 13018 400 13048
rect 4246 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4562 13088
rect 4246 13023 4562 13024
rect 11951 13088 12267 13089
rect 11951 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12267 13088
rect 11951 13023 12267 13024
rect 19656 13088 19972 13089
rect 19656 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19972 13088
rect 19656 13023 19972 13024
rect 27361 13088 27677 13089
rect 27361 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27677 13088
rect 27361 13023 27677 13024
rect 11329 13020 11395 13021
rect 11697 13020 11763 13021
rect 0 12958 2790 13018
rect 0 12928 400 12958
rect 2730 12882 2790 12958
rect 11278 12956 11284 13020
rect 11348 13018 11395 13020
rect 11348 13016 11440 13018
rect 11390 12960 11440 13016
rect 11348 12958 11440 12960
rect 11348 12956 11395 12958
rect 11646 12956 11652 13020
rect 11716 13018 11763 13020
rect 28257 13018 28323 13021
rect 31600 13018 32000 13048
rect 11716 13016 11808 13018
rect 11758 12960 11808 13016
rect 11716 12958 11808 12960
rect 28257 13016 32000 13018
rect 28257 12960 28262 13016
rect 28318 12960 32000 13016
rect 28257 12958 32000 12960
rect 11716 12956 11763 12958
rect 11329 12955 11395 12956
rect 11697 12955 11763 12956
rect 28257 12955 28323 12958
rect 31600 12928 32000 12958
rect 8937 12882 9003 12885
rect 2730 12880 9003 12882
rect 2730 12824 8942 12880
rect 8998 12824 9003 12880
rect 2730 12822 9003 12824
rect 8937 12819 9003 12822
rect 23238 12820 23244 12884
rect 23308 12882 23314 12884
rect 25589 12882 25655 12885
rect 23308 12880 25655 12882
rect 23308 12824 25594 12880
rect 25650 12824 25655 12880
rect 23308 12822 25655 12824
rect 23308 12820 23314 12822
rect 25589 12819 25655 12822
rect 23657 12746 23723 12749
rect 26141 12746 26207 12749
rect 23657 12744 26207 12746
rect 23657 12688 23662 12744
rect 23718 12688 26146 12744
rect 26202 12688 26207 12744
rect 23657 12686 26207 12688
rect 23657 12683 23723 12686
rect 26141 12683 26207 12686
rect 8098 12544 8414 12545
rect 8098 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8414 12544
rect 8098 12479 8414 12480
rect 15803 12544 16119 12545
rect 15803 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16119 12544
rect 15803 12479 16119 12480
rect 23508 12544 23824 12545
rect 23508 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23824 12544
rect 23508 12479 23824 12480
rect 31213 12544 31529 12545
rect 31213 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31529 12544
rect 31213 12479 31529 12480
rect 10041 12338 10107 12341
rect 13077 12338 13143 12341
rect 10041 12336 13143 12338
rect 10041 12280 10046 12336
rect 10102 12280 13082 12336
rect 13138 12280 13143 12336
rect 10041 12278 13143 12280
rect 10041 12275 10107 12278
rect 13077 12275 13143 12278
rect 18505 12338 18571 12341
rect 23974 12338 23980 12340
rect 18505 12336 23980 12338
rect 18505 12280 18510 12336
rect 18566 12280 23980 12336
rect 18505 12278 23980 12280
rect 18505 12275 18571 12278
rect 23974 12276 23980 12278
rect 24044 12276 24050 12340
rect 28257 12338 28323 12341
rect 31600 12338 32000 12368
rect 28257 12336 32000 12338
rect 28257 12280 28262 12336
rect 28318 12280 32000 12336
rect 28257 12278 32000 12280
rect 28257 12275 28323 12278
rect 31600 12248 32000 12278
rect 20345 12066 20411 12069
rect 25221 12066 25287 12069
rect 20345 12064 25287 12066
rect 20345 12008 20350 12064
rect 20406 12008 25226 12064
rect 25282 12008 25287 12064
rect 20345 12006 25287 12008
rect 20345 12003 20411 12006
rect 25221 12003 25287 12006
rect 4246 12000 4562 12001
rect 4246 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4562 12000
rect 4246 11935 4562 11936
rect 11951 12000 12267 12001
rect 11951 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12267 12000
rect 11951 11935 12267 11936
rect 19656 12000 19972 12001
rect 19656 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19972 12000
rect 19656 11935 19972 11936
rect 27361 12000 27677 12001
rect 27361 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27677 12000
rect 27361 11935 27677 11936
rect 15377 11930 15443 11933
rect 17125 11930 17191 11933
rect 15377 11928 17191 11930
rect 15377 11872 15382 11928
rect 15438 11872 17130 11928
rect 17186 11872 17191 11928
rect 15377 11870 17191 11872
rect 15377 11867 15443 11870
rect 17125 11867 17191 11870
rect 15193 11794 15259 11797
rect 15653 11794 15719 11797
rect 15193 11792 15719 11794
rect 15193 11736 15198 11792
rect 15254 11736 15658 11792
rect 15714 11736 15719 11792
rect 15193 11734 15719 11736
rect 15193 11731 15259 11734
rect 15653 11731 15719 11734
rect 15837 11794 15903 11797
rect 18229 11794 18295 11797
rect 15837 11792 18295 11794
rect 15837 11736 15842 11792
rect 15898 11736 18234 11792
rect 18290 11736 18295 11792
rect 15837 11734 18295 11736
rect 15837 11731 15903 11734
rect 18229 11731 18295 11734
rect 19333 11796 19399 11797
rect 19333 11792 19380 11796
rect 19444 11794 19450 11796
rect 23289 11794 23355 11797
rect 29637 11794 29703 11797
rect 19333 11736 19338 11792
rect 19333 11732 19380 11736
rect 19444 11734 19490 11794
rect 23289 11792 29703 11794
rect 23289 11736 23294 11792
rect 23350 11736 29642 11792
rect 29698 11736 29703 11792
rect 23289 11734 29703 11736
rect 19444 11732 19450 11734
rect 19333 11731 19399 11732
rect 23289 11731 23355 11734
rect 29637 11731 29703 11734
rect 14917 11658 14983 11661
rect 19425 11658 19491 11661
rect 14917 11656 19491 11658
rect 14917 11600 14922 11656
rect 14978 11600 19430 11656
rect 19486 11600 19491 11656
rect 14917 11598 19491 11600
rect 14917 11595 14983 11598
rect 19425 11595 19491 11598
rect 24485 11658 24551 11661
rect 25957 11658 26023 11661
rect 24485 11656 26023 11658
rect 24485 11600 24490 11656
rect 24546 11600 25962 11656
rect 26018 11600 26023 11656
rect 24485 11598 26023 11600
rect 24485 11595 24551 11598
rect 25957 11595 26023 11598
rect 28257 11658 28323 11661
rect 31600 11658 32000 11688
rect 28257 11656 32000 11658
rect 28257 11600 28262 11656
rect 28318 11600 32000 11656
rect 28257 11598 32000 11600
rect 28257 11595 28323 11598
rect 31600 11568 32000 11598
rect 8098 11456 8414 11457
rect 8098 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8414 11456
rect 8098 11391 8414 11392
rect 15803 11456 16119 11457
rect 15803 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16119 11456
rect 15803 11391 16119 11392
rect 23508 11456 23824 11457
rect 23508 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23824 11456
rect 23508 11391 23824 11392
rect 31213 11456 31529 11457
rect 31213 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31529 11456
rect 31213 11391 31529 11392
rect 9489 11250 9555 11253
rect 16113 11250 16179 11253
rect 9489 11248 16179 11250
rect 9489 11192 9494 11248
rect 9550 11192 16118 11248
rect 16174 11192 16179 11248
rect 9489 11190 16179 11192
rect 9489 11187 9555 11190
rect 16113 11187 16179 11190
rect 14825 11114 14891 11117
rect 16481 11114 16547 11117
rect 14825 11112 16547 11114
rect 14825 11056 14830 11112
rect 14886 11056 16486 11112
rect 16542 11056 16547 11112
rect 14825 11054 16547 11056
rect 14825 11051 14891 11054
rect 16481 11051 16547 11054
rect 0 10978 400 11008
rect 13261 10980 13327 10981
rect 13261 10978 13308 10980
rect 0 10918 2790 10978
rect 13216 10976 13308 10978
rect 13216 10920 13266 10976
rect 13216 10918 13308 10920
rect 0 10888 400 10918
rect 2730 10706 2790 10918
rect 13261 10916 13308 10918
rect 13372 10916 13378 10980
rect 28257 10978 28323 10981
rect 31600 10978 32000 11008
rect 28257 10976 32000 10978
rect 28257 10920 28262 10976
rect 28318 10920 32000 10976
rect 28257 10918 32000 10920
rect 13261 10915 13327 10916
rect 28257 10915 28323 10918
rect 4246 10912 4562 10913
rect 4246 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4562 10912
rect 4246 10847 4562 10848
rect 11951 10912 12267 10913
rect 11951 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12267 10912
rect 11951 10847 12267 10848
rect 19656 10912 19972 10913
rect 19656 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19972 10912
rect 19656 10847 19972 10848
rect 27361 10912 27677 10913
rect 27361 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27677 10912
rect 31600 10888 32000 10918
rect 27361 10847 27677 10848
rect 10225 10706 10291 10709
rect 2730 10704 10291 10706
rect 2730 10648 10230 10704
rect 10286 10648 10291 10704
rect 2730 10646 10291 10648
rect 10225 10643 10291 10646
rect 15653 10432 15719 10437
rect 15653 10376 15658 10432
rect 15714 10376 15719 10432
rect 15653 10371 15719 10376
rect 8098 10368 8414 10369
rect 0 10298 400 10328
rect 8098 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8414 10368
rect 8098 10303 8414 10304
rect 0 10238 2790 10298
rect 0 10208 400 10238
rect 2730 10162 2790 10238
rect 9121 10162 9187 10165
rect 2730 10160 9187 10162
rect 2730 10104 9126 10160
rect 9182 10104 9187 10160
rect 2730 10102 9187 10104
rect 15656 10162 15716 10371
rect 15803 10368 16119 10369
rect 15803 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16119 10368
rect 15803 10303 16119 10304
rect 23508 10368 23824 10369
rect 23508 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23824 10368
rect 23508 10303 23824 10304
rect 31213 10368 31529 10369
rect 31213 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31529 10368
rect 31213 10303 31529 10304
rect 31600 10296 32000 10328
rect 31600 10240 31666 10296
rect 31722 10240 32000 10296
rect 31600 10208 32000 10240
rect 15929 10162 15995 10165
rect 15656 10160 15995 10162
rect 15656 10104 15934 10160
rect 15990 10104 15995 10160
rect 15656 10102 15995 10104
rect 9121 10099 9187 10102
rect 15929 10099 15995 10102
rect 15469 10026 15535 10029
rect 15837 10026 15903 10029
rect 15469 10024 15903 10026
rect 15469 9968 15474 10024
rect 15530 9968 15842 10024
rect 15898 9968 15903 10024
rect 15469 9966 15903 9968
rect 15469 9963 15535 9966
rect 15837 9963 15903 9966
rect 4246 9824 4562 9825
rect 4246 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4562 9824
rect 4246 9759 4562 9760
rect 11951 9824 12267 9825
rect 11951 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12267 9824
rect 11951 9759 12267 9760
rect 19656 9824 19972 9825
rect 19656 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19972 9824
rect 19656 9759 19972 9760
rect 27361 9824 27677 9825
rect 27361 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27677 9824
rect 27361 9759 27677 9760
rect 0 9618 400 9648
rect 8661 9618 8727 9621
rect 0 9616 8727 9618
rect 0 9560 8666 9616
rect 8722 9560 8727 9616
rect 0 9558 8727 9560
rect 0 9528 400 9558
rect 8661 9555 8727 9558
rect 15561 9618 15627 9621
rect 17953 9618 18019 9621
rect 15561 9616 18019 9618
rect 15561 9560 15566 9616
rect 15622 9560 17958 9616
rect 18014 9560 18019 9616
rect 15561 9558 18019 9560
rect 15561 9555 15627 9558
rect 17953 9555 18019 9558
rect 21357 9618 21423 9621
rect 24025 9618 24091 9621
rect 21357 9616 24091 9618
rect 21357 9560 21362 9616
rect 21418 9560 24030 9616
rect 24086 9560 24091 9616
rect 21357 9558 24091 9560
rect 21357 9555 21423 9558
rect 24025 9555 24091 9558
rect 28257 9618 28323 9621
rect 31600 9618 32000 9648
rect 28257 9616 32000 9618
rect 28257 9560 28262 9616
rect 28318 9560 32000 9616
rect 28257 9558 32000 9560
rect 28257 9555 28323 9558
rect 31600 9528 32000 9558
rect 6453 9482 6519 9485
rect 9765 9482 9831 9485
rect 6453 9480 9831 9482
rect 6453 9424 6458 9480
rect 6514 9424 9770 9480
rect 9826 9424 9831 9480
rect 6453 9422 9831 9424
rect 6453 9419 6519 9422
rect 9765 9419 9831 9422
rect 8098 9280 8414 9281
rect 8098 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8414 9280
rect 8098 9215 8414 9216
rect 15803 9280 16119 9281
rect 15803 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16119 9280
rect 15803 9215 16119 9216
rect 23508 9280 23824 9281
rect 23508 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23824 9280
rect 23508 9215 23824 9216
rect 31213 9280 31529 9281
rect 31213 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31529 9280
rect 31213 9215 31529 9216
rect 11329 9210 11395 9213
rect 13445 9210 13511 9213
rect 11329 9208 13511 9210
rect 11329 9152 11334 9208
rect 11390 9152 13450 9208
rect 13506 9152 13511 9208
rect 11329 9150 13511 9152
rect 11329 9147 11395 9150
rect 13445 9147 13511 9150
rect 12709 9074 12775 9077
rect 17769 9074 17835 9077
rect 19333 9074 19399 9077
rect 22369 9074 22435 9077
rect 12709 9072 22435 9074
rect 12709 9016 12714 9072
rect 12770 9016 17774 9072
rect 17830 9016 19338 9072
rect 19394 9016 22374 9072
rect 22430 9016 22435 9072
rect 12709 9014 22435 9016
rect 12709 9011 12775 9014
rect 17769 9011 17835 9014
rect 19333 9011 19399 9014
rect 22369 9011 22435 9014
rect 23289 8938 23355 8941
rect 31600 8938 32000 8968
rect 23289 8936 32000 8938
rect 23289 8880 23294 8936
rect 23350 8880 32000 8936
rect 23289 8878 32000 8880
rect 23289 8875 23355 8878
rect 31600 8848 32000 8878
rect 22001 8802 22067 8805
rect 23933 8802 23999 8805
rect 22001 8800 23999 8802
rect 22001 8744 22006 8800
rect 22062 8744 23938 8800
rect 23994 8744 23999 8800
rect 22001 8742 23999 8744
rect 22001 8739 22067 8742
rect 23933 8739 23999 8742
rect 4246 8736 4562 8737
rect 4246 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4562 8736
rect 4246 8671 4562 8672
rect 11951 8736 12267 8737
rect 11951 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12267 8736
rect 11951 8671 12267 8672
rect 19656 8736 19972 8737
rect 19656 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19972 8736
rect 19656 8671 19972 8672
rect 27361 8736 27677 8737
rect 27361 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27677 8736
rect 27361 8671 27677 8672
rect 22829 8530 22895 8533
rect 25589 8530 25655 8533
rect 31661 8530 31727 8533
rect 22829 8528 24870 8530
rect 22829 8472 22834 8528
rect 22890 8472 24870 8528
rect 22829 8470 24870 8472
rect 22829 8467 22895 8470
rect 6729 8394 6795 8397
rect 9765 8394 9831 8397
rect 15193 8396 15259 8397
rect 15142 8394 15148 8396
rect 6729 8392 9831 8394
rect 6729 8336 6734 8392
rect 6790 8336 9770 8392
rect 9826 8336 9831 8392
rect 6729 8334 9831 8336
rect 15102 8334 15148 8394
rect 15212 8392 15259 8396
rect 15254 8336 15259 8392
rect 6729 8331 6795 8334
rect 9765 8331 9831 8334
rect 15142 8332 15148 8334
rect 15212 8332 15259 8336
rect 15193 8331 15259 8332
rect 20161 8394 20227 8397
rect 20662 8394 20668 8396
rect 20161 8392 20668 8394
rect 20161 8336 20166 8392
rect 20222 8336 20668 8392
rect 20161 8334 20668 8336
rect 20161 8331 20227 8334
rect 20662 8332 20668 8334
rect 20732 8332 20738 8396
rect 21909 8394 21975 8397
rect 24810 8394 24870 8470
rect 25589 8528 31727 8530
rect 25589 8472 25594 8528
rect 25650 8472 31666 8528
rect 31722 8472 31727 8528
rect 25589 8470 31727 8472
rect 25589 8467 25655 8470
rect 31661 8467 31727 8470
rect 21909 8392 24594 8394
rect 21909 8336 21914 8392
rect 21970 8336 24594 8392
rect 21909 8334 24594 8336
rect 24810 8334 28090 8394
rect 21909 8331 21975 8334
rect 0 8258 400 8288
rect 24534 8258 24594 8334
rect 24669 8258 24735 8261
rect 0 8198 2790 8258
rect 24534 8256 24735 8258
rect 24534 8200 24674 8256
rect 24730 8200 24735 8256
rect 24534 8198 24735 8200
rect 0 8168 400 8198
rect 2730 7986 2790 8198
rect 24669 8195 24735 8198
rect 8098 8192 8414 8193
rect 8098 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8414 8192
rect 8098 8127 8414 8128
rect 15803 8192 16119 8193
rect 15803 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16119 8192
rect 15803 8127 16119 8128
rect 23508 8192 23824 8193
rect 23508 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23824 8192
rect 23508 8127 23824 8128
rect 8845 7986 8911 7989
rect 2730 7984 8911 7986
rect 2730 7928 8850 7984
rect 8906 7928 8911 7984
rect 2730 7926 8911 7928
rect 8845 7923 8911 7926
rect 23749 7714 23815 7717
rect 25589 7714 25655 7717
rect 23749 7712 25655 7714
rect 23749 7656 23754 7712
rect 23810 7656 25594 7712
rect 25650 7656 25655 7712
rect 23749 7654 25655 7656
rect 23749 7651 23815 7654
rect 25589 7651 25655 7654
rect 4246 7648 4562 7649
rect 4246 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4562 7648
rect 4246 7583 4562 7584
rect 11951 7648 12267 7649
rect 11951 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12267 7648
rect 11951 7583 12267 7584
rect 19656 7648 19972 7649
rect 19656 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19972 7648
rect 19656 7583 19972 7584
rect 27361 7648 27677 7649
rect 27361 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27677 7648
rect 27361 7583 27677 7584
rect 24209 7578 24275 7581
rect 26325 7578 26391 7581
rect 24209 7576 26391 7578
rect 24209 7520 24214 7576
rect 24270 7520 26330 7576
rect 26386 7520 26391 7576
rect 24209 7518 26391 7520
rect 28030 7578 28090 8334
rect 31600 8256 32000 8288
rect 31600 8200 31666 8256
rect 31722 8200 32000 8256
rect 31213 8192 31529 8193
rect 31213 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31529 8192
rect 31600 8168 32000 8200
rect 31213 8127 31529 8128
rect 31600 7578 32000 7608
rect 28030 7518 32000 7578
rect 24209 7515 24275 7518
rect 26325 7515 26391 7518
rect 31600 7488 32000 7518
rect 7005 7442 7071 7445
rect 10133 7442 10199 7445
rect 7005 7440 10199 7442
rect 7005 7384 7010 7440
rect 7066 7384 10138 7440
rect 10194 7384 10199 7440
rect 7005 7382 10199 7384
rect 7005 7379 7071 7382
rect 10133 7379 10199 7382
rect 9213 7306 9279 7309
rect 9581 7306 9647 7309
rect 9213 7304 9647 7306
rect 9213 7248 9218 7304
rect 9274 7248 9586 7304
rect 9642 7248 9647 7304
rect 9213 7246 9647 7248
rect 9213 7243 9279 7246
rect 9581 7243 9647 7246
rect 19701 7306 19767 7309
rect 20161 7306 20227 7309
rect 31661 7306 31727 7309
rect 19701 7304 20227 7306
rect 19701 7248 19706 7304
rect 19762 7248 20166 7304
rect 20222 7248 20227 7304
rect 19701 7246 20227 7248
rect 19701 7243 19767 7246
rect 20161 7243 20227 7246
rect 23200 7304 31727 7306
rect 23200 7248 31666 7304
rect 31722 7248 31727 7304
rect 23200 7246 31727 7248
rect 23200 7173 23260 7246
rect 31661 7243 31727 7246
rect 14825 7170 14891 7173
rect 15469 7170 15535 7173
rect 14825 7168 15535 7170
rect 14825 7112 14830 7168
rect 14886 7112 15474 7168
rect 15530 7112 15535 7168
rect 14825 7110 15535 7112
rect 14825 7107 14891 7110
rect 15469 7107 15535 7110
rect 23197 7168 23263 7173
rect 23197 7112 23202 7168
rect 23258 7112 23263 7168
rect 23197 7107 23263 7112
rect 24485 7170 24551 7173
rect 25957 7170 26023 7173
rect 24485 7168 26023 7170
rect 24485 7112 24490 7168
rect 24546 7112 25962 7168
rect 26018 7112 26023 7168
rect 24485 7110 26023 7112
rect 24485 7107 24551 7110
rect 25957 7107 26023 7110
rect 8098 7104 8414 7105
rect 8098 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8414 7104
rect 8098 7039 8414 7040
rect 15803 7104 16119 7105
rect 15803 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16119 7104
rect 15803 7039 16119 7040
rect 23508 7104 23824 7105
rect 23508 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23824 7104
rect 23508 7039 23824 7040
rect 31213 7104 31529 7105
rect 31213 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31529 7104
rect 31213 7039 31529 7040
rect 11513 7034 11579 7037
rect 11513 7032 15394 7034
rect 11513 6976 11518 7032
rect 11574 6976 15394 7032
rect 11513 6974 15394 6976
rect 11513 6971 11579 6974
rect 15334 6901 15394 6974
rect 7649 6898 7715 6901
rect 10317 6898 10383 6901
rect 7649 6896 10383 6898
rect 7649 6840 7654 6896
rect 7710 6840 10322 6896
rect 10378 6840 10383 6896
rect 7649 6838 10383 6840
rect 15334 6896 15443 6901
rect 15334 6840 15382 6896
rect 15438 6840 15443 6896
rect 15334 6838 15443 6840
rect 7649 6835 7715 6838
rect 10317 6835 10383 6838
rect 15377 6835 15443 6838
rect 22645 6898 22711 6901
rect 24117 6898 24183 6901
rect 22645 6896 24183 6898
rect 22645 6840 22650 6896
rect 22706 6840 24122 6896
rect 24178 6840 24183 6896
rect 22645 6838 24183 6840
rect 22645 6835 22711 6838
rect 24117 6835 24183 6838
rect 25589 6898 25655 6901
rect 31600 6898 32000 6928
rect 25589 6896 32000 6898
rect 25589 6840 25594 6896
rect 25650 6840 32000 6896
rect 25589 6838 32000 6840
rect 25589 6835 25655 6838
rect 31600 6808 32000 6838
rect 23105 6762 23171 6765
rect 25037 6762 25103 6765
rect 23105 6760 25103 6762
rect 23105 6704 23110 6760
rect 23166 6704 25042 6760
rect 25098 6704 25103 6760
rect 23105 6702 25103 6704
rect 23105 6699 23171 6702
rect 25037 6699 25103 6702
rect 22001 6626 22067 6629
rect 24761 6626 24827 6629
rect 22001 6624 24827 6626
rect 22001 6568 22006 6624
rect 22062 6568 24766 6624
rect 24822 6568 24827 6624
rect 22001 6566 24827 6568
rect 22001 6563 22067 6566
rect 24761 6563 24827 6566
rect 4246 6560 4562 6561
rect 4246 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4562 6560
rect 4246 6495 4562 6496
rect 11951 6560 12267 6561
rect 11951 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12267 6560
rect 11951 6495 12267 6496
rect 19656 6560 19972 6561
rect 19656 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19972 6560
rect 19656 6495 19972 6496
rect 27361 6560 27677 6561
rect 27361 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27677 6560
rect 27361 6495 27677 6496
rect 21633 6354 21699 6357
rect 23473 6354 23539 6357
rect 21633 6352 23539 6354
rect 21633 6296 21638 6352
rect 21694 6296 23478 6352
rect 23534 6296 23539 6352
rect 21633 6294 23539 6296
rect 21633 6291 21699 6294
rect 23473 6291 23539 6294
rect 9029 6218 9095 6221
rect 9765 6218 9831 6221
rect 9029 6216 9831 6218
rect 9029 6160 9034 6216
rect 9090 6160 9770 6216
rect 9826 6160 9831 6216
rect 9029 6158 9831 6160
rect 9029 6155 9095 6158
rect 9765 6155 9831 6158
rect 18873 6218 18939 6221
rect 19241 6218 19307 6221
rect 18873 6216 19307 6218
rect 18873 6160 18878 6216
rect 18934 6160 19246 6216
rect 19302 6160 19307 6216
rect 18873 6158 19307 6160
rect 18873 6155 18939 6158
rect 19241 6155 19307 6158
rect 21725 6218 21791 6221
rect 22277 6218 22343 6221
rect 21725 6216 22343 6218
rect 21725 6160 21730 6216
rect 21786 6160 22282 6216
rect 22338 6160 22343 6216
rect 21725 6158 22343 6160
rect 21725 6155 21791 6158
rect 22277 6155 22343 6158
rect 22645 6218 22711 6221
rect 31600 6218 32000 6248
rect 22645 6216 32000 6218
rect 22645 6160 22650 6216
rect 22706 6160 32000 6216
rect 22645 6158 32000 6160
rect 22645 6155 22711 6158
rect 31600 6128 32000 6158
rect 21909 6082 21975 6085
rect 23105 6082 23171 6085
rect 21909 6080 23171 6082
rect 21909 6024 21914 6080
rect 21970 6024 23110 6080
rect 23166 6024 23171 6080
rect 21909 6022 23171 6024
rect 21909 6019 21975 6022
rect 23105 6019 23171 6022
rect 8098 6016 8414 6017
rect 8098 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8414 6016
rect 8098 5951 8414 5952
rect 15803 6016 16119 6017
rect 15803 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16119 6016
rect 15803 5951 16119 5952
rect 23508 6016 23824 6017
rect 23508 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23824 6016
rect 23508 5951 23824 5952
rect 31213 6016 31529 6017
rect 31213 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31529 6016
rect 31213 5951 31529 5952
rect 20069 5946 20135 5949
rect 22461 5946 22527 5949
rect 20069 5944 22527 5946
rect 20069 5888 20074 5944
rect 20130 5888 22466 5944
rect 22522 5888 22527 5944
rect 20069 5886 22527 5888
rect 20069 5883 20135 5886
rect 22461 5883 22527 5886
rect 20345 5810 20411 5813
rect 21541 5810 21607 5813
rect 20345 5808 21607 5810
rect 20345 5752 20350 5808
rect 20406 5752 21546 5808
rect 21602 5752 21607 5808
rect 20345 5750 21607 5752
rect 20345 5747 20411 5750
rect 21541 5747 21607 5750
rect 22001 5810 22067 5813
rect 23013 5810 23079 5813
rect 22001 5808 23079 5810
rect 22001 5752 22006 5808
rect 22062 5752 23018 5808
rect 23074 5752 23079 5808
rect 22001 5750 23079 5752
rect 22001 5747 22067 5750
rect 23013 5747 23079 5750
rect 19057 5674 19123 5677
rect 22185 5674 22251 5677
rect 19057 5672 22251 5674
rect 19057 5616 19062 5672
rect 19118 5616 22190 5672
rect 22246 5616 22251 5672
rect 19057 5614 22251 5616
rect 19057 5611 19123 5614
rect 22185 5611 22251 5614
rect 14549 5538 14615 5541
rect 15101 5538 15167 5541
rect 14549 5536 15167 5538
rect 14549 5480 14554 5536
rect 14610 5480 15106 5536
rect 15162 5480 15167 5536
rect 14549 5478 15167 5480
rect 14549 5475 14615 5478
rect 15101 5475 15167 5478
rect 20989 5538 21055 5541
rect 24025 5538 24091 5541
rect 31600 5538 32000 5568
rect 20989 5536 24091 5538
rect 20989 5480 20994 5536
rect 21050 5480 24030 5536
rect 24086 5480 24091 5536
rect 20989 5478 24091 5480
rect 20989 5475 21055 5478
rect 24025 5475 24091 5478
rect 28214 5478 32000 5538
rect 4246 5472 4562 5473
rect 4246 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4562 5472
rect 4246 5407 4562 5408
rect 11951 5472 12267 5473
rect 11951 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12267 5472
rect 11951 5407 12267 5408
rect 19656 5472 19972 5473
rect 19656 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19972 5472
rect 19656 5407 19972 5408
rect 27361 5472 27677 5473
rect 27361 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27677 5472
rect 27361 5407 27677 5408
rect 15009 5402 15075 5405
rect 14966 5400 15075 5402
rect 14966 5344 15014 5400
rect 15070 5344 15075 5400
rect 14966 5339 15075 5344
rect 21449 5402 21515 5405
rect 25129 5402 25195 5405
rect 21449 5400 25195 5402
rect 21449 5344 21454 5400
rect 21510 5344 25134 5400
rect 25190 5344 25195 5400
rect 21449 5342 25195 5344
rect 21449 5339 21515 5342
rect 25129 5339 25195 5342
rect 14966 4997 15026 5339
rect 20529 5266 20595 5269
rect 22277 5266 22343 5269
rect 20529 5264 22343 5266
rect 20529 5208 20534 5264
rect 20590 5208 22282 5264
rect 22338 5208 22343 5264
rect 20529 5206 22343 5208
rect 20529 5203 20595 5206
rect 22277 5203 22343 5206
rect 28214 5130 28274 5478
rect 31600 5448 32000 5478
rect 14917 4992 15026 4997
rect 14917 4936 14922 4992
rect 14978 4936 15026 4992
rect 14917 4934 15026 4936
rect 22050 5070 28274 5130
rect 14917 4931 14983 4934
rect 8098 4928 8414 4929
rect 8098 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8414 4928
rect 8098 4863 8414 4864
rect 15803 4928 16119 4929
rect 15803 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16119 4928
rect 15803 4863 16119 4864
rect 9305 4722 9371 4725
rect 10685 4722 10751 4725
rect 9305 4720 10751 4722
rect 9305 4664 9310 4720
rect 9366 4664 10690 4720
rect 10746 4664 10751 4720
rect 9305 4662 10751 4664
rect 9305 4659 9371 4662
rect 10685 4659 10751 4662
rect 20662 4524 20668 4588
rect 20732 4586 20738 4588
rect 22050 4586 22110 5070
rect 23508 4928 23824 4929
rect 23508 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23824 4928
rect 23508 4863 23824 4864
rect 31213 4928 31529 4929
rect 31213 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31529 4928
rect 31213 4863 31529 4864
rect 31600 4856 32000 4888
rect 31600 4800 31666 4856
rect 31722 4800 32000 4856
rect 31600 4768 32000 4800
rect 20732 4526 22110 4586
rect 20732 4524 20738 4526
rect 4246 4384 4562 4385
rect 4246 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4562 4384
rect 4246 4319 4562 4320
rect 11951 4384 12267 4385
rect 11951 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12267 4384
rect 11951 4319 12267 4320
rect 19656 4384 19972 4385
rect 19656 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19972 4384
rect 19656 4319 19972 4320
rect 27361 4384 27677 4385
rect 27361 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27677 4384
rect 27361 4319 27677 4320
rect 8098 3840 8414 3841
rect 8098 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8414 3840
rect 8098 3775 8414 3776
rect 15803 3840 16119 3841
rect 15803 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16119 3840
rect 15803 3775 16119 3776
rect 23508 3840 23824 3841
rect 23508 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23824 3840
rect 23508 3775 23824 3776
rect 31213 3840 31529 3841
rect 31213 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31529 3840
rect 31213 3775 31529 3776
rect 4246 3296 4562 3297
rect 4246 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4562 3296
rect 4246 3231 4562 3232
rect 11951 3296 12267 3297
rect 11951 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12267 3296
rect 11951 3231 12267 3232
rect 19656 3296 19972 3297
rect 19656 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19972 3296
rect 19656 3231 19972 3232
rect 27361 3296 27677 3297
rect 27361 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27677 3296
rect 27361 3231 27677 3232
rect 8098 2752 8414 2753
rect 8098 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8414 2752
rect 8098 2687 8414 2688
rect 15803 2752 16119 2753
rect 15803 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16119 2752
rect 15803 2687 16119 2688
rect 23508 2752 23824 2753
rect 23508 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23824 2752
rect 23508 2687 23824 2688
rect 31213 2752 31529 2753
rect 31213 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31529 2752
rect 31213 2687 31529 2688
rect 4246 2208 4562 2209
rect 4246 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4562 2208
rect 4246 2143 4562 2144
rect 11951 2208 12267 2209
rect 11951 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12267 2208
rect 11951 2143 12267 2144
rect 19656 2208 19972 2209
rect 19656 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19972 2208
rect 19656 2143 19972 2144
rect 27361 2208 27677 2209
rect 27361 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27677 2208
rect 27361 2143 27677 2144
rect 8098 1664 8414 1665
rect 8098 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8414 1664
rect 8098 1599 8414 1600
rect 15803 1664 16119 1665
rect 15803 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16119 1664
rect 15803 1599 16119 1600
rect 23508 1664 23824 1665
rect 23508 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23824 1664
rect 23508 1599 23824 1600
rect 31213 1664 31529 1665
rect 31213 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31529 1664
rect 31213 1599 31529 1600
rect 4246 1120 4562 1121
rect 4246 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4562 1120
rect 4246 1055 4562 1056
rect 11951 1120 12267 1121
rect 11951 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12267 1120
rect 11951 1055 12267 1056
rect 19656 1120 19972 1121
rect 19656 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19972 1120
rect 19656 1055 19972 1056
rect 27361 1120 27677 1121
rect 27361 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27677 1120
rect 27361 1055 27677 1056
rect 8098 576 8414 577
rect 8098 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8414 576
rect 8098 511 8414 512
rect 15803 576 16119 577
rect 15803 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16119 576
rect 15803 511 16119 512
rect 23508 576 23824 577
rect 23508 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23824 576
rect 23508 511 23824 512
rect 31213 576 31529 577
rect 31213 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31529 576
rect 31213 511 31529 512
rect 8293 370 8359 373
rect 15142 370 15148 372
rect 8293 368 15148 370
rect 8293 312 8298 368
rect 8354 312 15148 368
rect 8293 310 15148 312
rect 8293 307 8359 310
rect 15142 308 15148 310
rect 15212 308 15218 372
<< via3 >>
rect 8104 19068 8168 19072
rect 8104 19012 8108 19068
rect 8108 19012 8164 19068
rect 8164 19012 8168 19068
rect 8104 19008 8168 19012
rect 8184 19068 8248 19072
rect 8184 19012 8188 19068
rect 8188 19012 8244 19068
rect 8244 19012 8248 19068
rect 8184 19008 8248 19012
rect 8264 19068 8328 19072
rect 8264 19012 8268 19068
rect 8268 19012 8324 19068
rect 8324 19012 8328 19068
rect 8264 19008 8328 19012
rect 8344 19068 8408 19072
rect 8344 19012 8348 19068
rect 8348 19012 8404 19068
rect 8404 19012 8408 19068
rect 8344 19008 8408 19012
rect 15809 19068 15873 19072
rect 15809 19012 15813 19068
rect 15813 19012 15869 19068
rect 15869 19012 15873 19068
rect 15809 19008 15873 19012
rect 15889 19068 15953 19072
rect 15889 19012 15893 19068
rect 15893 19012 15949 19068
rect 15949 19012 15953 19068
rect 15889 19008 15953 19012
rect 15969 19068 16033 19072
rect 15969 19012 15973 19068
rect 15973 19012 16029 19068
rect 16029 19012 16033 19068
rect 15969 19008 16033 19012
rect 16049 19068 16113 19072
rect 16049 19012 16053 19068
rect 16053 19012 16109 19068
rect 16109 19012 16113 19068
rect 16049 19008 16113 19012
rect 23514 19068 23578 19072
rect 23514 19012 23518 19068
rect 23518 19012 23574 19068
rect 23574 19012 23578 19068
rect 23514 19008 23578 19012
rect 23594 19068 23658 19072
rect 23594 19012 23598 19068
rect 23598 19012 23654 19068
rect 23654 19012 23658 19068
rect 23594 19008 23658 19012
rect 23674 19068 23738 19072
rect 23674 19012 23678 19068
rect 23678 19012 23734 19068
rect 23734 19012 23738 19068
rect 23674 19008 23738 19012
rect 23754 19068 23818 19072
rect 23754 19012 23758 19068
rect 23758 19012 23814 19068
rect 23814 19012 23818 19068
rect 23754 19008 23818 19012
rect 31219 19068 31283 19072
rect 31219 19012 31223 19068
rect 31223 19012 31279 19068
rect 31279 19012 31283 19068
rect 31219 19008 31283 19012
rect 31299 19068 31363 19072
rect 31299 19012 31303 19068
rect 31303 19012 31359 19068
rect 31359 19012 31363 19068
rect 31299 19008 31363 19012
rect 31379 19068 31443 19072
rect 31379 19012 31383 19068
rect 31383 19012 31439 19068
rect 31439 19012 31443 19068
rect 31379 19008 31443 19012
rect 31459 19068 31523 19072
rect 31459 19012 31463 19068
rect 31463 19012 31519 19068
rect 31519 19012 31523 19068
rect 31459 19008 31523 19012
rect 11652 18668 11716 18732
rect 4252 18524 4316 18528
rect 4252 18468 4256 18524
rect 4256 18468 4312 18524
rect 4312 18468 4316 18524
rect 4252 18464 4316 18468
rect 4332 18524 4396 18528
rect 4332 18468 4336 18524
rect 4336 18468 4392 18524
rect 4392 18468 4396 18524
rect 4332 18464 4396 18468
rect 4412 18524 4476 18528
rect 4412 18468 4416 18524
rect 4416 18468 4472 18524
rect 4472 18468 4476 18524
rect 4412 18464 4476 18468
rect 4492 18524 4556 18528
rect 4492 18468 4496 18524
rect 4496 18468 4552 18524
rect 4552 18468 4556 18524
rect 4492 18464 4556 18468
rect 11957 18524 12021 18528
rect 11957 18468 11961 18524
rect 11961 18468 12017 18524
rect 12017 18468 12021 18524
rect 11957 18464 12021 18468
rect 12037 18524 12101 18528
rect 12037 18468 12041 18524
rect 12041 18468 12097 18524
rect 12097 18468 12101 18524
rect 12037 18464 12101 18468
rect 12117 18524 12181 18528
rect 12117 18468 12121 18524
rect 12121 18468 12177 18524
rect 12177 18468 12181 18524
rect 12117 18464 12181 18468
rect 12197 18524 12261 18528
rect 12197 18468 12201 18524
rect 12201 18468 12257 18524
rect 12257 18468 12261 18524
rect 12197 18464 12261 18468
rect 19662 18524 19726 18528
rect 19662 18468 19666 18524
rect 19666 18468 19722 18524
rect 19722 18468 19726 18524
rect 19662 18464 19726 18468
rect 19742 18524 19806 18528
rect 19742 18468 19746 18524
rect 19746 18468 19802 18524
rect 19802 18468 19806 18524
rect 19742 18464 19806 18468
rect 19822 18524 19886 18528
rect 19822 18468 19826 18524
rect 19826 18468 19882 18524
rect 19882 18468 19886 18524
rect 19822 18464 19886 18468
rect 19902 18524 19966 18528
rect 19902 18468 19906 18524
rect 19906 18468 19962 18524
rect 19962 18468 19966 18524
rect 19902 18464 19966 18468
rect 27367 18524 27431 18528
rect 27367 18468 27371 18524
rect 27371 18468 27427 18524
rect 27427 18468 27431 18524
rect 27367 18464 27431 18468
rect 27447 18524 27511 18528
rect 27447 18468 27451 18524
rect 27451 18468 27507 18524
rect 27507 18468 27511 18524
rect 27447 18464 27511 18468
rect 27527 18524 27591 18528
rect 27527 18468 27531 18524
rect 27531 18468 27587 18524
rect 27587 18468 27591 18524
rect 27527 18464 27591 18468
rect 27607 18524 27671 18528
rect 27607 18468 27611 18524
rect 27611 18468 27667 18524
rect 27667 18468 27671 18524
rect 27607 18464 27671 18468
rect 8104 17980 8168 17984
rect 8104 17924 8108 17980
rect 8108 17924 8164 17980
rect 8164 17924 8168 17980
rect 8104 17920 8168 17924
rect 8184 17980 8248 17984
rect 8184 17924 8188 17980
rect 8188 17924 8244 17980
rect 8244 17924 8248 17980
rect 8184 17920 8248 17924
rect 8264 17980 8328 17984
rect 8264 17924 8268 17980
rect 8268 17924 8324 17980
rect 8324 17924 8328 17980
rect 8264 17920 8328 17924
rect 8344 17980 8408 17984
rect 8344 17924 8348 17980
rect 8348 17924 8404 17980
rect 8404 17924 8408 17980
rect 8344 17920 8408 17924
rect 15809 17980 15873 17984
rect 15809 17924 15813 17980
rect 15813 17924 15869 17980
rect 15869 17924 15873 17980
rect 15809 17920 15873 17924
rect 15889 17980 15953 17984
rect 15889 17924 15893 17980
rect 15893 17924 15949 17980
rect 15949 17924 15953 17980
rect 15889 17920 15953 17924
rect 15969 17980 16033 17984
rect 15969 17924 15973 17980
rect 15973 17924 16029 17980
rect 16029 17924 16033 17980
rect 15969 17920 16033 17924
rect 16049 17980 16113 17984
rect 16049 17924 16053 17980
rect 16053 17924 16109 17980
rect 16109 17924 16113 17980
rect 16049 17920 16113 17924
rect 23514 17980 23578 17984
rect 23514 17924 23518 17980
rect 23518 17924 23574 17980
rect 23574 17924 23578 17980
rect 23514 17920 23578 17924
rect 23594 17980 23658 17984
rect 23594 17924 23598 17980
rect 23598 17924 23654 17980
rect 23654 17924 23658 17980
rect 23594 17920 23658 17924
rect 23674 17980 23738 17984
rect 23674 17924 23678 17980
rect 23678 17924 23734 17980
rect 23734 17924 23738 17980
rect 23674 17920 23738 17924
rect 23754 17980 23818 17984
rect 23754 17924 23758 17980
rect 23758 17924 23814 17980
rect 23814 17924 23818 17980
rect 23754 17920 23818 17924
rect 31219 17980 31283 17984
rect 31219 17924 31223 17980
rect 31223 17924 31279 17980
rect 31279 17924 31283 17980
rect 31219 17920 31283 17924
rect 31299 17980 31363 17984
rect 31299 17924 31303 17980
rect 31303 17924 31359 17980
rect 31359 17924 31363 17980
rect 31299 17920 31363 17924
rect 31379 17980 31443 17984
rect 31379 17924 31383 17980
rect 31383 17924 31439 17980
rect 31439 17924 31443 17980
rect 31379 17920 31443 17924
rect 31459 17980 31523 17984
rect 31459 17924 31463 17980
rect 31463 17924 31519 17980
rect 31519 17924 31523 17980
rect 31459 17920 31523 17924
rect 4252 17436 4316 17440
rect 4252 17380 4256 17436
rect 4256 17380 4312 17436
rect 4312 17380 4316 17436
rect 4252 17376 4316 17380
rect 4332 17436 4396 17440
rect 4332 17380 4336 17436
rect 4336 17380 4392 17436
rect 4392 17380 4396 17436
rect 4332 17376 4396 17380
rect 4412 17436 4476 17440
rect 4412 17380 4416 17436
rect 4416 17380 4472 17436
rect 4472 17380 4476 17436
rect 4412 17376 4476 17380
rect 4492 17436 4556 17440
rect 4492 17380 4496 17436
rect 4496 17380 4552 17436
rect 4552 17380 4556 17436
rect 4492 17376 4556 17380
rect 11957 17436 12021 17440
rect 11957 17380 11961 17436
rect 11961 17380 12017 17436
rect 12017 17380 12021 17436
rect 11957 17376 12021 17380
rect 12037 17436 12101 17440
rect 12037 17380 12041 17436
rect 12041 17380 12097 17436
rect 12097 17380 12101 17436
rect 12037 17376 12101 17380
rect 12117 17436 12181 17440
rect 12117 17380 12121 17436
rect 12121 17380 12177 17436
rect 12177 17380 12181 17436
rect 12117 17376 12181 17380
rect 12197 17436 12261 17440
rect 12197 17380 12201 17436
rect 12201 17380 12257 17436
rect 12257 17380 12261 17436
rect 12197 17376 12261 17380
rect 19662 17436 19726 17440
rect 19662 17380 19666 17436
rect 19666 17380 19722 17436
rect 19722 17380 19726 17436
rect 19662 17376 19726 17380
rect 19742 17436 19806 17440
rect 19742 17380 19746 17436
rect 19746 17380 19802 17436
rect 19802 17380 19806 17436
rect 19742 17376 19806 17380
rect 19822 17436 19886 17440
rect 19822 17380 19826 17436
rect 19826 17380 19882 17436
rect 19882 17380 19886 17436
rect 19822 17376 19886 17380
rect 19902 17436 19966 17440
rect 19902 17380 19906 17436
rect 19906 17380 19962 17436
rect 19962 17380 19966 17436
rect 19902 17376 19966 17380
rect 27367 17436 27431 17440
rect 27367 17380 27371 17436
rect 27371 17380 27427 17436
rect 27427 17380 27431 17436
rect 27367 17376 27431 17380
rect 27447 17436 27511 17440
rect 27447 17380 27451 17436
rect 27451 17380 27507 17436
rect 27507 17380 27511 17436
rect 27447 17376 27511 17380
rect 27527 17436 27591 17440
rect 27527 17380 27531 17436
rect 27531 17380 27587 17436
rect 27587 17380 27591 17436
rect 27527 17376 27591 17380
rect 27607 17436 27671 17440
rect 27607 17380 27611 17436
rect 27611 17380 27667 17436
rect 27667 17380 27671 17436
rect 27607 17376 27671 17380
rect 19380 17096 19444 17100
rect 19380 17040 19394 17096
rect 19394 17040 19444 17096
rect 19380 17036 19444 17040
rect 11284 16900 11348 16964
rect 8104 16892 8168 16896
rect 8104 16836 8108 16892
rect 8108 16836 8164 16892
rect 8164 16836 8168 16892
rect 8104 16832 8168 16836
rect 8184 16892 8248 16896
rect 8184 16836 8188 16892
rect 8188 16836 8244 16892
rect 8244 16836 8248 16892
rect 8184 16832 8248 16836
rect 8264 16892 8328 16896
rect 8264 16836 8268 16892
rect 8268 16836 8324 16892
rect 8324 16836 8328 16892
rect 8264 16832 8328 16836
rect 8344 16892 8408 16896
rect 8344 16836 8348 16892
rect 8348 16836 8404 16892
rect 8404 16836 8408 16892
rect 8344 16832 8408 16836
rect 15809 16892 15873 16896
rect 15809 16836 15813 16892
rect 15813 16836 15869 16892
rect 15869 16836 15873 16892
rect 15809 16832 15873 16836
rect 15889 16892 15953 16896
rect 15889 16836 15893 16892
rect 15893 16836 15949 16892
rect 15949 16836 15953 16892
rect 15889 16832 15953 16836
rect 15969 16892 16033 16896
rect 15969 16836 15973 16892
rect 15973 16836 16029 16892
rect 16029 16836 16033 16892
rect 15969 16832 16033 16836
rect 16049 16892 16113 16896
rect 16049 16836 16053 16892
rect 16053 16836 16109 16892
rect 16109 16836 16113 16892
rect 16049 16832 16113 16836
rect 23514 16892 23578 16896
rect 23514 16836 23518 16892
rect 23518 16836 23574 16892
rect 23574 16836 23578 16892
rect 23514 16832 23578 16836
rect 23594 16892 23658 16896
rect 23594 16836 23598 16892
rect 23598 16836 23654 16892
rect 23654 16836 23658 16892
rect 23594 16832 23658 16836
rect 23674 16892 23738 16896
rect 23674 16836 23678 16892
rect 23678 16836 23734 16892
rect 23734 16836 23738 16892
rect 23674 16832 23738 16836
rect 23754 16892 23818 16896
rect 23754 16836 23758 16892
rect 23758 16836 23814 16892
rect 23814 16836 23818 16892
rect 23754 16832 23818 16836
rect 31219 16892 31283 16896
rect 31219 16836 31223 16892
rect 31223 16836 31279 16892
rect 31279 16836 31283 16892
rect 31219 16832 31283 16836
rect 31299 16892 31363 16896
rect 31299 16836 31303 16892
rect 31303 16836 31359 16892
rect 31359 16836 31363 16892
rect 31299 16832 31363 16836
rect 31379 16892 31443 16896
rect 31379 16836 31383 16892
rect 31383 16836 31439 16892
rect 31439 16836 31443 16892
rect 31379 16832 31443 16836
rect 31459 16892 31523 16896
rect 31459 16836 31463 16892
rect 31463 16836 31519 16892
rect 31519 16836 31523 16892
rect 31459 16832 31523 16836
rect 10364 16764 10428 16828
rect 9996 16552 10060 16556
rect 9996 16496 10046 16552
rect 10046 16496 10060 16552
rect 9996 16492 10060 16496
rect 10548 16492 10612 16556
rect 10732 16492 10796 16556
rect 4252 16348 4316 16352
rect 4252 16292 4256 16348
rect 4256 16292 4312 16348
rect 4312 16292 4316 16348
rect 4252 16288 4316 16292
rect 4332 16348 4396 16352
rect 4332 16292 4336 16348
rect 4336 16292 4392 16348
rect 4392 16292 4396 16348
rect 4332 16288 4396 16292
rect 4412 16348 4476 16352
rect 4412 16292 4416 16348
rect 4416 16292 4472 16348
rect 4472 16292 4476 16348
rect 4412 16288 4476 16292
rect 4492 16348 4556 16352
rect 4492 16292 4496 16348
rect 4496 16292 4552 16348
rect 4552 16292 4556 16348
rect 4492 16288 4556 16292
rect 11957 16348 12021 16352
rect 11957 16292 11961 16348
rect 11961 16292 12017 16348
rect 12017 16292 12021 16348
rect 11957 16288 12021 16292
rect 12037 16348 12101 16352
rect 12037 16292 12041 16348
rect 12041 16292 12097 16348
rect 12097 16292 12101 16348
rect 12037 16288 12101 16292
rect 12117 16348 12181 16352
rect 12117 16292 12121 16348
rect 12121 16292 12177 16348
rect 12177 16292 12181 16348
rect 12117 16288 12181 16292
rect 12197 16348 12261 16352
rect 12197 16292 12201 16348
rect 12201 16292 12257 16348
rect 12257 16292 12261 16348
rect 12197 16288 12261 16292
rect 19662 16348 19726 16352
rect 19662 16292 19666 16348
rect 19666 16292 19722 16348
rect 19722 16292 19726 16348
rect 19662 16288 19726 16292
rect 19742 16348 19806 16352
rect 19742 16292 19746 16348
rect 19746 16292 19802 16348
rect 19802 16292 19806 16348
rect 19742 16288 19806 16292
rect 19822 16348 19886 16352
rect 19822 16292 19826 16348
rect 19826 16292 19882 16348
rect 19882 16292 19886 16348
rect 19822 16288 19886 16292
rect 19902 16348 19966 16352
rect 19902 16292 19906 16348
rect 19906 16292 19962 16348
rect 19962 16292 19966 16348
rect 19902 16288 19966 16292
rect 27367 16348 27431 16352
rect 27367 16292 27371 16348
rect 27371 16292 27427 16348
rect 27427 16292 27431 16348
rect 27367 16288 27431 16292
rect 27447 16348 27511 16352
rect 27447 16292 27451 16348
rect 27451 16292 27507 16348
rect 27507 16292 27511 16348
rect 27447 16288 27511 16292
rect 27527 16348 27591 16352
rect 27527 16292 27531 16348
rect 27531 16292 27587 16348
rect 27587 16292 27591 16348
rect 27527 16288 27591 16292
rect 27607 16348 27671 16352
rect 27607 16292 27611 16348
rect 27611 16292 27667 16348
rect 27667 16292 27671 16348
rect 27607 16288 27671 16292
rect 13308 15948 13372 16012
rect 22324 15948 22388 16012
rect 23980 15948 24044 16012
rect 8104 15804 8168 15808
rect 8104 15748 8108 15804
rect 8108 15748 8164 15804
rect 8164 15748 8168 15804
rect 8104 15744 8168 15748
rect 8184 15804 8248 15808
rect 8184 15748 8188 15804
rect 8188 15748 8244 15804
rect 8244 15748 8248 15804
rect 8184 15744 8248 15748
rect 8264 15804 8328 15808
rect 8264 15748 8268 15804
rect 8268 15748 8324 15804
rect 8324 15748 8328 15804
rect 8264 15744 8328 15748
rect 8344 15804 8408 15808
rect 8344 15748 8348 15804
rect 8348 15748 8404 15804
rect 8404 15748 8408 15804
rect 8344 15744 8408 15748
rect 15809 15804 15873 15808
rect 15809 15748 15813 15804
rect 15813 15748 15869 15804
rect 15869 15748 15873 15804
rect 15809 15744 15873 15748
rect 15889 15804 15953 15808
rect 15889 15748 15893 15804
rect 15893 15748 15949 15804
rect 15949 15748 15953 15804
rect 15889 15744 15953 15748
rect 15969 15804 16033 15808
rect 15969 15748 15973 15804
rect 15973 15748 16029 15804
rect 16029 15748 16033 15804
rect 15969 15744 16033 15748
rect 16049 15804 16113 15808
rect 16049 15748 16053 15804
rect 16053 15748 16109 15804
rect 16109 15748 16113 15804
rect 16049 15744 16113 15748
rect 23514 15804 23578 15808
rect 23514 15748 23518 15804
rect 23518 15748 23574 15804
rect 23574 15748 23578 15804
rect 23514 15744 23578 15748
rect 23594 15804 23658 15808
rect 23594 15748 23598 15804
rect 23598 15748 23654 15804
rect 23654 15748 23658 15804
rect 23594 15744 23658 15748
rect 23674 15804 23738 15808
rect 23674 15748 23678 15804
rect 23678 15748 23734 15804
rect 23734 15748 23738 15804
rect 23674 15744 23738 15748
rect 23754 15804 23818 15808
rect 23754 15748 23758 15804
rect 23758 15748 23814 15804
rect 23814 15748 23818 15804
rect 23754 15744 23818 15748
rect 31219 15804 31283 15808
rect 31219 15748 31223 15804
rect 31223 15748 31279 15804
rect 31279 15748 31283 15804
rect 31219 15744 31283 15748
rect 31299 15804 31363 15808
rect 31299 15748 31303 15804
rect 31303 15748 31359 15804
rect 31359 15748 31363 15804
rect 31299 15744 31363 15748
rect 31379 15804 31443 15808
rect 31379 15748 31383 15804
rect 31383 15748 31439 15804
rect 31439 15748 31443 15804
rect 31379 15744 31443 15748
rect 31459 15804 31523 15808
rect 31459 15748 31463 15804
rect 31463 15748 31519 15804
rect 31519 15748 31523 15804
rect 31459 15744 31523 15748
rect 9812 15676 9876 15740
rect 11100 15736 11164 15740
rect 11100 15680 11150 15736
rect 11150 15680 11164 15736
rect 11100 15676 11164 15680
rect 21956 15676 22020 15740
rect 24900 15540 24964 15604
rect 23244 15404 23308 15468
rect 10364 15268 10428 15332
rect 10732 15268 10796 15332
rect 4252 15260 4316 15264
rect 4252 15204 4256 15260
rect 4256 15204 4312 15260
rect 4312 15204 4316 15260
rect 4252 15200 4316 15204
rect 4332 15260 4396 15264
rect 4332 15204 4336 15260
rect 4336 15204 4392 15260
rect 4392 15204 4396 15260
rect 4332 15200 4396 15204
rect 4412 15260 4476 15264
rect 4412 15204 4416 15260
rect 4416 15204 4472 15260
rect 4472 15204 4476 15260
rect 4412 15200 4476 15204
rect 4492 15260 4556 15264
rect 4492 15204 4496 15260
rect 4496 15204 4552 15260
rect 4552 15204 4556 15260
rect 4492 15200 4556 15204
rect 11957 15260 12021 15264
rect 11957 15204 11961 15260
rect 11961 15204 12017 15260
rect 12017 15204 12021 15260
rect 11957 15200 12021 15204
rect 12037 15260 12101 15264
rect 12037 15204 12041 15260
rect 12041 15204 12097 15260
rect 12097 15204 12101 15260
rect 12037 15200 12101 15204
rect 12117 15260 12181 15264
rect 12117 15204 12121 15260
rect 12121 15204 12177 15260
rect 12177 15204 12181 15260
rect 12117 15200 12181 15204
rect 12197 15260 12261 15264
rect 12197 15204 12201 15260
rect 12201 15204 12257 15260
rect 12257 15204 12261 15260
rect 12197 15200 12261 15204
rect 19662 15260 19726 15264
rect 19662 15204 19666 15260
rect 19666 15204 19722 15260
rect 19722 15204 19726 15260
rect 19662 15200 19726 15204
rect 19742 15260 19806 15264
rect 19742 15204 19746 15260
rect 19746 15204 19802 15260
rect 19802 15204 19806 15260
rect 19742 15200 19806 15204
rect 19822 15260 19886 15264
rect 19822 15204 19826 15260
rect 19826 15204 19882 15260
rect 19882 15204 19886 15260
rect 19822 15200 19886 15204
rect 19902 15260 19966 15264
rect 19902 15204 19906 15260
rect 19906 15204 19962 15260
rect 19962 15204 19966 15260
rect 19902 15200 19966 15204
rect 27367 15260 27431 15264
rect 27367 15204 27371 15260
rect 27371 15204 27427 15260
rect 27427 15204 27431 15260
rect 27367 15200 27431 15204
rect 27447 15260 27511 15264
rect 27447 15204 27451 15260
rect 27451 15204 27507 15260
rect 27507 15204 27511 15260
rect 27447 15200 27511 15204
rect 27527 15260 27591 15264
rect 27527 15204 27531 15260
rect 27531 15204 27587 15260
rect 27587 15204 27591 15260
rect 27527 15200 27591 15204
rect 27607 15260 27671 15264
rect 27607 15204 27611 15260
rect 27611 15204 27667 15260
rect 27667 15204 27671 15260
rect 27607 15200 27671 15204
rect 9996 15132 10060 15196
rect 9812 15056 9876 15060
rect 9812 15000 9862 15056
rect 9862 15000 9876 15056
rect 9812 14996 9876 15000
rect 10548 14724 10612 14788
rect 8104 14716 8168 14720
rect 8104 14660 8108 14716
rect 8108 14660 8164 14716
rect 8164 14660 8168 14716
rect 8104 14656 8168 14660
rect 8184 14716 8248 14720
rect 8184 14660 8188 14716
rect 8188 14660 8244 14716
rect 8244 14660 8248 14716
rect 8184 14656 8248 14660
rect 8264 14716 8328 14720
rect 8264 14660 8268 14716
rect 8268 14660 8324 14716
rect 8324 14660 8328 14716
rect 8264 14656 8328 14660
rect 8344 14716 8408 14720
rect 8344 14660 8348 14716
rect 8348 14660 8404 14716
rect 8404 14660 8408 14716
rect 8344 14656 8408 14660
rect 15809 14716 15873 14720
rect 15809 14660 15813 14716
rect 15813 14660 15869 14716
rect 15869 14660 15873 14716
rect 15809 14656 15873 14660
rect 15889 14716 15953 14720
rect 15889 14660 15893 14716
rect 15893 14660 15949 14716
rect 15949 14660 15953 14716
rect 15889 14656 15953 14660
rect 15969 14716 16033 14720
rect 15969 14660 15973 14716
rect 15973 14660 16029 14716
rect 16029 14660 16033 14716
rect 15969 14656 16033 14660
rect 16049 14716 16113 14720
rect 16049 14660 16053 14716
rect 16053 14660 16109 14716
rect 16109 14660 16113 14716
rect 16049 14656 16113 14660
rect 23514 14716 23578 14720
rect 23514 14660 23518 14716
rect 23518 14660 23574 14716
rect 23574 14660 23578 14716
rect 23514 14656 23578 14660
rect 23594 14716 23658 14720
rect 23594 14660 23598 14716
rect 23598 14660 23654 14716
rect 23654 14660 23658 14716
rect 23594 14656 23658 14660
rect 23674 14716 23738 14720
rect 23674 14660 23678 14716
rect 23678 14660 23734 14716
rect 23734 14660 23738 14716
rect 23674 14656 23738 14660
rect 23754 14716 23818 14720
rect 23754 14660 23758 14716
rect 23758 14660 23814 14716
rect 23814 14660 23818 14716
rect 23754 14656 23818 14660
rect 31219 14716 31283 14720
rect 31219 14660 31223 14716
rect 31223 14660 31279 14716
rect 31279 14660 31283 14716
rect 31219 14656 31283 14660
rect 31299 14716 31363 14720
rect 31299 14660 31303 14716
rect 31303 14660 31359 14716
rect 31359 14660 31363 14716
rect 31299 14656 31363 14660
rect 31379 14716 31443 14720
rect 31379 14660 31383 14716
rect 31383 14660 31439 14716
rect 31439 14660 31443 14716
rect 31379 14656 31443 14660
rect 31459 14716 31523 14720
rect 31459 14660 31463 14716
rect 31463 14660 31519 14716
rect 31519 14660 31523 14716
rect 31459 14656 31523 14660
rect 4252 14172 4316 14176
rect 4252 14116 4256 14172
rect 4256 14116 4312 14172
rect 4312 14116 4316 14172
rect 4252 14112 4316 14116
rect 4332 14172 4396 14176
rect 4332 14116 4336 14172
rect 4336 14116 4392 14172
rect 4392 14116 4396 14172
rect 4332 14112 4396 14116
rect 4412 14172 4476 14176
rect 4412 14116 4416 14172
rect 4416 14116 4472 14172
rect 4472 14116 4476 14172
rect 4412 14112 4476 14116
rect 4492 14172 4556 14176
rect 4492 14116 4496 14172
rect 4496 14116 4552 14172
rect 4552 14116 4556 14172
rect 4492 14112 4556 14116
rect 11957 14172 12021 14176
rect 11957 14116 11961 14172
rect 11961 14116 12017 14172
rect 12017 14116 12021 14172
rect 11957 14112 12021 14116
rect 12037 14172 12101 14176
rect 12037 14116 12041 14172
rect 12041 14116 12097 14172
rect 12097 14116 12101 14172
rect 12037 14112 12101 14116
rect 12117 14172 12181 14176
rect 12117 14116 12121 14172
rect 12121 14116 12177 14172
rect 12177 14116 12181 14172
rect 12117 14112 12181 14116
rect 12197 14172 12261 14176
rect 12197 14116 12201 14172
rect 12201 14116 12257 14172
rect 12257 14116 12261 14172
rect 12197 14112 12261 14116
rect 19662 14172 19726 14176
rect 19662 14116 19666 14172
rect 19666 14116 19722 14172
rect 19722 14116 19726 14172
rect 19662 14112 19726 14116
rect 19742 14172 19806 14176
rect 19742 14116 19746 14172
rect 19746 14116 19802 14172
rect 19802 14116 19806 14172
rect 19742 14112 19806 14116
rect 19822 14172 19886 14176
rect 19822 14116 19826 14172
rect 19826 14116 19882 14172
rect 19882 14116 19886 14172
rect 19822 14112 19886 14116
rect 19902 14172 19966 14176
rect 19902 14116 19906 14172
rect 19906 14116 19962 14172
rect 19962 14116 19966 14172
rect 19902 14112 19966 14116
rect 27367 14172 27431 14176
rect 27367 14116 27371 14172
rect 27371 14116 27427 14172
rect 27427 14116 27431 14172
rect 27367 14112 27431 14116
rect 27447 14172 27511 14176
rect 27447 14116 27451 14172
rect 27451 14116 27507 14172
rect 27507 14116 27511 14172
rect 27447 14112 27511 14116
rect 27527 14172 27591 14176
rect 27527 14116 27531 14172
rect 27531 14116 27587 14172
rect 27587 14116 27591 14172
rect 27527 14112 27591 14116
rect 27607 14172 27671 14176
rect 27607 14116 27611 14172
rect 27611 14116 27667 14172
rect 27667 14116 27671 14172
rect 27607 14112 27671 14116
rect 22324 13636 22388 13700
rect 8104 13628 8168 13632
rect 8104 13572 8108 13628
rect 8108 13572 8164 13628
rect 8164 13572 8168 13628
rect 8104 13568 8168 13572
rect 8184 13628 8248 13632
rect 8184 13572 8188 13628
rect 8188 13572 8244 13628
rect 8244 13572 8248 13628
rect 8184 13568 8248 13572
rect 8264 13628 8328 13632
rect 8264 13572 8268 13628
rect 8268 13572 8324 13628
rect 8324 13572 8328 13628
rect 8264 13568 8328 13572
rect 8344 13628 8408 13632
rect 8344 13572 8348 13628
rect 8348 13572 8404 13628
rect 8404 13572 8408 13628
rect 8344 13568 8408 13572
rect 15809 13628 15873 13632
rect 15809 13572 15813 13628
rect 15813 13572 15869 13628
rect 15869 13572 15873 13628
rect 15809 13568 15873 13572
rect 15889 13628 15953 13632
rect 15889 13572 15893 13628
rect 15893 13572 15949 13628
rect 15949 13572 15953 13628
rect 15889 13568 15953 13572
rect 15969 13628 16033 13632
rect 15969 13572 15973 13628
rect 15973 13572 16029 13628
rect 16029 13572 16033 13628
rect 15969 13568 16033 13572
rect 16049 13628 16113 13632
rect 16049 13572 16053 13628
rect 16053 13572 16109 13628
rect 16109 13572 16113 13628
rect 16049 13568 16113 13572
rect 23514 13628 23578 13632
rect 23514 13572 23518 13628
rect 23518 13572 23574 13628
rect 23574 13572 23578 13628
rect 23514 13568 23578 13572
rect 23594 13628 23658 13632
rect 23594 13572 23598 13628
rect 23598 13572 23654 13628
rect 23654 13572 23658 13628
rect 23594 13568 23658 13572
rect 23674 13628 23738 13632
rect 23674 13572 23678 13628
rect 23678 13572 23734 13628
rect 23734 13572 23738 13628
rect 23674 13568 23738 13572
rect 23754 13628 23818 13632
rect 23754 13572 23758 13628
rect 23758 13572 23814 13628
rect 23814 13572 23818 13628
rect 23754 13568 23818 13572
rect 31219 13628 31283 13632
rect 31219 13572 31223 13628
rect 31223 13572 31279 13628
rect 31279 13572 31283 13628
rect 31219 13568 31283 13572
rect 31299 13628 31363 13632
rect 31299 13572 31303 13628
rect 31303 13572 31359 13628
rect 31359 13572 31363 13628
rect 31299 13568 31363 13572
rect 31379 13628 31443 13632
rect 31379 13572 31383 13628
rect 31383 13572 31439 13628
rect 31439 13572 31443 13628
rect 31379 13568 31443 13572
rect 31459 13628 31523 13632
rect 31459 13572 31463 13628
rect 31463 13572 31519 13628
rect 31519 13572 31523 13628
rect 31459 13568 31523 13572
rect 11100 13364 11164 13428
rect 21956 13364 22020 13428
rect 24900 13152 24964 13156
rect 24900 13096 24914 13152
rect 24914 13096 24964 13152
rect 24900 13092 24964 13096
rect 4252 13084 4316 13088
rect 4252 13028 4256 13084
rect 4256 13028 4312 13084
rect 4312 13028 4316 13084
rect 4252 13024 4316 13028
rect 4332 13084 4396 13088
rect 4332 13028 4336 13084
rect 4336 13028 4392 13084
rect 4392 13028 4396 13084
rect 4332 13024 4396 13028
rect 4412 13084 4476 13088
rect 4412 13028 4416 13084
rect 4416 13028 4472 13084
rect 4472 13028 4476 13084
rect 4412 13024 4476 13028
rect 4492 13084 4556 13088
rect 4492 13028 4496 13084
rect 4496 13028 4552 13084
rect 4552 13028 4556 13084
rect 4492 13024 4556 13028
rect 11957 13084 12021 13088
rect 11957 13028 11961 13084
rect 11961 13028 12017 13084
rect 12017 13028 12021 13084
rect 11957 13024 12021 13028
rect 12037 13084 12101 13088
rect 12037 13028 12041 13084
rect 12041 13028 12097 13084
rect 12097 13028 12101 13084
rect 12037 13024 12101 13028
rect 12117 13084 12181 13088
rect 12117 13028 12121 13084
rect 12121 13028 12177 13084
rect 12177 13028 12181 13084
rect 12117 13024 12181 13028
rect 12197 13084 12261 13088
rect 12197 13028 12201 13084
rect 12201 13028 12257 13084
rect 12257 13028 12261 13084
rect 12197 13024 12261 13028
rect 19662 13084 19726 13088
rect 19662 13028 19666 13084
rect 19666 13028 19722 13084
rect 19722 13028 19726 13084
rect 19662 13024 19726 13028
rect 19742 13084 19806 13088
rect 19742 13028 19746 13084
rect 19746 13028 19802 13084
rect 19802 13028 19806 13084
rect 19742 13024 19806 13028
rect 19822 13084 19886 13088
rect 19822 13028 19826 13084
rect 19826 13028 19882 13084
rect 19882 13028 19886 13084
rect 19822 13024 19886 13028
rect 19902 13084 19966 13088
rect 19902 13028 19906 13084
rect 19906 13028 19962 13084
rect 19962 13028 19966 13084
rect 19902 13024 19966 13028
rect 27367 13084 27431 13088
rect 27367 13028 27371 13084
rect 27371 13028 27427 13084
rect 27427 13028 27431 13084
rect 27367 13024 27431 13028
rect 27447 13084 27511 13088
rect 27447 13028 27451 13084
rect 27451 13028 27507 13084
rect 27507 13028 27511 13084
rect 27447 13024 27511 13028
rect 27527 13084 27591 13088
rect 27527 13028 27531 13084
rect 27531 13028 27587 13084
rect 27587 13028 27591 13084
rect 27527 13024 27591 13028
rect 27607 13084 27671 13088
rect 27607 13028 27611 13084
rect 27611 13028 27667 13084
rect 27667 13028 27671 13084
rect 27607 13024 27671 13028
rect 11284 13016 11348 13020
rect 11284 12960 11334 13016
rect 11334 12960 11348 13016
rect 11284 12956 11348 12960
rect 11652 13016 11716 13020
rect 11652 12960 11702 13016
rect 11702 12960 11716 13016
rect 11652 12956 11716 12960
rect 23244 12820 23308 12884
rect 8104 12540 8168 12544
rect 8104 12484 8108 12540
rect 8108 12484 8164 12540
rect 8164 12484 8168 12540
rect 8104 12480 8168 12484
rect 8184 12540 8248 12544
rect 8184 12484 8188 12540
rect 8188 12484 8244 12540
rect 8244 12484 8248 12540
rect 8184 12480 8248 12484
rect 8264 12540 8328 12544
rect 8264 12484 8268 12540
rect 8268 12484 8324 12540
rect 8324 12484 8328 12540
rect 8264 12480 8328 12484
rect 8344 12540 8408 12544
rect 8344 12484 8348 12540
rect 8348 12484 8404 12540
rect 8404 12484 8408 12540
rect 8344 12480 8408 12484
rect 15809 12540 15873 12544
rect 15809 12484 15813 12540
rect 15813 12484 15869 12540
rect 15869 12484 15873 12540
rect 15809 12480 15873 12484
rect 15889 12540 15953 12544
rect 15889 12484 15893 12540
rect 15893 12484 15949 12540
rect 15949 12484 15953 12540
rect 15889 12480 15953 12484
rect 15969 12540 16033 12544
rect 15969 12484 15973 12540
rect 15973 12484 16029 12540
rect 16029 12484 16033 12540
rect 15969 12480 16033 12484
rect 16049 12540 16113 12544
rect 16049 12484 16053 12540
rect 16053 12484 16109 12540
rect 16109 12484 16113 12540
rect 16049 12480 16113 12484
rect 23514 12540 23578 12544
rect 23514 12484 23518 12540
rect 23518 12484 23574 12540
rect 23574 12484 23578 12540
rect 23514 12480 23578 12484
rect 23594 12540 23658 12544
rect 23594 12484 23598 12540
rect 23598 12484 23654 12540
rect 23654 12484 23658 12540
rect 23594 12480 23658 12484
rect 23674 12540 23738 12544
rect 23674 12484 23678 12540
rect 23678 12484 23734 12540
rect 23734 12484 23738 12540
rect 23674 12480 23738 12484
rect 23754 12540 23818 12544
rect 23754 12484 23758 12540
rect 23758 12484 23814 12540
rect 23814 12484 23818 12540
rect 23754 12480 23818 12484
rect 31219 12540 31283 12544
rect 31219 12484 31223 12540
rect 31223 12484 31279 12540
rect 31279 12484 31283 12540
rect 31219 12480 31283 12484
rect 31299 12540 31363 12544
rect 31299 12484 31303 12540
rect 31303 12484 31359 12540
rect 31359 12484 31363 12540
rect 31299 12480 31363 12484
rect 31379 12540 31443 12544
rect 31379 12484 31383 12540
rect 31383 12484 31439 12540
rect 31439 12484 31443 12540
rect 31379 12480 31443 12484
rect 31459 12540 31523 12544
rect 31459 12484 31463 12540
rect 31463 12484 31519 12540
rect 31519 12484 31523 12540
rect 31459 12480 31523 12484
rect 23980 12276 24044 12340
rect 4252 11996 4316 12000
rect 4252 11940 4256 11996
rect 4256 11940 4312 11996
rect 4312 11940 4316 11996
rect 4252 11936 4316 11940
rect 4332 11996 4396 12000
rect 4332 11940 4336 11996
rect 4336 11940 4392 11996
rect 4392 11940 4396 11996
rect 4332 11936 4396 11940
rect 4412 11996 4476 12000
rect 4412 11940 4416 11996
rect 4416 11940 4472 11996
rect 4472 11940 4476 11996
rect 4412 11936 4476 11940
rect 4492 11996 4556 12000
rect 4492 11940 4496 11996
rect 4496 11940 4552 11996
rect 4552 11940 4556 11996
rect 4492 11936 4556 11940
rect 11957 11996 12021 12000
rect 11957 11940 11961 11996
rect 11961 11940 12017 11996
rect 12017 11940 12021 11996
rect 11957 11936 12021 11940
rect 12037 11996 12101 12000
rect 12037 11940 12041 11996
rect 12041 11940 12097 11996
rect 12097 11940 12101 11996
rect 12037 11936 12101 11940
rect 12117 11996 12181 12000
rect 12117 11940 12121 11996
rect 12121 11940 12177 11996
rect 12177 11940 12181 11996
rect 12117 11936 12181 11940
rect 12197 11996 12261 12000
rect 12197 11940 12201 11996
rect 12201 11940 12257 11996
rect 12257 11940 12261 11996
rect 12197 11936 12261 11940
rect 19662 11996 19726 12000
rect 19662 11940 19666 11996
rect 19666 11940 19722 11996
rect 19722 11940 19726 11996
rect 19662 11936 19726 11940
rect 19742 11996 19806 12000
rect 19742 11940 19746 11996
rect 19746 11940 19802 11996
rect 19802 11940 19806 11996
rect 19742 11936 19806 11940
rect 19822 11996 19886 12000
rect 19822 11940 19826 11996
rect 19826 11940 19882 11996
rect 19882 11940 19886 11996
rect 19822 11936 19886 11940
rect 19902 11996 19966 12000
rect 19902 11940 19906 11996
rect 19906 11940 19962 11996
rect 19962 11940 19966 11996
rect 19902 11936 19966 11940
rect 27367 11996 27431 12000
rect 27367 11940 27371 11996
rect 27371 11940 27427 11996
rect 27427 11940 27431 11996
rect 27367 11936 27431 11940
rect 27447 11996 27511 12000
rect 27447 11940 27451 11996
rect 27451 11940 27507 11996
rect 27507 11940 27511 11996
rect 27447 11936 27511 11940
rect 27527 11996 27591 12000
rect 27527 11940 27531 11996
rect 27531 11940 27587 11996
rect 27587 11940 27591 11996
rect 27527 11936 27591 11940
rect 27607 11996 27671 12000
rect 27607 11940 27611 11996
rect 27611 11940 27667 11996
rect 27667 11940 27671 11996
rect 27607 11936 27671 11940
rect 19380 11792 19444 11796
rect 19380 11736 19394 11792
rect 19394 11736 19444 11792
rect 19380 11732 19444 11736
rect 8104 11452 8168 11456
rect 8104 11396 8108 11452
rect 8108 11396 8164 11452
rect 8164 11396 8168 11452
rect 8104 11392 8168 11396
rect 8184 11452 8248 11456
rect 8184 11396 8188 11452
rect 8188 11396 8244 11452
rect 8244 11396 8248 11452
rect 8184 11392 8248 11396
rect 8264 11452 8328 11456
rect 8264 11396 8268 11452
rect 8268 11396 8324 11452
rect 8324 11396 8328 11452
rect 8264 11392 8328 11396
rect 8344 11452 8408 11456
rect 8344 11396 8348 11452
rect 8348 11396 8404 11452
rect 8404 11396 8408 11452
rect 8344 11392 8408 11396
rect 15809 11452 15873 11456
rect 15809 11396 15813 11452
rect 15813 11396 15869 11452
rect 15869 11396 15873 11452
rect 15809 11392 15873 11396
rect 15889 11452 15953 11456
rect 15889 11396 15893 11452
rect 15893 11396 15949 11452
rect 15949 11396 15953 11452
rect 15889 11392 15953 11396
rect 15969 11452 16033 11456
rect 15969 11396 15973 11452
rect 15973 11396 16029 11452
rect 16029 11396 16033 11452
rect 15969 11392 16033 11396
rect 16049 11452 16113 11456
rect 16049 11396 16053 11452
rect 16053 11396 16109 11452
rect 16109 11396 16113 11452
rect 16049 11392 16113 11396
rect 23514 11452 23578 11456
rect 23514 11396 23518 11452
rect 23518 11396 23574 11452
rect 23574 11396 23578 11452
rect 23514 11392 23578 11396
rect 23594 11452 23658 11456
rect 23594 11396 23598 11452
rect 23598 11396 23654 11452
rect 23654 11396 23658 11452
rect 23594 11392 23658 11396
rect 23674 11452 23738 11456
rect 23674 11396 23678 11452
rect 23678 11396 23734 11452
rect 23734 11396 23738 11452
rect 23674 11392 23738 11396
rect 23754 11452 23818 11456
rect 23754 11396 23758 11452
rect 23758 11396 23814 11452
rect 23814 11396 23818 11452
rect 23754 11392 23818 11396
rect 31219 11452 31283 11456
rect 31219 11396 31223 11452
rect 31223 11396 31279 11452
rect 31279 11396 31283 11452
rect 31219 11392 31283 11396
rect 31299 11452 31363 11456
rect 31299 11396 31303 11452
rect 31303 11396 31359 11452
rect 31359 11396 31363 11452
rect 31299 11392 31363 11396
rect 31379 11452 31443 11456
rect 31379 11396 31383 11452
rect 31383 11396 31439 11452
rect 31439 11396 31443 11452
rect 31379 11392 31443 11396
rect 31459 11452 31523 11456
rect 31459 11396 31463 11452
rect 31463 11396 31519 11452
rect 31519 11396 31523 11452
rect 31459 11392 31523 11396
rect 13308 10976 13372 10980
rect 13308 10920 13322 10976
rect 13322 10920 13372 10976
rect 13308 10916 13372 10920
rect 4252 10908 4316 10912
rect 4252 10852 4256 10908
rect 4256 10852 4312 10908
rect 4312 10852 4316 10908
rect 4252 10848 4316 10852
rect 4332 10908 4396 10912
rect 4332 10852 4336 10908
rect 4336 10852 4392 10908
rect 4392 10852 4396 10908
rect 4332 10848 4396 10852
rect 4412 10908 4476 10912
rect 4412 10852 4416 10908
rect 4416 10852 4472 10908
rect 4472 10852 4476 10908
rect 4412 10848 4476 10852
rect 4492 10908 4556 10912
rect 4492 10852 4496 10908
rect 4496 10852 4552 10908
rect 4552 10852 4556 10908
rect 4492 10848 4556 10852
rect 11957 10908 12021 10912
rect 11957 10852 11961 10908
rect 11961 10852 12017 10908
rect 12017 10852 12021 10908
rect 11957 10848 12021 10852
rect 12037 10908 12101 10912
rect 12037 10852 12041 10908
rect 12041 10852 12097 10908
rect 12097 10852 12101 10908
rect 12037 10848 12101 10852
rect 12117 10908 12181 10912
rect 12117 10852 12121 10908
rect 12121 10852 12177 10908
rect 12177 10852 12181 10908
rect 12117 10848 12181 10852
rect 12197 10908 12261 10912
rect 12197 10852 12201 10908
rect 12201 10852 12257 10908
rect 12257 10852 12261 10908
rect 12197 10848 12261 10852
rect 19662 10908 19726 10912
rect 19662 10852 19666 10908
rect 19666 10852 19722 10908
rect 19722 10852 19726 10908
rect 19662 10848 19726 10852
rect 19742 10908 19806 10912
rect 19742 10852 19746 10908
rect 19746 10852 19802 10908
rect 19802 10852 19806 10908
rect 19742 10848 19806 10852
rect 19822 10908 19886 10912
rect 19822 10852 19826 10908
rect 19826 10852 19882 10908
rect 19882 10852 19886 10908
rect 19822 10848 19886 10852
rect 19902 10908 19966 10912
rect 19902 10852 19906 10908
rect 19906 10852 19962 10908
rect 19962 10852 19966 10908
rect 19902 10848 19966 10852
rect 27367 10908 27431 10912
rect 27367 10852 27371 10908
rect 27371 10852 27427 10908
rect 27427 10852 27431 10908
rect 27367 10848 27431 10852
rect 27447 10908 27511 10912
rect 27447 10852 27451 10908
rect 27451 10852 27507 10908
rect 27507 10852 27511 10908
rect 27447 10848 27511 10852
rect 27527 10908 27591 10912
rect 27527 10852 27531 10908
rect 27531 10852 27587 10908
rect 27587 10852 27591 10908
rect 27527 10848 27591 10852
rect 27607 10908 27671 10912
rect 27607 10852 27611 10908
rect 27611 10852 27667 10908
rect 27667 10852 27671 10908
rect 27607 10848 27671 10852
rect 8104 10364 8168 10368
rect 8104 10308 8108 10364
rect 8108 10308 8164 10364
rect 8164 10308 8168 10364
rect 8104 10304 8168 10308
rect 8184 10364 8248 10368
rect 8184 10308 8188 10364
rect 8188 10308 8244 10364
rect 8244 10308 8248 10364
rect 8184 10304 8248 10308
rect 8264 10364 8328 10368
rect 8264 10308 8268 10364
rect 8268 10308 8324 10364
rect 8324 10308 8328 10364
rect 8264 10304 8328 10308
rect 8344 10364 8408 10368
rect 8344 10308 8348 10364
rect 8348 10308 8404 10364
rect 8404 10308 8408 10364
rect 8344 10304 8408 10308
rect 15809 10364 15873 10368
rect 15809 10308 15813 10364
rect 15813 10308 15869 10364
rect 15869 10308 15873 10364
rect 15809 10304 15873 10308
rect 15889 10364 15953 10368
rect 15889 10308 15893 10364
rect 15893 10308 15949 10364
rect 15949 10308 15953 10364
rect 15889 10304 15953 10308
rect 15969 10364 16033 10368
rect 15969 10308 15973 10364
rect 15973 10308 16029 10364
rect 16029 10308 16033 10364
rect 15969 10304 16033 10308
rect 16049 10364 16113 10368
rect 16049 10308 16053 10364
rect 16053 10308 16109 10364
rect 16109 10308 16113 10364
rect 16049 10304 16113 10308
rect 23514 10364 23578 10368
rect 23514 10308 23518 10364
rect 23518 10308 23574 10364
rect 23574 10308 23578 10364
rect 23514 10304 23578 10308
rect 23594 10364 23658 10368
rect 23594 10308 23598 10364
rect 23598 10308 23654 10364
rect 23654 10308 23658 10364
rect 23594 10304 23658 10308
rect 23674 10364 23738 10368
rect 23674 10308 23678 10364
rect 23678 10308 23734 10364
rect 23734 10308 23738 10364
rect 23674 10304 23738 10308
rect 23754 10364 23818 10368
rect 23754 10308 23758 10364
rect 23758 10308 23814 10364
rect 23814 10308 23818 10364
rect 23754 10304 23818 10308
rect 31219 10364 31283 10368
rect 31219 10308 31223 10364
rect 31223 10308 31279 10364
rect 31279 10308 31283 10364
rect 31219 10304 31283 10308
rect 31299 10364 31363 10368
rect 31299 10308 31303 10364
rect 31303 10308 31359 10364
rect 31359 10308 31363 10364
rect 31299 10304 31363 10308
rect 31379 10364 31443 10368
rect 31379 10308 31383 10364
rect 31383 10308 31439 10364
rect 31439 10308 31443 10364
rect 31379 10304 31443 10308
rect 31459 10364 31523 10368
rect 31459 10308 31463 10364
rect 31463 10308 31519 10364
rect 31519 10308 31523 10364
rect 31459 10304 31523 10308
rect 4252 9820 4316 9824
rect 4252 9764 4256 9820
rect 4256 9764 4312 9820
rect 4312 9764 4316 9820
rect 4252 9760 4316 9764
rect 4332 9820 4396 9824
rect 4332 9764 4336 9820
rect 4336 9764 4392 9820
rect 4392 9764 4396 9820
rect 4332 9760 4396 9764
rect 4412 9820 4476 9824
rect 4412 9764 4416 9820
rect 4416 9764 4472 9820
rect 4472 9764 4476 9820
rect 4412 9760 4476 9764
rect 4492 9820 4556 9824
rect 4492 9764 4496 9820
rect 4496 9764 4552 9820
rect 4552 9764 4556 9820
rect 4492 9760 4556 9764
rect 11957 9820 12021 9824
rect 11957 9764 11961 9820
rect 11961 9764 12017 9820
rect 12017 9764 12021 9820
rect 11957 9760 12021 9764
rect 12037 9820 12101 9824
rect 12037 9764 12041 9820
rect 12041 9764 12097 9820
rect 12097 9764 12101 9820
rect 12037 9760 12101 9764
rect 12117 9820 12181 9824
rect 12117 9764 12121 9820
rect 12121 9764 12177 9820
rect 12177 9764 12181 9820
rect 12117 9760 12181 9764
rect 12197 9820 12261 9824
rect 12197 9764 12201 9820
rect 12201 9764 12257 9820
rect 12257 9764 12261 9820
rect 12197 9760 12261 9764
rect 19662 9820 19726 9824
rect 19662 9764 19666 9820
rect 19666 9764 19722 9820
rect 19722 9764 19726 9820
rect 19662 9760 19726 9764
rect 19742 9820 19806 9824
rect 19742 9764 19746 9820
rect 19746 9764 19802 9820
rect 19802 9764 19806 9820
rect 19742 9760 19806 9764
rect 19822 9820 19886 9824
rect 19822 9764 19826 9820
rect 19826 9764 19882 9820
rect 19882 9764 19886 9820
rect 19822 9760 19886 9764
rect 19902 9820 19966 9824
rect 19902 9764 19906 9820
rect 19906 9764 19962 9820
rect 19962 9764 19966 9820
rect 19902 9760 19966 9764
rect 27367 9820 27431 9824
rect 27367 9764 27371 9820
rect 27371 9764 27427 9820
rect 27427 9764 27431 9820
rect 27367 9760 27431 9764
rect 27447 9820 27511 9824
rect 27447 9764 27451 9820
rect 27451 9764 27507 9820
rect 27507 9764 27511 9820
rect 27447 9760 27511 9764
rect 27527 9820 27591 9824
rect 27527 9764 27531 9820
rect 27531 9764 27587 9820
rect 27587 9764 27591 9820
rect 27527 9760 27591 9764
rect 27607 9820 27671 9824
rect 27607 9764 27611 9820
rect 27611 9764 27667 9820
rect 27667 9764 27671 9820
rect 27607 9760 27671 9764
rect 8104 9276 8168 9280
rect 8104 9220 8108 9276
rect 8108 9220 8164 9276
rect 8164 9220 8168 9276
rect 8104 9216 8168 9220
rect 8184 9276 8248 9280
rect 8184 9220 8188 9276
rect 8188 9220 8244 9276
rect 8244 9220 8248 9276
rect 8184 9216 8248 9220
rect 8264 9276 8328 9280
rect 8264 9220 8268 9276
rect 8268 9220 8324 9276
rect 8324 9220 8328 9276
rect 8264 9216 8328 9220
rect 8344 9276 8408 9280
rect 8344 9220 8348 9276
rect 8348 9220 8404 9276
rect 8404 9220 8408 9276
rect 8344 9216 8408 9220
rect 15809 9276 15873 9280
rect 15809 9220 15813 9276
rect 15813 9220 15869 9276
rect 15869 9220 15873 9276
rect 15809 9216 15873 9220
rect 15889 9276 15953 9280
rect 15889 9220 15893 9276
rect 15893 9220 15949 9276
rect 15949 9220 15953 9276
rect 15889 9216 15953 9220
rect 15969 9276 16033 9280
rect 15969 9220 15973 9276
rect 15973 9220 16029 9276
rect 16029 9220 16033 9276
rect 15969 9216 16033 9220
rect 16049 9276 16113 9280
rect 16049 9220 16053 9276
rect 16053 9220 16109 9276
rect 16109 9220 16113 9276
rect 16049 9216 16113 9220
rect 23514 9276 23578 9280
rect 23514 9220 23518 9276
rect 23518 9220 23574 9276
rect 23574 9220 23578 9276
rect 23514 9216 23578 9220
rect 23594 9276 23658 9280
rect 23594 9220 23598 9276
rect 23598 9220 23654 9276
rect 23654 9220 23658 9276
rect 23594 9216 23658 9220
rect 23674 9276 23738 9280
rect 23674 9220 23678 9276
rect 23678 9220 23734 9276
rect 23734 9220 23738 9276
rect 23674 9216 23738 9220
rect 23754 9276 23818 9280
rect 23754 9220 23758 9276
rect 23758 9220 23814 9276
rect 23814 9220 23818 9276
rect 23754 9216 23818 9220
rect 31219 9276 31283 9280
rect 31219 9220 31223 9276
rect 31223 9220 31279 9276
rect 31279 9220 31283 9276
rect 31219 9216 31283 9220
rect 31299 9276 31363 9280
rect 31299 9220 31303 9276
rect 31303 9220 31359 9276
rect 31359 9220 31363 9276
rect 31299 9216 31363 9220
rect 31379 9276 31443 9280
rect 31379 9220 31383 9276
rect 31383 9220 31439 9276
rect 31439 9220 31443 9276
rect 31379 9216 31443 9220
rect 31459 9276 31523 9280
rect 31459 9220 31463 9276
rect 31463 9220 31519 9276
rect 31519 9220 31523 9276
rect 31459 9216 31523 9220
rect 4252 8732 4316 8736
rect 4252 8676 4256 8732
rect 4256 8676 4312 8732
rect 4312 8676 4316 8732
rect 4252 8672 4316 8676
rect 4332 8732 4396 8736
rect 4332 8676 4336 8732
rect 4336 8676 4392 8732
rect 4392 8676 4396 8732
rect 4332 8672 4396 8676
rect 4412 8732 4476 8736
rect 4412 8676 4416 8732
rect 4416 8676 4472 8732
rect 4472 8676 4476 8732
rect 4412 8672 4476 8676
rect 4492 8732 4556 8736
rect 4492 8676 4496 8732
rect 4496 8676 4552 8732
rect 4552 8676 4556 8732
rect 4492 8672 4556 8676
rect 11957 8732 12021 8736
rect 11957 8676 11961 8732
rect 11961 8676 12017 8732
rect 12017 8676 12021 8732
rect 11957 8672 12021 8676
rect 12037 8732 12101 8736
rect 12037 8676 12041 8732
rect 12041 8676 12097 8732
rect 12097 8676 12101 8732
rect 12037 8672 12101 8676
rect 12117 8732 12181 8736
rect 12117 8676 12121 8732
rect 12121 8676 12177 8732
rect 12177 8676 12181 8732
rect 12117 8672 12181 8676
rect 12197 8732 12261 8736
rect 12197 8676 12201 8732
rect 12201 8676 12257 8732
rect 12257 8676 12261 8732
rect 12197 8672 12261 8676
rect 19662 8732 19726 8736
rect 19662 8676 19666 8732
rect 19666 8676 19722 8732
rect 19722 8676 19726 8732
rect 19662 8672 19726 8676
rect 19742 8732 19806 8736
rect 19742 8676 19746 8732
rect 19746 8676 19802 8732
rect 19802 8676 19806 8732
rect 19742 8672 19806 8676
rect 19822 8732 19886 8736
rect 19822 8676 19826 8732
rect 19826 8676 19882 8732
rect 19882 8676 19886 8732
rect 19822 8672 19886 8676
rect 19902 8732 19966 8736
rect 19902 8676 19906 8732
rect 19906 8676 19962 8732
rect 19962 8676 19966 8732
rect 19902 8672 19966 8676
rect 27367 8732 27431 8736
rect 27367 8676 27371 8732
rect 27371 8676 27427 8732
rect 27427 8676 27431 8732
rect 27367 8672 27431 8676
rect 27447 8732 27511 8736
rect 27447 8676 27451 8732
rect 27451 8676 27507 8732
rect 27507 8676 27511 8732
rect 27447 8672 27511 8676
rect 27527 8732 27591 8736
rect 27527 8676 27531 8732
rect 27531 8676 27587 8732
rect 27587 8676 27591 8732
rect 27527 8672 27591 8676
rect 27607 8732 27671 8736
rect 27607 8676 27611 8732
rect 27611 8676 27667 8732
rect 27667 8676 27671 8732
rect 27607 8672 27671 8676
rect 15148 8392 15212 8396
rect 15148 8336 15198 8392
rect 15198 8336 15212 8392
rect 15148 8332 15212 8336
rect 20668 8332 20732 8396
rect 8104 8188 8168 8192
rect 8104 8132 8108 8188
rect 8108 8132 8164 8188
rect 8164 8132 8168 8188
rect 8104 8128 8168 8132
rect 8184 8188 8248 8192
rect 8184 8132 8188 8188
rect 8188 8132 8244 8188
rect 8244 8132 8248 8188
rect 8184 8128 8248 8132
rect 8264 8188 8328 8192
rect 8264 8132 8268 8188
rect 8268 8132 8324 8188
rect 8324 8132 8328 8188
rect 8264 8128 8328 8132
rect 8344 8188 8408 8192
rect 8344 8132 8348 8188
rect 8348 8132 8404 8188
rect 8404 8132 8408 8188
rect 8344 8128 8408 8132
rect 15809 8188 15873 8192
rect 15809 8132 15813 8188
rect 15813 8132 15869 8188
rect 15869 8132 15873 8188
rect 15809 8128 15873 8132
rect 15889 8188 15953 8192
rect 15889 8132 15893 8188
rect 15893 8132 15949 8188
rect 15949 8132 15953 8188
rect 15889 8128 15953 8132
rect 15969 8188 16033 8192
rect 15969 8132 15973 8188
rect 15973 8132 16029 8188
rect 16029 8132 16033 8188
rect 15969 8128 16033 8132
rect 16049 8188 16113 8192
rect 16049 8132 16053 8188
rect 16053 8132 16109 8188
rect 16109 8132 16113 8188
rect 16049 8128 16113 8132
rect 23514 8188 23578 8192
rect 23514 8132 23518 8188
rect 23518 8132 23574 8188
rect 23574 8132 23578 8188
rect 23514 8128 23578 8132
rect 23594 8188 23658 8192
rect 23594 8132 23598 8188
rect 23598 8132 23654 8188
rect 23654 8132 23658 8188
rect 23594 8128 23658 8132
rect 23674 8188 23738 8192
rect 23674 8132 23678 8188
rect 23678 8132 23734 8188
rect 23734 8132 23738 8188
rect 23674 8128 23738 8132
rect 23754 8188 23818 8192
rect 23754 8132 23758 8188
rect 23758 8132 23814 8188
rect 23814 8132 23818 8188
rect 23754 8128 23818 8132
rect 4252 7644 4316 7648
rect 4252 7588 4256 7644
rect 4256 7588 4312 7644
rect 4312 7588 4316 7644
rect 4252 7584 4316 7588
rect 4332 7644 4396 7648
rect 4332 7588 4336 7644
rect 4336 7588 4392 7644
rect 4392 7588 4396 7644
rect 4332 7584 4396 7588
rect 4412 7644 4476 7648
rect 4412 7588 4416 7644
rect 4416 7588 4472 7644
rect 4472 7588 4476 7644
rect 4412 7584 4476 7588
rect 4492 7644 4556 7648
rect 4492 7588 4496 7644
rect 4496 7588 4552 7644
rect 4552 7588 4556 7644
rect 4492 7584 4556 7588
rect 11957 7644 12021 7648
rect 11957 7588 11961 7644
rect 11961 7588 12017 7644
rect 12017 7588 12021 7644
rect 11957 7584 12021 7588
rect 12037 7644 12101 7648
rect 12037 7588 12041 7644
rect 12041 7588 12097 7644
rect 12097 7588 12101 7644
rect 12037 7584 12101 7588
rect 12117 7644 12181 7648
rect 12117 7588 12121 7644
rect 12121 7588 12177 7644
rect 12177 7588 12181 7644
rect 12117 7584 12181 7588
rect 12197 7644 12261 7648
rect 12197 7588 12201 7644
rect 12201 7588 12257 7644
rect 12257 7588 12261 7644
rect 12197 7584 12261 7588
rect 19662 7644 19726 7648
rect 19662 7588 19666 7644
rect 19666 7588 19722 7644
rect 19722 7588 19726 7644
rect 19662 7584 19726 7588
rect 19742 7644 19806 7648
rect 19742 7588 19746 7644
rect 19746 7588 19802 7644
rect 19802 7588 19806 7644
rect 19742 7584 19806 7588
rect 19822 7644 19886 7648
rect 19822 7588 19826 7644
rect 19826 7588 19882 7644
rect 19882 7588 19886 7644
rect 19822 7584 19886 7588
rect 19902 7644 19966 7648
rect 19902 7588 19906 7644
rect 19906 7588 19962 7644
rect 19962 7588 19966 7644
rect 19902 7584 19966 7588
rect 27367 7644 27431 7648
rect 27367 7588 27371 7644
rect 27371 7588 27427 7644
rect 27427 7588 27431 7644
rect 27367 7584 27431 7588
rect 27447 7644 27511 7648
rect 27447 7588 27451 7644
rect 27451 7588 27507 7644
rect 27507 7588 27511 7644
rect 27447 7584 27511 7588
rect 27527 7644 27591 7648
rect 27527 7588 27531 7644
rect 27531 7588 27587 7644
rect 27587 7588 27591 7644
rect 27527 7584 27591 7588
rect 27607 7644 27671 7648
rect 27607 7588 27611 7644
rect 27611 7588 27667 7644
rect 27667 7588 27671 7644
rect 27607 7584 27671 7588
rect 31219 8188 31283 8192
rect 31219 8132 31223 8188
rect 31223 8132 31279 8188
rect 31279 8132 31283 8188
rect 31219 8128 31283 8132
rect 31299 8188 31363 8192
rect 31299 8132 31303 8188
rect 31303 8132 31359 8188
rect 31359 8132 31363 8188
rect 31299 8128 31363 8132
rect 31379 8188 31443 8192
rect 31379 8132 31383 8188
rect 31383 8132 31439 8188
rect 31439 8132 31443 8188
rect 31379 8128 31443 8132
rect 31459 8188 31523 8192
rect 31459 8132 31463 8188
rect 31463 8132 31519 8188
rect 31519 8132 31523 8188
rect 31459 8128 31523 8132
rect 8104 7100 8168 7104
rect 8104 7044 8108 7100
rect 8108 7044 8164 7100
rect 8164 7044 8168 7100
rect 8104 7040 8168 7044
rect 8184 7100 8248 7104
rect 8184 7044 8188 7100
rect 8188 7044 8244 7100
rect 8244 7044 8248 7100
rect 8184 7040 8248 7044
rect 8264 7100 8328 7104
rect 8264 7044 8268 7100
rect 8268 7044 8324 7100
rect 8324 7044 8328 7100
rect 8264 7040 8328 7044
rect 8344 7100 8408 7104
rect 8344 7044 8348 7100
rect 8348 7044 8404 7100
rect 8404 7044 8408 7100
rect 8344 7040 8408 7044
rect 15809 7100 15873 7104
rect 15809 7044 15813 7100
rect 15813 7044 15869 7100
rect 15869 7044 15873 7100
rect 15809 7040 15873 7044
rect 15889 7100 15953 7104
rect 15889 7044 15893 7100
rect 15893 7044 15949 7100
rect 15949 7044 15953 7100
rect 15889 7040 15953 7044
rect 15969 7100 16033 7104
rect 15969 7044 15973 7100
rect 15973 7044 16029 7100
rect 16029 7044 16033 7100
rect 15969 7040 16033 7044
rect 16049 7100 16113 7104
rect 16049 7044 16053 7100
rect 16053 7044 16109 7100
rect 16109 7044 16113 7100
rect 16049 7040 16113 7044
rect 23514 7100 23578 7104
rect 23514 7044 23518 7100
rect 23518 7044 23574 7100
rect 23574 7044 23578 7100
rect 23514 7040 23578 7044
rect 23594 7100 23658 7104
rect 23594 7044 23598 7100
rect 23598 7044 23654 7100
rect 23654 7044 23658 7100
rect 23594 7040 23658 7044
rect 23674 7100 23738 7104
rect 23674 7044 23678 7100
rect 23678 7044 23734 7100
rect 23734 7044 23738 7100
rect 23674 7040 23738 7044
rect 23754 7100 23818 7104
rect 23754 7044 23758 7100
rect 23758 7044 23814 7100
rect 23814 7044 23818 7100
rect 23754 7040 23818 7044
rect 31219 7100 31283 7104
rect 31219 7044 31223 7100
rect 31223 7044 31279 7100
rect 31279 7044 31283 7100
rect 31219 7040 31283 7044
rect 31299 7100 31363 7104
rect 31299 7044 31303 7100
rect 31303 7044 31359 7100
rect 31359 7044 31363 7100
rect 31299 7040 31363 7044
rect 31379 7100 31443 7104
rect 31379 7044 31383 7100
rect 31383 7044 31439 7100
rect 31439 7044 31443 7100
rect 31379 7040 31443 7044
rect 31459 7100 31523 7104
rect 31459 7044 31463 7100
rect 31463 7044 31519 7100
rect 31519 7044 31523 7100
rect 31459 7040 31523 7044
rect 4252 6556 4316 6560
rect 4252 6500 4256 6556
rect 4256 6500 4312 6556
rect 4312 6500 4316 6556
rect 4252 6496 4316 6500
rect 4332 6556 4396 6560
rect 4332 6500 4336 6556
rect 4336 6500 4392 6556
rect 4392 6500 4396 6556
rect 4332 6496 4396 6500
rect 4412 6556 4476 6560
rect 4412 6500 4416 6556
rect 4416 6500 4472 6556
rect 4472 6500 4476 6556
rect 4412 6496 4476 6500
rect 4492 6556 4556 6560
rect 4492 6500 4496 6556
rect 4496 6500 4552 6556
rect 4552 6500 4556 6556
rect 4492 6496 4556 6500
rect 11957 6556 12021 6560
rect 11957 6500 11961 6556
rect 11961 6500 12017 6556
rect 12017 6500 12021 6556
rect 11957 6496 12021 6500
rect 12037 6556 12101 6560
rect 12037 6500 12041 6556
rect 12041 6500 12097 6556
rect 12097 6500 12101 6556
rect 12037 6496 12101 6500
rect 12117 6556 12181 6560
rect 12117 6500 12121 6556
rect 12121 6500 12177 6556
rect 12177 6500 12181 6556
rect 12117 6496 12181 6500
rect 12197 6556 12261 6560
rect 12197 6500 12201 6556
rect 12201 6500 12257 6556
rect 12257 6500 12261 6556
rect 12197 6496 12261 6500
rect 19662 6556 19726 6560
rect 19662 6500 19666 6556
rect 19666 6500 19722 6556
rect 19722 6500 19726 6556
rect 19662 6496 19726 6500
rect 19742 6556 19806 6560
rect 19742 6500 19746 6556
rect 19746 6500 19802 6556
rect 19802 6500 19806 6556
rect 19742 6496 19806 6500
rect 19822 6556 19886 6560
rect 19822 6500 19826 6556
rect 19826 6500 19882 6556
rect 19882 6500 19886 6556
rect 19822 6496 19886 6500
rect 19902 6556 19966 6560
rect 19902 6500 19906 6556
rect 19906 6500 19962 6556
rect 19962 6500 19966 6556
rect 19902 6496 19966 6500
rect 27367 6556 27431 6560
rect 27367 6500 27371 6556
rect 27371 6500 27427 6556
rect 27427 6500 27431 6556
rect 27367 6496 27431 6500
rect 27447 6556 27511 6560
rect 27447 6500 27451 6556
rect 27451 6500 27507 6556
rect 27507 6500 27511 6556
rect 27447 6496 27511 6500
rect 27527 6556 27591 6560
rect 27527 6500 27531 6556
rect 27531 6500 27587 6556
rect 27587 6500 27591 6556
rect 27527 6496 27591 6500
rect 27607 6556 27671 6560
rect 27607 6500 27611 6556
rect 27611 6500 27667 6556
rect 27667 6500 27671 6556
rect 27607 6496 27671 6500
rect 8104 6012 8168 6016
rect 8104 5956 8108 6012
rect 8108 5956 8164 6012
rect 8164 5956 8168 6012
rect 8104 5952 8168 5956
rect 8184 6012 8248 6016
rect 8184 5956 8188 6012
rect 8188 5956 8244 6012
rect 8244 5956 8248 6012
rect 8184 5952 8248 5956
rect 8264 6012 8328 6016
rect 8264 5956 8268 6012
rect 8268 5956 8324 6012
rect 8324 5956 8328 6012
rect 8264 5952 8328 5956
rect 8344 6012 8408 6016
rect 8344 5956 8348 6012
rect 8348 5956 8404 6012
rect 8404 5956 8408 6012
rect 8344 5952 8408 5956
rect 15809 6012 15873 6016
rect 15809 5956 15813 6012
rect 15813 5956 15869 6012
rect 15869 5956 15873 6012
rect 15809 5952 15873 5956
rect 15889 6012 15953 6016
rect 15889 5956 15893 6012
rect 15893 5956 15949 6012
rect 15949 5956 15953 6012
rect 15889 5952 15953 5956
rect 15969 6012 16033 6016
rect 15969 5956 15973 6012
rect 15973 5956 16029 6012
rect 16029 5956 16033 6012
rect 15969 5952 16033 5956
rect 16049 6012 16113 6016
rect 16049 5956 16053 6012
rect 16053 5956 16109 6012
rect 16109 5956 16113 6012
rect 16049 5952 16113 5956
rect 23514 6012 23578 6016
rect 23514 5956 23518 6012
rect 23518 5956 23574 6012
rect 23574 5956 23578 6012
rect 23514 5952 23578 5956
rect 23594 6012 23658 6016
rect 23594 5956 23598 6012
rect 23598 5956 23654 6012
rect 23654 5956 23658 6012
rect 23594 5952 23658 5956
rect 23674 6012 23738 6016
rect 23674 5956 23678 6012
rect 23678 5956 23734 6012
rect 23734 5956 23738 6012
rect 23674 5952 23738 5956
rect 23754 6012 23818 6016
rect 23754 5956 23758 6012
rect 23758 5956 23814 6012
rect 23814 5956 23818 6012
rect 23754 5952 23818 5956
rect 31219 6012 31283 6016
rect 31219 5956 31223 6012
rect 31223 5956 31279 6012
rect 31279 5956 31283 6012
rect 31219 5952 31283 5956
rect 31299 6012 31363 6016
rect 31299 5956 31303 6012
rect 31303 5956 31359 6012
rect 31359 5956 31363 6012
rect 31299 5952 31363 5956
rect 31379 6012 31443 6016
rect 31379 5956 31383 6012
rect 31383 5956 31439 6012
rect 31439 5956 31443 6012
rect 31379 5952 31443 5956
rect 31459 6012 31523 6016
rect 31459 5956 31463 6012
rect 31463 5956 31519 6012
rect 31519 5956 31523 6012
rect 31459 5952 31523 5956
rect 4252 5468 4316 5472
rect 4252 5412 4256 5468
rect 4256 5412 4312 5468
rect 4312 5412 4316 5468
rect 4252 5408 4316 5412
rect 4332 5468 4396 5472
rect 4332 5412 4336 5468
rect 4336 5412 4392 5468
rect 4392 5412 4396 5468
rect 4332 5408 4396 5412
rect 4412 5468 4476 5472
rect 4412 5412 4416 5468
rect 4416 5412 4472 5468
rect 4472 5412 4476 5468
rect 4412 5408 4476 5412
rect 4492 5468 4556 5472
rect 4492 5412 4496 5468
rect 4496 5412 4552 5468
rect 4552 5412 4556 5468
rect 4492 5408 4556 5412
rect 11957 5468 12021 5472
rect 11957 5412 11961 5468
rect 11961 5412 12017 5468
rect 12017 5412 12021 5468
rect 11957 5408 12021 5412
rect 12037 5468 12101 5472
rect 12037 5412 12041 5468
rect 12041 5412 12097 5468
rect 12097 5412 12101 5468
rect 12037 5408 12101 5412
rect 12117 5468 12181 5472
rect 12117 5412 12121 5468
rect 12121 5412 12177 5468
rect 12177 5412 12181 5468
rect 12117 5408 12181 5412
rect 12197 5468 12261 5472
rect 12197 5412 12201 5468
rect 12201 5412 12257 5468
rect 12257 5412 12261 5468
rect 12197 5408 12261 5412
rect 19662 5468 19726 5472
rect 19662 5412 19666 5468
rect 19666 5412 19722 5468
rect 19722 5412 19726 5468
rect 19662 5408 19726 5412
rect 19742 5468 19806 5472
rect 19742 5412 19746 5468
rect 19746 5412 19802 5468
rect 19802 5412 19806 5468
rect 19742 5408 19806 5412
rect 19822 5468 19886 5472
rect 19822 5412 19826 5468
rect 19826 5412 19882 5468
rect 19882 5412 19886 5468
rect 19822 5408 19886 5412
rect 19902 5468 19966 5472
rect 19902 5412 19906 5468
rect 19906 5412 19962 5468
rect 19962 5412 19966 5468
rect 19902 5408 19966 5412
rect 27367 5468 27431 5472
rect 27367 5412 27371 5468
rect 27371 5412 27427 5468
rect 27427 5412 27431 5468
rect 27367 5408 27431 5412
rect 27447 5468 27511 5472
rect 27447 5412 27451 5468
rect 27451 5412 27507 5468
rect 27507 5412 27511 5468
rect 27447 5408 27511 5412
rect 27527 5468 27591 5472
rect 27527 5412 27531 5468
rect 27531 5412 27587 5468
rect 27587 5412 27591 5468
rect 27527 5408 27591 5412
rect 27607 5468 27671 5472
rect 27607 5412 27611 5468
rect 27611 5412 27667 5468
rect 27667 5412 27671 5468
rect 27607 5408 27671 5412
rect 8104 4924 8168 4928
rect 8104 4868 8108 4924
rect 8108 4868 8164 4924
rect 8164 4868 8168 4924
rect 8104 4864 8168 4868
rect 8184 4924 8248 4928
rect 8184 4868 8188 4924
rect 8188 4868 8244 4924
rect 8244 4868 8248 4924
rect 8184 4864 8248 4868
rect 8264 4924 8328 4928
rect 8264 4868 8268 4924
rect 8268 4868 8324 4924
rect 8324 4868 8328 4924
rect 8264 4864 8328 4868
rect 8344 4924 8408 4928
rect 8344 4868 8348 4924
rect 8348 4868 8404 4924
rect 8404 4868 8408 4924
rect 8344 4864 8408 4868
rect 15809 4924 15873 4928
rect 15809 4868 15813 4924
rect 15813 4868 15869 4924
rect 15869 4868 15873 4924
rect 15809 4864 15873 4868
rect 15889 4924 15953 4928
rect 15889 4868 15893 4924
rect 15893 4868 15949 4924
rect 15949 4868 15953 4924
rect 15889 4864 15953 4868
rect 15969 4924 16033 4928
rect 15969 4868 15973 4924
rect 15973 4868 16029 4924
rect 16029 4868 16033 4924
rect 15969 4864 16033 4868
rect 16049 4924 16113 4928
rect 16049 4868 16053 4924
rect 16053 4868 16109 4924
rect 16109 4868 16113 4924
rect 16049 4864 16113 4868
rect 20668 4524 20732 4588
rect 23514 4924 23578 4928
rect 23514 4868 23518 4924
rect 23518 4868 23574 4924
rect 23574 4868 23578 4924
rect 23514 4864 23578 4868
rect 23594 4924 23658 4928
rect 23594 4868 23598 4924
rect 23598 4868 23654 4924
rect 23654 4868 23658 4924
rect 23594 4864 23658 4868
rect 23674 4924 23738 4928
rect 23674 4868 23678 4924
rect 23678 4868 23734 4924
rect 23734 4868 23738 4924
rect 23674 4864 23738 4868
rect 23754 4924 23818 4928
rect 23754 4868 23758 4924
rect 23758 4868 23814 4924
rect 23814 4868 23818 4924
rect 23754 4864 23818 4868
rect 31219 4924 31283 4928
rect 31219 4868 31223 4924
rect 31223 4868 31279 4924
rect 31279 4868 31283 4924
rect 31219 4864 31283 4868
rect 31299 4924 31363 4928
rect 31299 4868 31303 4924
rect 31303 4868 31359 4924
rect 31359 4868 31363 4924
rect 31299 4864 31363 4868
rect 31379 4924 31443 4928
rect 31379 4868 31383 4924
rect 31383 4868 31439 4924
rect 31439 4868 31443 4924
rect 31379 4864 31443 4868
rect 31459 4924 31523 4928
rect 31459 4868 31463 4924
rect 31463 4868 31519 4924
rect 31519 4868 31523 4924
rect 31459 4864 31523 4868
rect 4252 4380 4316 4384
rect 4252 4324 4256 4380
rect 4256 4324 4312 4380
rect 4312 4324 4316 4380
rect 4252 4320 4316 4324
rect 4332 4380 4396 4384
rect 4332 4324 4336 4380
rect 4336 4324 4392 4380
rect 4392 4324 4396 4380
rect 4332 4320 4396 4324
rect 4412 4380 4476 4384
rect 4412 4324 4416 4380
rect 4416 4324 4472 4380
rect 4472 4324 4476 4380
rect 4412 4320 4476 4324
rect 4492 4380 4556 4384
rect 4492 4324 4496 4380
rect 4496 4324 4552 4380
rect 4552 4324 4556 4380
rect 4492 4320 4556 4324
rect 11957 4380 12021 4384
rect 11957 4324 11961 4380
rect 11961 4324 12017 4380
rect 12017 4324 12021 4380
rect 11957 4320 12021 4324
rect 12037 4380 12101 4384
rect 12037 4324 12041 4380
rect 12041 4324 12097 4380
rect 12097 4324 12101 4380
rect 12037 4320 12101 4324
rect 12117 4380 12181 4384
rect 12117 4324 12121 4380
rect 12121 4324 12177 4380
rect 12177 4324 12181 4380
rect 12117 4320 12181 4324
rect 12197 4380 12261 4384
rect 12197 4324 12201 4380
rect 12201 4324 12257 4380
rect 12257 4324 12261 4380
rect 12197 4320 12261 4324
rect 19662 4380 19726 4384
rect 19662 4324 19666 4380
rect 19666 4324 19722 4380
rect 19722 4324 19726 4380
rect 19662 4320 19726 4324
rect 19742 4380 19806 4384
rect 19742 4324 19746 4380
rect 19746 4324 19802 4380
rect 19802 4324 19806 4380
rect 19742 4320 19806 4324
rect 19822 4380 19886 4384
rect 19822 4324 19826 4380
rect 19826 4324 19882 4380
rect 19882 4324 19886 4380
rect 19822 4320 19886 4324
rect 19902 4380 19966 4384
rect 19902 4324 19906 4380
rect 19906 4324 19962 4380
rect 19962 4324 19966 4380
rect 19902 4320 19966 4324
rect 27367 4380 27431 4384
rect 27367 4324 27371 4380
rect 27371 4324 27427 4380
rect 27427 4324 27431 4380
rect 27367 4320 27431 4324
rect 27447 4380 27511 4384
rect 27447 4324 27451 4380
rect 27451 4324 27507 4380
rect 27507 4324 27511 4380
rect 27447 4320 27511 4324
rect 27527 4380 27591 4384
rect 27527 4324 27531 4380
rect 27531 4324 27587 4380
rect 27587 4324 27591 4380
rect 27527 4320 27591 4324
rect 27607 4380 27671 4384
rect 27607 4324 27611 4380
rect 27611 4324 27667 4380
rect 27667 4324 27671 4380
rect 27607 4320 27671 4324
rect 8104 3836 8168 3840
rect 8104 3780 8108 3836
rect 8108 3780 8164 3836
rect 8164 3780 8168 3836
rect 8104 3776 8168 3780
rect 8184 3836 8248 3840
rect 8184 3780 8188 3836
rect 8188 3780 8244 3836
rect 8244 3780 8248 3836
rect 8184 3776 8248 3780
rect 8264 3836 8328 3840
rect 8264 3780 8268 3836
rect 8268 3780 8324 3836
rect 8324 3780 8328 3836
rect 8264 3776 8328 3780
rect 8344 3836 8408 3840
rect 8344 3780 8348 3836
rect 8348 3780 8404 3836
rect 8404 3780 8408 3836
rect 8344 3776 8408 3780
rect 15809 3836 15873 3840
rect 15809 3780 15813 3836
rect 15813 3780 15869 3836
rect 15869 3780 15873 3836
rect 15809 3776 15873 3780
rect 15889 3836 15953 3840
rect 15889 3780 15893 3836
rect 15893 3780 15949 3836
rect 15949 3780 15953 3836
rect 15889 3776 15953 3780
rect 15969 3836 16033 3840
rect 15969 3780 15973 3836
rect 15973 3780 16029 3836
rect 16029 3780 16033 3836
rect 15969 3776 16033 3780
rect 16049 3836 16113 3840
rect 16049 3780 16053 3836
rect 16053 3780 16109 3836
rect 16109 3780 16113 3836
rect 16049 3776 16113 3780
rect 23514 3836 23578 3840
rect 23514 3780 23518 3836
rect 23518 3780 23574 3836
rect 23574 3780 23578 3836
rect 23514 3776 23578 3780
rect 23594 3836 23658 3840
rect 23594 3780 23598 3836
rect 23598 3780 23654 3836
rect 23654 3780 23658 3836
rect 23594 3776 23658 3780
rect 23674 3836 23738 3840
rect 23674 3780 23678 3836
rect 23678 3780 23734 3836
rect 23734 3780 23738 3836
rect 23674 3776 23738 3780
rect 23754 3836 23818 3840
rect 23754 3780 23758 3836
rect 23758 3780 23814 3836
rect 23814 3780 23818 3836
rect 23754 3776 23818 3780
rect 31219 3836 31283 3840
rect 31219 3780 31223 3836
rect 31223 3780 31279 3836
rect 31279 3780 31283 3836
rect 31219 3776 31283 3780
rect 31299 3836 31363 3840
rect 31299 3780 31303 3836
rect 31303 3780 31359 3836
rect 31359 3780 31363 3836
rect 31299 3776 31363 3780
rect 31379 3836 31443 3840
rect 31379 3780 31383 3836
rect 31383 3780 31439 3836
rect 31439 3780 31443 3836
rect 31379 3776 31443 3780
rect 31459 3836 31523 3840
rect 31459 3780 31463 3836
rect 31463 3780 31519 3836
rect 31519 3780 31523 3836
rect 31459 3776 31523 3780
rect 4252 3292 4316 3296
rect 4252 3236 4256 3292
rect 4256 3236 4312 3292
rect 4312 3236 4316 3292
rect 4252 3232 4316 3236
rect 4332 3292 4396 3296
rect 4332 3236 4336 3292
rect 4336 3236 4392 3292
rect 4392 3236 4396 3292
rect 4332 3232 4396 3236
rect 4412 3292 4476 3296
rect 4412 3236 4416 3292
rect 4416 3236 4472 3292
rect 4472 3236 4476 3292
rect 4412 3232 4476 3236
rect 4492 3292 4556 3296
rect 4492 3236 4496 3292
rect 4496 3236 4552 3292
rect 4552 3236 4556 3292
rect 4492 3232 4556 3236
rect 11957 3292 12021 3296
rect 11957 3236 11961 3292
rect 11961 3236 12017 3292
rect 12017 3236 12021 3292
rect 11957 3232 12021 3236
rect 12037 3292 12101 3296
rect 12037 3236 12041 3292
rect 12041 3236 12097 3292
rect 12097 3236 12101 3292
rect 12037 3232 12101 3236
rect 12117 3292 12181 3296
rect 12117 3236 12121 3292
rect 12121 3236 12177 3292
rect 12177 3236 12181 3292
rect 12117 3232 12181 3236
rect 12197 3292 12261 3296
rect 12197 3236 12201 3292
rect 12201 3236 12257 3292
rect 12257 3236 12261 3292
rect 12197 3232 12261 3236
rect 19662 3292 19726 3296
rect 19662 3236 19666 3292
rect 19666 3236 19722 3292
rect 19722 3236 19726 3292
rect 19662 3232 19726 3236
rect 19742 3292 19806 3296
rect 19742 3236 19746 3292
rect 19746 3236 19802 3292
rect 19802 3236 19806 3292
rect 19742 3232 19806 3236
rect 19822 3292 19886 3296
rect 19822 3236 19826 3292
rect 19826 3236 19882 3292
rect 19882 3236 19886 3292
rect 19822 3232 19886 3236
rect 19902 3292 19966 3296
rect 19902 3236 19906 3292
rect 19906 3236 19962 3292
rect 19962 3236 19966 3292
rect 19902 3232 19966 3236
rect 27367 3292 27431 3296
rect 27367 3236 27371 3292
rect 27371 3236 27427 3292
rect 27427 3236 27431 3292
rect 27367 3232 27431 3236
rect 27447 3292 27511 3296
rect 27447 3236 27451 3292
rect 27451 3236 27507 3292
rect 27507 3236 27511 3292
rect 27447 3232 27511 3236
rect 27527 3292 27591 3296
rect 27527 3236 27531 3292
rect 27531 3236 27587 3292
rect 27587 3236 27591 3292
rect 27527 3232 27591 3236
rect 27607 3292 27671 3296
rect 27607 3236 27611 3292
rect 27611 3236 27667 3292
rect 27667 3236 27671 3292
rect 27607 3232 27671 3236
rect 8104 2748 8168 2752
rect 8104 2692 8108 2748
rect 8108 2692 8164 2748
rect 8164 2692 8168 2748
rect 8104 2688 8168 2692
rect 8184 2748 8248 2752
rect 8184 2692 8188 2748
rect 8188 2692 8244 2748
rect 8244 2692 8248 2748
rect 8184 2688 8248 2692
rect 8264 2748 8328 2752
rect 8264 2692 8268 2748
rect 8268 2692 8324 2748
rect 8324 2692 8328 2748
rect 8264 2688 8328 2692
rect 8344 2748 8408 2752
rect 8344 2692 8348 2748
rect 8348 2692 8404 2748
rect 8404 2692 8408 2748
rect 8344 2688 8408 2692
rect 15809 2748 15873 2752
rect 15809 2692 15813 2748
rect 15813 2692 15869 2748
rect 15869 2692 15873 2748
rect 15809 2688 15873 2692
rect 15889 2748 15953 2752
rect 15889 2692 15893 2748
rect 15893 2692 15949 2748
rect 15949 2692 15953 2748
rect 15889 2688 15953 2692
rect 15969 2748 16033 2752
rect 15969 2692 15973 2748
rect 15973 2692 16029 2748
rect 16029 2692 16033 2748
rect 15969 2688 16033 2692
rect 16049 2748 16113 2752
rect 16049 2692 16053 2748
rect 16053 2692 16109 2748
rect 16109 2692 16113 2748
rect 16049 2688 16113 2692
rect 23514 2748 23578 2752
rect 23514 2692 23518 2748
rect 23518 2692 23574 2748
rect 23574 2692 23578 2748
rect 23514 2688 23578 2692
rect 23594 2748 23658 2752
rect 23594 2692 23598 2748
rect 23598 2692 23654 2748
rect 23654 2692 23658 2748
rect 23594 2688 23658 2692
rect 23674 2748 23738 2752
rect 23674 2692 23678 2748
rect 23678 2692 23734 2748
rect 23734 2692 23738 2748
rect 23674 2688 23738 2692
rect 23754 2748 23818 2752
rect 23754 2692 23758 2748
rect 23758 2692 23814 2748
rect 23814 2692 23818 2748
rect 23754 2688 23818 2692
rect 31219 2748 31283 2752
rect 31219 2692 31223 2748
rect 31223 2692 31279 2748
rect 31279 2692 31283 2748
rect 31219 2688 31283 2692
rect 31299 2748 31363 2752
rect 31299 2692 31303 2748
rect 31303 2692 31359 2748
rect 31359 2692 31363 2748
rect 31299 2688 31363 2692
rect 31379 2748 31443 2752
rect 31379 2692 31383 2748
rect 31383 2692 31439 2748
rect 31439 2692 31443 2748
rect 31379 2688 31443 2692
rect 31459 2748 31523 2752
rect 31459 2692 31463 2748
rect 31463 2692 31519 2748
rect 31519 2692 31523 2748
rect 31459 2688 31523 2692
rect 4252 2204 4316 2208
rect 4252 2148 4256 2204
rect 4256 2148 4312 2204
rect 4312 2148 4316 2204
rect 4252 2144 4316 2148
rect 4332 2204 4396 2208
rect 4332 2148 4336 2204
rect 4336 2148 4392 2204
rect 4392 2148 4396 2204
rect 4332 2144 4396 2148
rect 4412 2204 4476 2208
rect 4412 2148 4416 2204
rect 4416 2148 4472 2204
rect 4472 2148 4476 2204
rect 4412 2144 4476 2148
rect 4492 2204 4556 2208
rect 4492 2148 4496 2204
rect 4496 2148 4552 2204
rect 4552 2148 4556 2204
rect 4492 2144 4556 2148
rect 11957 2204 12021 2208
rect 11957 2148 11961 2204
rect 11961 2148 12017 2204
rect 12017 2148 12021 2204
rect 11957 2144 12021 2148
rect 12037 2204 12101 2208
rect 12037 2148 12041 2204
rect 12041 2148 12097 2204
rect 12097 2148 12101 2204
rect 12037 2144 12101 2148
rect 12117 2204 12181 2208
rect 12117 2148 12121 2204
rect 12121 2148 12177 2204
rect 12177 2148 12181 2204
rect 12117 2144 12181 2148
rect 12197 2204 12261 2208
rect 12197 2148 12201 2204
rect 12201 2148 12257 2204
rect 12257 2148 12261 2204
rect 12197 2144 12261 2148
rect 19662 2204 19726 2208
rect 19662 2148 19666 2204
rect 19666 2148 19722 2204
rect 19722 2148 19726 2204
rect 19662 2144 19726 2148
rect 19742 2204 19806 2208
rect 19742 2148 19746 2204
rect 19746 2148 19802 2204
rect 19802 2148 19806 2204
rect 19742 2144 19806 2148
rect 19822 2204 19886 2208
rect 19822 2148 19826 2204
rect 19826 2148 19882 2204
rect 19882 2148 19886 2204
rect 19822 2144 19886 2148
rect 19902 2204 19966 2208
rect 19902 2148 19906 2204
rect 19906 2148 19962 2204
rect 19962 2148 19966 2204
rect 19902 2144 19966 2148
rect 27367 2204 27431 2208
rect 27367 2148 27371 2204
rect 27371 2148 27427 2204
rect 27427 2148 27431 2204
rect 27367 2144 27431 2148
rect 27447 2204 27511 2208
rect 27447 2148 27451 2204
rect 27451 2148 27507 2204
rect 27507 2148 27511 2204
rect 27447 2144 27511 2148
rect 27527 2204 27591 2208
rect 27527 2148 27531 2204
rect 27531 2148 27587 2204
rect 27587 2148 27591 2204
rect 27527 2144 27591 2148
rect 27607 2204 27671 2208
rect 27607 2148 27611 2204
rect 27611 2148 27667 2204
rect 27667 2148 27671 2204
rect 27607 2144 27671 2148
rect 8104 1660 8168 1664
rect 8104 1604 8108 1660
rect 8108 1604 8164 1660
rect 8164 1604 8168 1660
rect 8104 1600 8168 1604
rect 8184 1660 8248 1664
rect 8184 1604 8188 1660
rect 8188 1604 8244 1660
rect 8244 1604 8248 1660
rect 8184 1600 8248 1604
rect 8264 1660 8328 1664
rect 8264 1604 8268 1660
rect 8268 1604 8324 1660
rect 8324 1604 8328 1660
rect 8264 1600 8328 1604
rect 8344 1660 8408 1664
rect 8344 1604 8348 1660
rect 8348 1604 8404 1660
rect 8404 1604 8408 1660
rect 8344 1600 8408 1604
rect 15809 1660 15873 1664
rect 15809 1604 15813 1660
rect 15813 1604 15869 1660
rect 15869 1604 15873 1660
rect 15809 1600 15873 1604
rect 15889 1660 15953 1664
rect 15889 1604 15893 1660
rect 15893 1604 15949 1660
rect 15949 1604 15953 1660
rect 15889 1600 15953 1604
rect 15969 1660 16033 1664
rect 15969 1604 15973 1660
rect 15973 1604 16029 1660
rect 16029 1604 16033 1660
rect 15969 1600 16033 1604
rect 16049 1660 16113 1664
rect 16049 1604 16053 1660
rect 16053 1604 16109 1660
rect 16109 1604 16113 1660
rect 16049 1600 16113 1604
rect 23514 1660 23578 1664
rect 23514 1604 23518 1660
rect 23518 1604 23574 1660
rect 23574 1604 23578 1660
rect 23514 1600 23578 1604
rect 23594 1660 23658 1664
rect 23594 1604 23598 1660
rect 23598 1604 23654 1660
rect 23654 1604 23658 1660
rect 23594 1600 23658 1604
rect 23674 1660 23738 1664
rect 23674 1604 23678 1660
rect 23678 1604 23734 1660
rect 23734 1604 23738 1660
rect 23674 1600 23738 1604
rect 23754 1660 23818 1664
rect 23754 1604 23758 1660
rect 23758 1604 23814 1660
rect 23814 1604 23818 1660
rect 23754 1600 23818 1604
rect 31219 1660 31283 1664
rect 31219 1604 31223 1660
rect 31223 1604 31279 1660
rect 31279 1604 31283 1660
rect 31219 1600 31283 1604
rect 31299 1660 31363 1664
rect 31299 1604 31303 1660
rect 31303 1604 31359 1660
rect 31359 1604 31363 1660
rect 31299 1600 31363 1604
rect 31379 1660 31443 1664
rect 31379 1604 31383 1660
rect 31383 1604 31439 1660
rect 31439 1604 31443 1660
rect 31379 1600 31443 1604
rect 31459 1660 31523 1664
rect 31459 1604 31463 1660
rect 31463 1604 31519 1660
rect 31519 1604 31523 1660
rect 31459 1600 31523 1604
rect 4252 1116 4316 1120
rect 4252 1060 4256 1116
rect 4256 1060 4312 1116
rect 4312 1060 4316 1116
rect 4252 1056 4316 1060
rect 4332 1116 4396 1120
rect 4332 1060 4336 1116
rect 4336 1060 4392 1116
rect 4392 1060 4396 1116
rect 4332 1056 4396 1060
rect 4412 1116 4476 1120
rect 4412 1060 4416 1116
rect 4416 1060 4472 1116
rect 4472 1060 4476 1116
rect 4412 1056 4476 1060
rect 4492 1116 4556 1120
rect 4492 1060 4496 1116
rect 4496 1060 4552 1116
rect 4552 1060 4556 1116
rect 4492 1056 4556 1060
rect 11957 1116 12021 1120
rect 11957 1060 11961 1116
rect 11961 1060 12017 1116
rect 12017 1060 12021 1116
rect 11957 1056 12021 1060
rect 12037 1116 12101 1120
rect 12037 1060 12041 1116
rect 12041 1060 12097 1116
rect 12097 1060 12101 1116
rect 12037 1056 12101 1060
rect 12117 1116 12181 1120
rect 12117 1060 12121 1116
rect 12121 1060 12177 1116
rect 12177 1060 12181 1116
rect 12117 1056 12181 1060
rect 12197 1116 12261 1120
rect 12197 1060 12201 1116
rect 12201 1060 12257 1116
rect 12257 1060 12261 1116
rect 12197 1056 12261 1060
rect 19662 1116 19726 1120
rect 19662 1060 19666 1116
rect 19666 1060 19722 1116
rect 19722 1060 19726 1116
rect 19662 1056 19726 1060
rect 19742 1116 19806 1120
rect 19742 1060 19746 1116
rect 19746 1060 19802 1116
rect 19802 1060 19806 1116
rect 19742 1056 19806 1060
rect 19822 1116 19886 1120
rect 19822 1060 19826 1116
rect 19826 1060 19882 1116
rect 19882 1060 19886 1116
rect 19822 1056 19886 1060
rect 19902 1116 19966 1120
rect 19902 1060 19906 1116
rect 19906 1060 19962 1116
rect 19962 1060 19966 1116
rect 19902 1056 19966 1060
rect 27367 1116 27431 1120
rect 27367 1060 27371 1116
rect 27371 1060 27427 1116
rect 27427 1060 27431 1116
rect 27367 1056 27431 1060
rect 27447 1116 27511 1120
rect 27447 1060 27451 1116
rect 27451 1060 27507 1116
rect 27507 1060 27511 1116
rect 27447 1056 27511 1060
rect 27527 1116 27591 1120
rect 27527 1060 27531 1116
rect 27531 1060 27587 1116
rect 27587 1060 27591 1116
rect 27527 1056 27591 1060
rect 27607 1116 27671 1120
rect 27607 1060 27611 1116
rect 27611 1060 27667 1116
rect 27667 1060 27671 1116
rect 27607 1056 27671 1060
rect 8104 572 8168 576
rect 8104 516 8108 572
rect 8108 516 8164 572
rect 8164 516 8168 572
rect 8104 512 8168 516
rect 8184 572 8248 576
rect 8184 516 8188 572
rect 8188 516 8244 572
rect 8244 516 8248 572
rect 8184 512 8248 516
rect 8264 572 8328 576
rect 8264 516 8268 572
rect 8268 516 8324 572
rect 8324 516 8328 572
rect 8264 512 8328 516
rect 8344 572 8408 576
rect 8344 516 8348 572
rect 8348 516 8404 572
rect 8404 516 8408 572
rect 8344 512 8408 516
rect 15809 572 15873 576
rect 15809 516 15813 572
rect 15813 516 15869 572
rect 15869 516 15873 572
rect 15809 512 15873 516
rect 15889 572 15953 576
rect 15889 516 15893 572
rect 15893 516 15949 572
rect 15949 516 15953 572
rect 15889 512 15953 516
rect 15969 572 16033 576
rect 15969 516 15973 572
rect 15973 516 16029 572
rect 16029 516 16033 572
rect 15969 512 16033 516
rect 16049 572 16113 576
rect 16049 516 16053 572
rect 16053 516 16109 572
rect 16109 516 16113 572
rect 16049 512 16113 516
rect 23514 572 23578 576
rect 23514 516 23518 572
rect 23518 516 23574 572
rect 23574 516 23578 572
rect 23514 512 23578 516
rect 23594 572 23658 576
rect 23594 516 23598 572
rect 23598 516 23654 572
rect 23654 516 23658 572
rect 23594 512 23658 516
rect 23674 572 23738 576
rect 23674 516 23678 572
rect 23678 516 23734 572
rect 23734 516 23738 572
rect 23674 512 23738 516
rect 23754 572 23818 576
rect 23754 516 23758 572
rect 23758 516 23814 572
rect 23814 516 23818 572
rect 23754 512 23818 516
rect 31219 572 31283 576
rect 31219 516 31223 572
rect 31223 516 31279 572
rect 31279 516 31283 572
rect 31219 512 31283 516
rect 31299 572 31363 576
rect 31299 516 31303 572
rect 31303 516 31359 572
rect 31359 516 31363 572
rect 31299 512 31363 516
rect 31379 572 31443 576
rect 31379 516 31383 572
rect 31383 516 31439 572
rect 31439 516 31443 572
rect 31379 512 31443 516
rect 31459 572 31523 576
rect 31459 516 31463 572
rect 31463 516 31519 572
rect 31519 516 31523 572
rect 31459 512 31523 516
rect 15148 308 15212 372
<< metal4 >>
rect 4244 18528 4564 19088
rect 4244 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4564 18528
rect 4244 17440 4564 18464
rect 4244 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4564 17440
rect 4244 16352 4564 17376
rect 4244 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4564 16352
rect 4244 15264 4564 16288
rect 4244 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4564 15264
rect 4244 14176 4564 15200
rect 4244 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4564 14176
rect 4244 13088 4564 14112
rect 4244 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4564 13088
rect 4244 12000 4564 13024
rect 4244 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4564 12000
rect 4244 10912 4564 11936
rect 4244 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4564 10912
rect 4244 9824 4564 10848
rect 4244 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4564 9824
rect 4244 8736 4564 9760
rect 4244 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4564 8736
rect 4244 7648 4564 8672
rect 4244 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4564 7648
rect 4244 6560 4564 7584
rect 4244 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4564 6560
rect 4244 5472 4564 6496
rect 4244 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4564 5472
rect 4244 4384 4564 5408
rect 4244 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4564 4384
rect 4244 3296 4564 4320
rect 4244 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4564 3296
rect 4244 2208 4564 3232
rect 4244 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4564 2208
rect 4244 1120 4564 2144
rect 4244 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4564 1120
rect 4244 496 4564 1056
rect 8096 19072 8416 19088
rect 8096 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8416 19072
rect 8096 17984 8416 19008
rect 11651 18732 11717 18733
rect 11651 18668 11652 18732
rect 11716 18668 11717 18732
rect 11651 18667 11717 18668
rect 8096 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8416 17984
rect 8096 16896 8416 17920
rect 11283 16964 11349 16965
rect 11283 16900 11284 16964
rect 11348 16900 11349 16964
rect 11283 16899 11349 16900
rect 8096 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8416 16896
rect 8096 15808 8416 16832
rect 10363 16828 10429 16829
rect 10363 16764 10364 16828
rect 10428 16764 10429 16828
rect 10363 16763 10429 16764
rect 9995 16556 10061 16557
rect 9995 16492 9996 16556
rect 10060 16492 10061 16556
rect 9995 16491 10061 16492
rect 8096 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8416 15808
rect 8096 14720 8416 15744
rect 9811 15740 9877 15741
rect 9811 15676 9812 15740
rect 9876 15676 9877 15740
rect 9811 15675 9877 15676
rect 9814 15061 9874 15675
rect 9998 15197 10058 16491
rect 10366 15333 10426 16763
rect 10547 16556 10613 16557
rect 10547 16492 10548 16556
rect 10612 16492 10613 16556
rect 10547 16491 10613 16492
rect 10731 16556 10797 16557
rect 10731 16492 10732 16556
rect 10796 16492 10797 16556
rect 10731 16491 10797 16492
rect 10363 15332 10429 15333
rect 10363 15268 10364 15332
rect 10428 15268 10429 15332
rect 10363 15267 10429 15268
rect 9995 15196 10061 15197
rect 9995 15132 9996 15196
rect 10060 15132 10061 15196
rect 9995 15131 10061 15132
rect 9811 15060 9877 15061
rect 9811 14996 9812 15060
rect 9876 14996 9877 15060
rect 9811 14995 9877 14996
rect 10550 14789 10610 16491
rect 10734 15333 10794 16491
rect 11099 15740 11165 15741
rect 11099 15676 11100 15740
rect 11164 15676 11165 15740
rect 11099 15675 11165 15676
rect 10731 15332 10797 15333
rect 10731 15268 10732 15332
rect 10796 15268 10797 15332
rect 10731 15267 10797 15268
rect 10547 14788 10613 14789
rect 10547 14724 10548 14788
rect 10612 14724 10613 14788
rect 10547 14723 10613 14724
rect 8096 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8416 14720
rect 8096 13632 8416 14656
rect 8096 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8416 13632
rect 8096 12544 8416 13568
rect 11102 13429 11162 15675
rect 11099 13428 11165 13429
rect 11099 13364 11100 13428
rect 11164 13364 11165 13428
rect 11099 13363 11165 13364
rect 11286 13021 11346 16899
rect 11654 13021 11714 18667
rect 11949 18528 12269 19088
rect 11949 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12269 18528
rect 11949 17440 12269 18464
rect 11949 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12269 17440
rect 11949 16352 12269 17376
rect 11949 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12269 16352
rect 11949 15264 12269 16288
rect 15801 19072 16121 19088
rect 15801 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16121 19072
rect 15801 17984 16121 19008
rect 15801 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16121 17984
rect 15801 16896 16121 17920
rect 19654 18528 19974 19088
rect 19654 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19974 18528
rect 19654 17440 19974 18464
rect 19654 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19974 17440
rect 19379 17100 19445 17101
rect 19379 17036 19380 17100
rect 19444 17036 19445 17100
rect 19379 17035 19445 17036
rect 15801 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16121 16896
rect 13307 16012 13373 16013
rect 13307 15948 13308 16012
rect 13372 15948 13373 16012
rect 13307 15947 13373 15948
rect 11949 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12269 15264
rect 11949 14176 12269 15200
rect 11949 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12269 14176
rect 11949 13088 12269 14112
rect 11949 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12269 13088
rect 11283 13020 11349 13021
rect 11283 12956 11284 13020
rect 11348 12956 11349 13020
rect 11283 12955 11349 12956
rect 11651 13020 11717 13021
rect 11651 12956 11652 13020
rect 11716 12956 11717 13020
rect 11651 12955 11717 12956
rect 8096 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8416 12544
rect 8096 11456 8416 12480
rect 8096 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8416 11456
rect 8096 10368 8416 11392
rect 8096 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8416 10368
rect 8096 9280 8416 10304
rect 8096 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8416 9280
rect 8096 8192 8416 9216
rect 8096 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8416 8192
rect 8096 7104 8416 8128
rect 8096 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8416 7104
rect 8096 6016 8416 7040
rect 8096 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8416 6016
rect 8096 4928 8416 5952
rect 8096 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8416 4928
rect 8096 3840 8416 4864
rect 8096 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8416 3840
rect 8096 2752 8416 3776
rect 8096 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8416 2752
rect 8096 1664 8416 2688
rect 8096 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8416 1664
rect 8096 576 8416 1600
rect 8096 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8416 576
rect 8096 496 8416 512
rect 11949 12000 12269 13024
rect 11949 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12269 12000
rect 11949 10912 12269 11936
rect 13310 10981 13370 15947
rect 15801 15808 16121 16832
rect 15801 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16121 15808
rect 15801 14720 16121 15744
rect 15801 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16121 14720
rect 15801 13632 16121 14656
rect 15801 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16121 13632
rect 15801 12544 16121 13568
rect 15801 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16121 12544
rect 15801 11456 16121 12480
rect 19382 11797 19442 17035
rect 19654 16352 19974 17376
rect 19654 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19974 16352
rect 19654 15264 19974 16288
rect 23506 19072 23826 19088
rect 23506 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23826 19072
rect 23506 17984 23826 19008
rect 23506 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23826 17984
rect 23506 16896 23826 17920
rect 23506 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23826 16896
rect 22323 16012 22389 16013
rect 22323 15948 22324 16012
rect 22388 15948 22389 16012
rect 22323 15947 22389 15948
rect 21955 15740 22021 15741
rect 21955 15676 21956 15740
rect 22020 15676 22021 15740
rect 21955 15675 22021 15676
rect 19654 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19974 15264
rect 19654 14176 19974 15200
rect 19654 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19974 14176
rect 19654 13088 19974 14112
rect 21958 13429 22018 15675
rect 22326 13701 22386 15947
rect 23506 15808 23826 16832
rect 27359 18528 27679 19088
rect 27359 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27679 18528
rect 27359 17440 27679 18464
rect 27359 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27679 17440
rect 27359 16352 27679 17376
rect 27359 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27679 16352
rect 23979 16012 24045 16013
rect 23979 15948 23980 16012
rect 24044 15948 24045 16012
rect 23979 15947 24045 15948
rect 23506 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23826 15808
rect 23243 15468 23309 15469
rect 23243 15404 23244 15468
rect 23308 15404 23309 15468
rect 23243 15403 23309 15404
rect 22323 13700 22389 13701
rect 22323 13636 22324 13700
rect 22388 13636 22389 13700
rect 22323 13635 22389 13636
rect 21955 13428 22021 13429
rect 21955 13364 21956 13428
rect 22020 13364 22021 13428
rect 21955 13363 22021 13364
rect 19654 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19974 13088
rect 19654 12000 19974 13024
rect 23246 12885 23306 15403
rect 23506 14720 23826 15744
rect 23506 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23826 14720
rect 23506 13632 23826 14656
rect 23506 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23826 13632
rect 23243 12884 23309 12885
rect 23243 12820 23244 12884
rect 23308 12820 23309 12884
rect 23243 12819 23309 12820
rect 19654 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19974 12000
rect 19379 11796 19445 11797
rect 19379 11732 19380 11796
rect 19444 11732 19445 11796
rect 19379 11731 19445 11732
rect 15801 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16121 11456
rect 13307 10980 13373 10981
rect 13307 10916 13308 10980
rect 13372 10916 13373 10980
rect 13307 10915 13373 10916
rect 11949 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12269 10912
rect 11949 9824 12269 10848
rect 11949 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12269 9824
rect 11949 8736 12269 9760
rect 11949 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12269 8736
rect 11949 7648 12269 8672
rect 15801 10368 16121 11392
rect 15801 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16121 10368
rect 15801 9280 16121 10304
rect 15801 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16121 9280
rect 15147 8396 15213 8397
rect 15147 8332 15148 8396
rect 15212 8332 15213 8396
rect 15147 8331 15213 8332
rect 11949 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12269 7648
rect 11949 6560 12269 7584
rect 11949 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12269 6560
rect 11949 5472 12269 6496
rect 11949 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12269 5472
rect 11949 4384 12269 5408
rect 11949 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12269 4384
rect 11949 3296 12269 4320
rect 11949 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12269 3296
rect 11949 2208 12269 3232
rect 11949 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12269 2208
rect 11949 1120 12269 2144
rect 11949 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12269 1120
rect 11949 496 12269 1056
rect 15150 373 15210 8331
rect 15801 8192 16121 9216
rect 15801 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16121 8192
rect 15801 7104 16121 8128
rect 15801 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16121 7104
rect 15801 6016 16121 7040
rect 15801 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16121 6016
rect 15801 4928 16121 5952
rect 15801 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16121 4928
rect 15801 3840 16121 4864
rect 15801 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16121 3840
rect 15801 2752 16121 3776
rect 15801 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16121 2752
rect 15801 1664 16121 2688
rect 15801 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16121 1664
rect 15801 576 16121 1600
rect 15801 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16121 576
rect 15801 496 16121 512
rect 19654 10912 19974 11936
rect 19654 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19974 10912
rect 19654 9824 19974 10848
rect 19654 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19974 9824
rect 19654 8736 19974 9760
rect 19654 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19974 8736
rect 19654 7648 19974 8672
rect 23506 12544 23826 13568
rect 23506 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23826 12544
rect 23506 11456 23826 12480
rect 23982 12341 24042 15947
rect 24899 15604 24965 15605
rect 24899 15540 24900 15604
rect 24964 15540 24965 15604
rect 24899 15539 24965 15540
rect 24902 13157 24962 15539
rect 27359 15264 27679 16288
rect 27359 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27679 15264
rect 27359 14176 27679 15200
rect 27359 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27679 14176
rect 24899 13156 24965 13157
rect 24899 13092 24900 13156
rect 24964 13092 24965 13156
rect 24899 13091 24965 13092
rect 27359 13088 27679 14112
rect 27359 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27679 13088
rect 23979 12340 24045 12341
rect 23979 12276 23980 12340
rect 24044 12276 24045 12340
rect 23979 12275 24045 12276
rect 23506 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23826 11456
rect 23506 10368 23826 11392
rect 23506 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23826 10368
rect 23506 9280 23826 10304
rect 23506 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23826 9280
rect 20667 8396 20733 8397
rect 20667 8332 20668 8396
rect 20732 8332 20733 8396
rect 20667 8331 20733 8332
rect 19654 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19974 7648
rect 19654 6560 19974 7584
rect 19654 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19974 6560
rect 19654 5472 19974 6496
rect 19654 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19974 5472
rect 19654 4384 19974 5408
rect 20670 4589 20730 8331
rect 23506 8192 23826 9216
rect 23506 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23826 8192
rect 23506 7104 23826 8128
rect 23506 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23826 7104
rect 23506 6016 23826 7040
rect 23506 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23826 6016
rect 23506 4928 23826 5952
rect 23506 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23826 4928
rect 20667 4588 20733 4589
rect 20667 4524 20668 4588
rect 20732 4524 20733 4588
rect 20667 4523 20733 4524
rect 19654 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19974 4384
rect 19654 3296 19974 4320
rect 19654 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19974 3296
rect 19654 2208 19974 3232
rect 19654 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19974 2208
rect 19654 1120 19974 2144
rect 19654 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19974 1120
rect 19654 496 19974 1056
rect 23506 3840 23826 4864
rect 23506 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23826 3840
rect 23506 2752 23826 3776
rect 23506 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23826 2752
rect 23506 1664 23826 2688
rect 23506 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23826 1664
rect 23506 576 23826 1600
rect 23506 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23826 576
rect 23506 496 23826 512
rect 27359 12000 27679 13024
rect 27359 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27679 12000
rect 27359 10912 27679 11936
rect 27359 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27679 10912
rect 27359 9824 27679 10848
rect 27359 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27679 9824
rect 27359 8736 27679 9760
rect 27359 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27679 8736
rect 27359 7648 27679 8672
rect 27359 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27679 7648
rect 27359 6560 27679 7584
rect 27359 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27679 6560
rect 27359 5472 27679 6496
rect 27359 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27679 5472
rect 27359 4384 27679 5408
rect 27359 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27679 4384
rect 27359 3296 27679 4320
rect 27359 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27679 3296
rect 27359 2208 27679 3232
rect 27359 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27679 2208
rect 27359 1120 27679 2144
rect 27359 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27679 1120
rect 27359 496 27679 1056
rect 31211 19072 31531 19088
rect 31211 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31531 19072
rect 31211 17984 31531 19008
rect 31211 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31531 17984
rect 31211 16896 31531 17920
rect 31211 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31531 16896
rect 31211 15808 31531 16832
rect 31211 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31531 15808
rect 31211 14720 31531 15744
rect 31211 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31531 14720
rect 31211 13632 31531 14656
rect 31211 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31531 13632
rect 31211 12544 31531 13568
rect 31211 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31531 12544
rect 31211 11456 31531 12480
rect 31211 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31531 11456
rect 31211 10368 31531 11392
rect 31211 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31531 10368
rect 31211 9280 31531 10304
rect 31211 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31531 9280
rect 31211 8192 31531 9216
rect 31211 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31531 8192
rect 31211 7104 31531 8128
rect 31211 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31531 7104
rect 31211 6016 31531 7040
rect 31211 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31531 6016
rect 31211 4928 31531 5952
rect 31211 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31531 4928
rect 31211 3840 31531 4864
rect 31211 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31531 3840
rect 31211 2752 31531 3776
rect 31211 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31531 2752
rect 31211 1664 31531 2688
rect 31211 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31531 1664
rect 31211 576 31531 1600
rect 31211 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31531 576
rect 31211 496 31531 512
rect 15147 372 15213 373
rect 15147 308 15148 372
rect 15212 308 15213 372
rect 15147 307 15213 308
use sky130_fd_sc_hd__inv_2  _026__9 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__10
timestamp 1701704242
transform 1 0 24656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__11
timestamp 1701704242
transform 1 0 19136 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__12
timestamp 1701704242
transform 1 0 19228 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__13
timestamp 1701704242
transform 1 0 7176 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__14
timestamp 1701704242
transform -1 0 10028 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__15
timestamp 1701704242
transform 1 0 7452 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__16
timestamp 1701704242
transform 1 0 19044 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__17
timestamp 1701704242
transform -1 0 7268 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__18
timestamp 1701704242
transform -1 0 7176 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__19
timestamp 1701704242
transform -1 0 9752 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__20
timestamp 1701704242
transform 1 0 8648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__21
timestamp 1701704242
transform -1 0 11868 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__22
timestamp 1701704242
transform -1 0 13064 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__23
timestamp 1701704242
transform -1 0 14536 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__24
timestamp 1701704242
transform -1 0 15456 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__25
timestamp 1701704242
transform 1 0 15180 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__26
timestamp 1701704242
transform 1 0 17204 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__27
timestamp 1701704242
transform -1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__28
timestamp 1701704242
transform -1 0 16652 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__29
timestamp 1701704242
transform 1 0 14168 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__30
timestamp 1701704242
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__31
timestamp 1701704242
transform -1 0 15548 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__32
timestamp 1701704242
transform -1 0 12880 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__33
timestamp 1701704242
transform -1 0 11500 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__34
timestamp 1701704242
transform -1 0 11224 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__35
timestamp 1701704242
transform -1 0 8924 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__36
timestamp 1701704242
transform -1 0 8648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__37
timestamp 1701704242
transform -1 0 10304 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__38
timestamp 1701704242
transform 1 0 16192 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__39
timestamp 1701704242
transform -1 0 7176 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__40
timestamp 1701704242
transform -1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__41
timestamp 1701704242
transform -1 0 12052 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__42
timestamp 1701704242
transform 1 0 12696 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__43
timestamp 1701704242
transform 1 0 12512 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__44
timestamp 1701704242
transform -1 0 15640 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__45
timestamp 1701704242
transform 1 0 16284 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__46
timestamp 1701704242
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__47
timestamp 1701704242
transform -1 0 19964 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__48
timestamp 1701704242
transform -1 0 19688 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__49
timestamp 1701704242
transform 1 0 13984 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__50
timestamp 1701704242
transform 1 0 19320 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__51
timestamp 1701704242
transform 1 0 20700 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__52
timestamp 1701704242
transform 1 0 21528 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__53
timestamp 1701704242
transform -1 0 25208 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__54
timestamp 1701704242
transform 1 0 21436 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__55
timestamp 1701704242
transform 1 0 20792 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__56
timestamp 1701704242
transform 1 0 25852 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__57
timestamp 1701704242
transform 1 0 21252 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026__58
timestamp 1701704242
transform -1 0 25760 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _027_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _028_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 7820 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _029_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8924 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _030_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 9384 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _031_
timestamp 1701704242
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp 1701704242
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _033_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14168 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _034_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 14352 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _035_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16376 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _036_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15640 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _037_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16928 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1701704242
transform -1 0 15640 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _039_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 14904 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _040_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13524 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _041_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12696 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1701704242
transform 1 0 13432 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _043_
timestamp 1701704242
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _044_
timestamp 1701704242
transform -1 0 11316 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _045_
timestamp 1701704242
transform -1 0 10304 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _046_
timestamp 1701704242
transform 1 0 10120 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _047_
timestamp 1701704242
transform -1 0 10120 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1701704242
transform 1 0 8740 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _049_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10580 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _050_
timestamp 1701704242
transform 1 0 9476 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _051_
timestamp 1701704242
transform -1 0 10580 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _052_
timestamp 1701704242
transform -1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _053_
timestamp 1701704242
transform 1 0 10028 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _054_
timestamp 1701704242
transform -1 0 9752 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _055_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15640 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _056_
timestamp 1701704242
transform 1 0 13892 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _057_
timestamp 1701704242
transform 1 0 16100 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _058_
timestamp 1701704242
transform 1 0 12972 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _059_
timestamp 1701704242
transform 1 0 11592 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _060_
timestamp 1701704242
transform 1 0 8372 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _061_
timestamp 1701704242
transform 1 0 8372 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _062_
timestamp 1701704242
transform 1 0 9384 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _063_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12420 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _064_
timestamp 1701704242
transform 1 0 13248 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _065_
timestamp 1701704242
transform 1 0 14168 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _066_
timestamp 1701704242
transform 1 0 14536 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _067_
timestamp 1701704242
transform 1 0 16744 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _068_
timestamp 1701704242
transform 1 0 17020 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _069_
timestamp 1701704242
transform 1 0 16100 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _070_
timestamp 1701704242
transform 1 0 17664 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _071_
timestamp 1701704242
transform 1 0 19504 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _072_
timestamp 1701704242
transform 1 0 21252 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _073_
timestamp 1701704242
transform 1 0 21896 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _074_
timestamp 1701704242
transform 1 0 23092 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _075_
timestamp 1701704242
transform 1 0 21436 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _076_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18492 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _077_
timestamp 1701704242
transform 1 0 24196 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _078_
timestamp 1701704242
transform 1 0 21988 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _079_
timestamp 1701704242
transform 1 0 22448 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _080_
timestamp 1701704242
transform 1 0 22172 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _081_
timestamp 1701704242
transform 1 0 18768 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _082_
timestamp 1701704242
transform 1 0 21620 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _083_
timestamp 1701704242
transform 1 0 18676 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _084_
timestamp 1701704242
transform 1 0 22172 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _085_
timestamp 1701704242
transform 1 0 18676 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _086_
timestamp 1701704242
transform 1 0 23092 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _087_
timestamp 1701704242
transform 1 0 22172 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _088_
timestamp 1701704242
transform 1 0 23736 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _089_
timestamp 1701704242
transform 1 0 22172 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _090_
timestamp 1701704242
transform 1 0 22356 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _091_
timestamp 1701704242
transform 1 0 21804 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _092_
timestamp 1701704242
transform -1 0 21804 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _093_
timestamp 1701704242
transform 1 0 18676 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _094_
timestamp 1701704242
transform 1 0 19228 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _095_
timestamp 1701704242
transform 1 0 16744 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _096_
timestamp 1701704242
transform 1 0 17664 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _097_
timestamp 1701704242
transform 1 0 15180 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _098_
timestamp 1701704242
transform -1 0 15272 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _099_
timestamp 1701704242
transform 1 0 14352 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _100_
timestamp 1701704242
transform -1 0 15088 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _101_
timestamp 1701704242
transform 1 0 10856 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _102_
timestamp 1701704242
transform 1 0 9200 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _103_
timestamp 1701704242
transform 1 0 8648 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _104_
timestamp 1701704242
transform 1 0 11960 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _105_
timestamp 1701704242
transform -1 0 10396 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _106_
timestamp 1701704242
transform 1 0 10028 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _107_
timestamp 1701704242
transform -1 0 13156 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _108_
timestamp 1701704242
transform 1 0 13616 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _109_
timestamp 1701704242
transform 1 0 13156 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _110_
timestamp 1701704242
transform 1 0 16100 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _111_
timestamp 1701704242
transform 1 0 17020 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _112_
timestamp 1701704242
transform 1 0 16836 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _113_
timestamp 1701704242
transform 1 0 17020 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _114_
timestamp 1701704242
transform 1 0 17204 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _115_
timestamp 1701704242
transform 1 0 18676 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _116_
timestamp 1701704242
transform 1 0 16100 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _117_
timestamp 1701704242
transform 1 0 13340 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _118_
timestamp 1701704242
transform 1 0 13892 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _119_
timestamp 1701704242
transform 1 0 11868 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _120_
timestamp 1701704242
transform -1 0 11868 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _121_
timestamp 1701704242
transform -1 0 10580 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _122_
timestamp 1701704242
transform -1 0 10120 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _123_
timestamp 1701704242
transform 1 0 11592 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _124_
timestamp 1701704242
transform -1 0 10304 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _125_
timestamp 1701704242
transform -1 0 13248 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _126_
timestamp 1701704242
transform 1 0 11040 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _127_
timestamp 1701704242
transform 1 0 16928 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _128_
timestamp 1701704242
transform 1 0 16928 0 -1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _129_
timestamp 1701704242
transform 1 0 17020 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _130_
timestamp 1701704242
transform 1 0 14444 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _131_
timestamp 1701704242
transform -1 0 14076 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _132_
timestamp 1701704242
transform -1 0 12512 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _133_
timestamp 1701704242
transform 1 0 10856 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _134_
timestamp 1701704242
transform -1 0 12880 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_i_stop pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16008 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net9
timestamp 1701704242
transform 1 0 16100 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_i_stop
timestamp 1701704242
transform -1 0 12788 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_net9
timestamp 1701704242
transform -1 0 12788 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_i_stop
timestamp 1701704242
transform -1 0 15732 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_net9
timestamp 1701704242
transform -1 0 17940 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_i_stop
timestamp 1701704242
transform -1 0 12788 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_net9
timestamp 1701704242
transform -1 0 13064 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_i_stop
timestamp 1701704242
transform -1 0 16008 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_net9
timestamp 1701704242
transform 1 0 15180 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_i_stop
timestamp 1701704242
transform 1 0 16928 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_net9
timestamp 1701704242
transform -1 0 20148 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_i_stop
timestamp 1701704242
transform 1 0 21252 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_net9
timestamp 1701704242
transform 1 0 22356 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_i_stop
timestamp 1701704242
transform 1 0 17572 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_net9
timestamp 1701704242
transform 1 0 18676 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_i_stop
timestamp 1701704242
transform 1 0 21252 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_net9
timestamp 1701704242
transform 1 0 21896 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__nor2_1  dly_stg1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg2
timestamp 1701704242
transform -1 0 9844 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  dly_stg5 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7728 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg6_774
timestamp 1701704242
transform -1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg9_316
timestamp 1701704242
transform -1 0 10672 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg9_317
timestamp 1701704242
transform -1 0 9384 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg9_318
timestamp 1701704242
transform 1 0 10580 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_466
timestamp 1701704242
transform 1 0 11592 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_467
timestamp 1701704242
transform 1 0 9292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_468
timestamp 1701704242
transform -1 0 11408 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_469
timestamp 1701704242
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_470
timestamp 1701704242
transform -1 0 10856 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_471
timestamp 1701704242
transform -1 0 8464 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_472
timestamp 1701704242
transform 1 0 9200 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_473
timestamp 1701704242
transform -1 0 12972 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_474
timestamp 1701704242
transform 1 0 13064 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_475
timestamp 1701704242
transform 1 0 16468 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_476
timestamp 1701704242
transform -1 0 15088 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_477
timestamp 1701704242
transform 1 0 16376 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_478
timestamp 1701704242
transform 1 0 8464 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg11_629
timestamp 1701704242
transform 1 0 10580 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg11_630
timestamp 1701704242
transform -1 0 10580 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg11_631
timestamp 1701704242
transform 1 0 11408 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_319
timestamp 1701704242
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_320
timestamp 1701704242
transform -1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_321
timestamp 1701704242
transform -1 0 11316 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_322
timestamp 1701704242
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  fanout1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10396 0 1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1701704242
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1701704242
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6900 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_77 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7636 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1701704242
transform 1 0 8096 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1701704242
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1701704242
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1701704242
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1701704242
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1701704242
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1701704242
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1701704242
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1701704242
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1701704242
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1701704242
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1701704242
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1701704242
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1701704242
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1701704242
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1701704242
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1701704242
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1701704242
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1701704242
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1701704242
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1701704242
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1701704242
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1701704242
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1701704242
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1701704242
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_321
timestamp 1701704242
transform 1 0 30084 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_329
timestamp 1701704242
transform 1 0 30820 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1701704242
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1701704242
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1701704242
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1701704242
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1701704242
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1701704242
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1701704242
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1701704242
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1701704242
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1701704242
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1701704242
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1701704242
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1701704242
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1701704242
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1701704242
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1701704242
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1701704242
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1701704242
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1701704242
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1701704242
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1701704242
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1701704242
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1701704242
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1701704242
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1701704242
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1701704242
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1701704242
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1701704242
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_329
timestamp 1701704242
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1701704242
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1701704242
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1701704242
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1701704242
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1701704242
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1701704242
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1701704242
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1701704242
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1701704242
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1701704242
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1701704242
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1701704242
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1701704242
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1701704242
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1701704242
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1701704242
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1701704242
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1701704242
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1701704242
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1701704242
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1701704242
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1701704242
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1701704242
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1701704242
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1701704242
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1701704242
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1701704242
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1701704242
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1701704242
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1701704242
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1701704242
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1701704242
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1701704242
transform 1 0 30084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_329
timestamp 1701704242
transform 1 0 30820 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1701704242
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1701704242
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1701704242
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1701704242
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1701704242
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1701704242
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1701704242
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1701704242
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1701704242
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1701704242
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1701704242
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1701704242
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1701704242
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1701704242
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1701704242
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1701704242
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1701704242
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1701704242
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1701704242
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1701704242
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1701704242
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1701704242
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1701704242
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1701704242
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1701704242
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1701704242
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1701704242
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1701704242
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1701704242
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1701704242
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1701704242
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_329
timestamp 1701704242
transform 1 0 30820 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1701704242
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1701704242
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1701704242
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1701704242
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1701704242
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1701704242
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1701704242
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1701704242
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1701704242
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1701704242
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1701704242
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1701704242
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1701704242
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1701704242
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1701704242
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1701704242
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1701704242
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1701704242
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1701704242
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1701704242
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1701704242
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1701704242
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1701704242
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1701704242
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1701704242
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1701704242
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1701704242
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1701704242
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1701704242
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_321
timestamp 1701704242
transform 1 0 30084 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_329
timestamp 1701704242
transform 1 0 30820 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1701704242
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1701704242
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1701704242
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1701704242
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1701704242
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1701704242
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_81
timestamp 1701704242
transform 1 0 8004 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_106
timestamp 1701704242
transform 1 0 10304 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_147
timestamp 1701704242
transform 1 0 14076 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_152
timestamp 1701704242
transform 1 0 14536 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_158
timestamp 1701704242
transform 1 0 15088 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_175
timestamp 1701704242
transform 1 0 16652 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_195
timestamp 1701704242
transform 1 0 18492 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_207
timestamp 1701704242
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_219
timestamp 1701704242
transform 1 0 20700 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1701704242
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1701704242
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1701704242
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1701704242
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1701704242
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1701704242
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1701704242
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1701704242
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1701704242
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1701704242
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1701704242
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_329
timestamp 1701704242
transform 1 0 30820 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1701704242
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1701704242
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1701704242
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1701704242
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1701704242
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1701704242
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1701704242
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_92
timestamp 1701704242
transform 1 0 9016 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_96
timestamp 1701704242
transform 1 0 9384 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_110
timestamp 1701704242
transform 1 0 10672 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_117
timestamp 1701704242
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_136
timestamp 1701704242
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_141
timestamp 1701704242
transform 1 0 13524 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_161
timestamp 1701704242
transform 1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_180
timestamp 1701704242
transform 1 0 17112 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_192
timestamp 1701704242
transform 1 0 18216 0 1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1701704242
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1701704242
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1701704242
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1701704242
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1701704242
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1701704242
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1701704242
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1701704242
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1701704242
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1701704242
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1701704242
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1701704242
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1701704242
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_321
timestamp 1701704242
transform 1 0 30084 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_329
timestamp 1701704242
transform 1 0 30820 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1701704242
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1701704242
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1701704242
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1701704242
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1701704242
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1701704242
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1701704242
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1701704242
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_93
timestamp 1701704242
transform 1 0 9108 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1701704242
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_124
timestamp 1701704242
transform 1 0 11960 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_129
timestamp 1701704242
transform 1 0 12420 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_135
timestamp 1701704242
transform 1 0 12972 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_139
timestamp 1701704242
transform 1 0 13340 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_143
timestamp 1701704242
transform 1 0 13708 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_150
timestamp 1701704242
transform 1 0 14352 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_156
timestamp 1701704242
transform 1 0 14904 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_160
timestamp 1701704242
transform 1 0 15272 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_172
timestamp 1701704242
transform 1 0 16376 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_176
timestamp 1701704242
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_195
timestamp 1701704242
transform 1 0 18492 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_207
timestamp 1701704242
transform 1 0 19596 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_213
timestamp 1701704242
transform 1 0 20148 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1701704242
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1701704242
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1701704242
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1701704242
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1701704242
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1701704242
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1701704242
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1701704242
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1701704242
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1701704242
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1701704242
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_329
timestamp 1701704242
transform 1 0 30820 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1701704242
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1701704242
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1701704242
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1701704242
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1701704242
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_77
timestamp 1701704242
transform 1 0 7636 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_101
timestamp 1701704242
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1701704242
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_162
timestamp 1701704242
transform 1 0 15456 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_172
timestamp 1701704242
transform 1 0 16376 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_178
timestamp 1701704242
transform 1 0 16928 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_200
timestamp 1701704242
transform 1 0 18952 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_238
timestamp 1701704242
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_250
timestamp 1701704242
transform 1 0 23552 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1701704242
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1701704242
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1701704242
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1701704242
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1701704242
transform 1 0 28244 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1701704242
transform 1 0 28796 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1701704242
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_321
timestamp 1701704242
transform 1 0 30084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_329
timestamp 1701704242
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1701704242
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1701704242
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1701704242
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1701704242
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1701704242
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1701704242
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1701704242
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_69
timestamp 1701704242
transform 1 0 6900 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1701704242
transform 1 0 10948 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_134
timestamp 1701704242
transform 1 0 12880 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_185
timestamp 1701704242
transform 1 0 17572 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1701704242
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1701704242
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1701704242
transform 1 0 25668 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1701704242
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1701704242
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1701704242
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1701704242
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1701704242
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_329
timestamp 1701704242
transform 1 0 30820 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1701704242
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1701704242
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1701704242
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1701704242
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1701704242
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_65
timestamp 1701704242
transform 1 0 6532 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_71
timestamp 1701704242
transform 1 0 7084 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_100
timestamp 1701704242
transform 1 0 9752 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_110
timestamp 1701704242
transform 1 0 10672 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1701704242
transform 1 0 13524 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_165
timestamp 1701704242
transform 1 0 15732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1701704242
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1701704242
transform 1 0 23552 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_259
timestamp 1701704242
transform 1 0 24380 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_271
timestamp 1701704242
transform 1 0 25484 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_283
timestamp 1701704242
transform 1 0 26588 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_295
timestamp 1701704242
transform 1 0 27692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1701704242
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1701704242
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_321
timestamp 1701704242
transform 1 0 30084 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_329
timestamp 1701704242
transform 1 0 30820 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1701704242
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1701704242
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1701704242
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1701704242
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1701704242
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_91
timestamp 1701704242
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_105
timestamp 1701704242
transform 1 0 10212 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1701704242
transform 1 0 10948 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_146
timestamp 1701704242
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 1701704242
transform 1 0 16100 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_176
timestamp 1701704242
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1701704242
transform 1 0 20976 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_266
timestamp 1701704242
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 1701704242
transform 1 0 26128 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1701704242
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1701704242
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1701704242
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1701704242
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_329
timestamp 1701704242
transform 1 0 30820 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1701704242
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1701704242
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1701704242
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_53
timestamp 1701704242
transform 1 0 5428 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_59
timestamp 1701704242
transform 1 0 5980 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1701704242
transform 1 0 8372 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_107
timestamp 1701704242
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1701704242
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1701704242
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_230
timestamp 1701704242
transform 1 0 21712 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_274
timestamp 1701704242
transform 1 0 25760 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_286
timestamp 1701704242
transform 1 0 26864 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_298
timestamp 1701704242
transform 1 0 27968 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_306
timestamp 1701704242
transform 1 0 28704 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1701704242
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_321
timestamp 1701704242
transform 1 0 30084 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_329
timestamp 1701704242
transform 1 0 30820 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1701704242
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1701704242
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1701704242
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1701704242
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1701704242
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1701704242
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1701704242
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_69
timestamp 1701704242
transform 1 0 6900 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_133
timestamp 1701704242
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_155
timestamp 1701704242
transform 1 0 14812 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_169
timestamp 1701704242
transform 1 0 16100 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_219
timestamp 1701704242
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1701704242
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1701704242
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1701704242
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1701704242
transform 1 0 28612 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1701704242
transform 1 0 29716 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_329
timestamp 1701704242
transform 1 0 30820 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1701704242
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1701704242
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1701704242
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1701704242
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_65
timestamp 1701704242
transform 1 0 6532 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1701704242
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_106
timestamp 1701704242
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1701704242
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1701704242
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1701704242
transform 1 0 23552 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_286
timestamp 1701704242
transform 1 0 26864 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_298
timestamp 1701704242
transform 1 0 27968 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_306
timestamp 1701704242
transform 1 0 28704 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1701704242
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_321
timestamp 1701704242
transform 1 0 30084 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_329
timestamp 1701704242
transform 1 0 30820 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1701704242
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1701704242
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1701704242
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1701704242
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1701704242
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_57
timestamp 1701704242
transform 1 0 5796 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_63
timestamp 1701704242
transform 1 0 6348 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_220
timestamp 1701704242
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_284
timestamp 1701704242
transform 1 0 26680 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_296
timestamp 1701704242
transform 1 0 27784 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_308
timestamp 1701704242
transform 1 0 28888 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_320
timestamp 1701704242
transform 1 0 29992 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1701704242
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1701704242
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1701704242
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_53
timestamp 1701704242
transform 1 0 5428 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_59
timestamp 1701704242
transform 1 0 5980 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1701704242
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1701704242
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_223
timestamp 1701704242
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1701704242
transform 1 0 23552 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1701704242
transform 1 0 27140 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1701704242
transform 1 0 28244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1701704242
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1701704242
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_321
timestamp 1701704242
transform 1 0 30084 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_329
timestamp 1701704242
transform 1 0 30820 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1701704242
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1701704242
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1701704242
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1701704242
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1701704242
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_57
timestamp 1701704242
transform 1 0 5796 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_65
timestamp 1701704242
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_113
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_215
timestamp 1701704242
transform 1 0 20332 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1701704242
transform 1 0 21068 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_225
timestamp 1701704242
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1701704242
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1701704242
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1701704242
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1701704242
transform 1 0 28612 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1701704242
transform 1 0 29716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_329
timestamp 1701704242
transform 1 0 30820 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1701704242
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1701704242
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1701704242
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1701704242
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1701704242
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_65
timestamp 1701704242
transform 1 0 6532 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_73
timestamp 1701704242
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1701704242
transform 1 0 13524 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_162
timestamp 1701704242
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_212
timestamp 1701704242
transform 1 0 20056 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_234
timestamp 1701704242
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_274
timestamp 1701704242
transform 1 0 25760 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_286
timestamp 1701704242
transform 1 0 26864 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_298
timestamp 1701704242
transform 1 0 27968 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_306
timestamp 1701704242
transform 1 0 28704 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1701704242
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_321
timestamp 1701704242
transform 1 0 30084 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_329
timestamp 1701704242
transform 1 0 30820 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1701704242
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1701704242
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1701704242
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1701704242
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1701704242
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1701704242
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_81
timestamp 1701704242
transform 1 0 8004 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_154
timestamp 1701704242
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_210
timestamp 1701704242
transform 1 0 19872 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_220
timestamp 1701704242
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_228
timestamp 1701704242
transform 1 0 21528 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_272
timestamp 1701704242
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1701704242
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1701704242
transform 1 0 27508 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1701704242
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1701704242
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_329
timestamp 1701704242
transform 1 0 30820 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1701704242
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1701704242
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1701704242
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1701704242
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1701704242
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1701704242
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_65
timestamp 1701704242
transform 1 0 6532 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_73
timestamp 1701704242
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1701704242
transform 1 0 13524 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_169
timestamp 1701704242
transform 1 0 16100 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_176
timestamp 1701704242
transform 1 0 16744 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_234
timestamp 1701704242
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_280
timestamp 1701704242
transform 1 0 26312 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_292
timestamp 1701704242
transform 1 0 27416 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_304
timestamp 1701704242
transform 1 0 28520 0 1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1701704242
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_321
timestamp 1701704242
transform 1 0 30084 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_329
timestamp 1701704242
transform 1 0 30820 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1701704242
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1701704242
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1701704242
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1701704242
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1701704242
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1701704242
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1701704242
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_69
timestamp 1701704242
transform 1 0 6900 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_77
timestamp 1701704242
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_113
timestamp 1701704242
transform 1 0 10948 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_184
timestamp 1701704242
transform 1 0 17480 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_214
timestamp 1701704242
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1701704242
transform 1 0 20976 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1701704242
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1701704242
transform 1 0 27508 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1701704242
transform 1 0 28612 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1701704242
transform 1 0 29716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_329
timestamp 1701704242
transform 1 0 30820 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1701704242
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1701704242
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1701704242
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1701704242
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1701704242
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1701704242
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_65
timestamp 1701704242
transform 1 0 6532 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_73
timestamp 1701704242
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1701704242
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_133
timestamp 1701704242
transform 1 0 12788 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 1701704242
transform 1 0 13524 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_286
timestamp 1701704242
transform 1 0 26864 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_298
timestamp 1701704242
transform 1 0 27968 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_306
timestamp 1701704242
transform 1 0 28704 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1701704242
transform 1 0 28980 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_321
timestamp 1701704242
transform 1 0 30084 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_329
timestamp 1701704242
transform 1 0 30820 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1701704242
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1701704242
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1701704242
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1701704242
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1701704242
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1701704242
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1701704242
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_69
timestamp 1701704242
transform 1 0 6900 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_113
timestamp 1701704242
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_141
timestamp 1701704242
transform 1 0 13524 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1701704242
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_225
timestamp 1701704242
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_278
timestamp 1701704242
transform 1 0 26128 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_284
timestamp 1701704242
transform 1 0 26680 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_296
timestamp 1701704242
transform 1 0 27784 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_308
timestamp 1701704242
transform 1 0 28888 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_320
timestamp 1701704242
transform 1 0 29992 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1701704242
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1701704242
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1701704242
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1701704242
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1701704242
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1701704242
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_65
timestamp 1701704242
transform 1 0 6532 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_105
timestamp 1701704242
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 1701704242
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_163
timestamp 1701704242
transform 1 0 15548 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_176
timestamp 1701704242
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_286
timestamp 1701704242
transform 1 0 26864 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_298
timestamp 1701704242
transform 1 0 27968 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1701704242
transform 1 0 28704 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1701704242
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_321
timestamp 1701704242
transform 1 0 30084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_329
timestamp 1701704242
transform 1 0 30820 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1701704242
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1701704242
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1701704242
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1701704242
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1701704242
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1701704242
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1701704242
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_69
timestamp 1701704242
transform 1 0 6900 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1701704242
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_136
timestamp 1701704242
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1701704242
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1701704242
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_278
timestamp 1701704242
transform 1 0 26128 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1701704242
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1701704242
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1701704242
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1701704242
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_329
timestamp 1701704242
transform 1 0 30820 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1701704242
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1701704242
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1701704242
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1701704242
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1701704242
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1701704242
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1701704242
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_77
timestamp 1701704242
transform 1 0 7636 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_129
timestamp 1701704242
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1701704242
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_158
timestamp 1701704242
transform 1 0 15088 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1701704242
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_274
timestamp 1701704242
transform 1 0 25760 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_286
timestamp 1701704242
transform 1 0 26864 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_298
timestamp 1701704242
transform 1 0 27968 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_306
timestamp 1701704242
transform 1 0 28704 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1701704242
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1701704242
transform 1 0 30084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_329
timestamp 1701704242
transform 1 0 30820 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1701704242
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1701704242
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1701704242
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1701704242
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1701704242
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1701704242
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1701704242
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1701704242
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_81
timestamp 1701704242
transform 1 0 8004 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_87
timestamp 1701704242
transform 1 0 8556 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_113
timestamp 1701704242
transform 1 0 10948 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_135
timestamp 1701704242
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_155
timestamp 1701704242
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1701704242
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1701704242
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_267
timestamp 1701704242
transform 1 0 25116 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1701704242
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1701704242
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1701704242
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1701704242
transform 1 0 28612 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1701704242
transform 1 0 29716 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_329
timestamp 1701704242
transform 1 0 30820 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1701704242
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1701704242
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1701704242
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1701704242
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1701704242
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1701704242
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1701704242
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1701704242
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1701704242
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1701704242
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_130
timestamp 1701704242
transform 1 0 12512 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1701704242
transform 1 0 13524 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_160
timestamp 1701704242
transform 1 0 15272 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_164
timestamp 1701704242
transform 1 0 15640 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_177
timestamp 1701704242
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_185
timestamp 1701704242
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_189
timestamp 1701704242
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1701704242
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_262
timestamp 1701704242
transform 1 0 24656 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_274
timestamp 1701704242
transform 1 0 25760 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_286
timestamp 1701704242
transform 1 0 26864 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_298
timestamp 1701704242
transform 1 0 27968 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_306
timestamp 1701704242
transform 1 0 28704 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1701704242
transform 1 0 28980 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_321
timestamp 1701704242
transform 1 0 30084 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_329
timestamp 1701704242
transform 1 0 30820 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1701704242
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1701704242
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1701704242
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1701704242
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1701704242
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1701704242
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1701704242
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1701704242
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1701704242
transform 1 0 8004 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_93
timestamp 1701704242
transform 1 0 9108 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_101
timestamp 1701704242
transform 1 0 9844 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_105
timestamp 1701704242
transform 1 0 10212 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_131
timestamp 1701704242
transform 1 0 12604 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_141
timestamp 1701704242
transform 1 0 13524 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_152
timestamp 1701704242
transform 1 0 14536 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_172
timestamp 1701704242
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_184
timestamp 1701704242
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_196
timestamp 1701704242
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_213
timestamp 1701704242
transform 1 0 20148 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1701704242
transform 1 0 21068 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_252
timestamp 1701704242
transform 1 0 23736 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_264
timestamp 1701704242
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_276
timestamp 1701704242
transform 1 0 25944 0 -1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1701704242
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1701704242
transform 1 0 27508 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1701704242
transform 1 0 28612 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1701704242
transform 1 0 29716 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_329
timestamp 1701704242
transform 1 0 30820 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1701704242
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1701704242
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1701704242
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1701704242
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1701704242
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1701704242
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1701704242
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1701704242
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1701704242
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1701704242
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_109
timestamp 1701704242
transform 1 0 10580 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_128
timestamp 1701704242
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_138
timestamp 1701704242
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_147
timestamp 1701704242
transform 1 0 14076 0 1 16864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_158
timestamp 1701704242
transform 1 0 15088 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_170
timestamp 1701704242
transform 1 0 16192 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_182
timestamp 1701704242
transform 1 0 17296 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1701704242
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1701704242
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_209
timestamp 1701704242
transform 1 0 19780 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_246
timestamp 1701704242
transform 1 0 23184 0 1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1701704242
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1701704242
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1701704242
transform 1 0 26036 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1701704242
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1701704242
transform 1 0 28244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1701704242
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1701704242
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_321
timestamp 1701704242
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_329
timestamp 1701704242
transform 1 0 30820 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1701704242
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1701704242
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1701704242
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1701704242
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1701704242
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1701704242
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1701704242
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1701704242
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1701704242
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1701704242
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1701704242
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1701704242
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1701704242
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1701704242
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1701704242
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1701704242
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1701704242
transform 1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1701704242
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1701704242
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1701704242
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1701704242
transform 1 0 18308 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1701704242
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_217
timestamp 1701704242
transform 1 0 20516 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_221
timestamp 1701704242
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1701704242
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1701704242
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1701704242
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1701704242
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1701704242
transform 1 0 25668 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1701704242
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1701704242
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1701704242
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1701704242
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1701704242
transform 1 0 29716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_329
timestamp 1701704242
transform 1 0 30820 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1701704242
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1701704242
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1701704242
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1701704242
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1701704242
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1701704242
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1701704242
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1701704242
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1701704242
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1701704242
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1701704242
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1701704242
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1701704242
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1701704242
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1701704242
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1701704242
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1701704242
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1701704242
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1701704242
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1701704242
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1701704242
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1701704242
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1701704242
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1701704242
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1701704242
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1701704242
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1701704242
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1701704242
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1701704242
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1701704242
transform 1 0 26036 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1701704242
transform 1 0 27140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1701704242
transform 1 0 28244 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1701704242
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1701704242
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1701704242
transform 1 0 30084 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_329
timestamp 1701704242
transform 1 0 30820 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1701704242
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1701704242
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_27
timestamp 1701704242
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1701704242
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1701704242
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1701704242
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1701704242
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1701704242
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1701704242
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_85
timestamp 1701704242
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1701704242
transform 1 0 9476 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1701704242
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1701704242
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1701704242
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_137
timestamp 1701704242
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_141
timestamp 1701704242
transform 1 0 13524 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_153
timestamp 1701704242
transform 1 0 14628 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1701704242
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1701704242
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1701704242
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_193
timestamp 1701704242
transform 1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_197
timestamp 1701704242
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_209
timestamp 1701704242
transform 1 0 19780 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1701704242
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1701704242
transform 1 0 21252 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1701704242
transform 1 0 22356 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_249
timestamp 1701704242
transform 1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1701704242
transform 1 0 23828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_265
timestamp 1701704242
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1701704242
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1701704242
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1701704242
transform 1 0 27508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_305
timestamp 1701704242
transform 1 0 28612 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_309
timestamp 1701704242
transform 1 0 28980 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_321
timestamp 1701704242
transform 1 0 30084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_329
timestamp 1701704242
transform 1 0 30820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[1\].dly_stg3
timestamp 1701704242
transform 1 0 10856 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_72
timestamp 1701704242
transform 1 0 14904 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_73
timestamp 1701704242
transform 1 0 11316 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_74
timestamp 1701704242
transform 1 0 15548 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_75
timestamp 1701704242
transform 1 0 14628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[2\].dly_stg3
timestamp 1701704242
transform -1 0 16376 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_76
timestamp 1701704242
transform -1 0 15088 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_77
timestamp 1701704242
transform -1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_78
timestamp 1701704242
transform -1 0 16744 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_79
timestamp 1701704242
transform -1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[3\].dly_stg3
timestamp 1701704242
transform -1 0 16468 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_80
timestamp 1701704242
transform -1 0 18492 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_81
timestamp 1701704242
transform -1 0 15916 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_82
timestamp 1701704242
transform -1 0 16744 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_83
timestamp 1701704242
transform 1 0 18676 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[4\].dly_stg3
timestamp 1701704242
transform 1 0 14536 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_84
timestamp 1701704242
transform -1 0 20148 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_85
timestamp 1701704242
transform 1 0 19228 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_86
timestamp 1701704242
transform -1 0 18952 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_87
timestamp 1701704242
transform 1 0 19780 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[5\].dly_stg3
timestamp 1701704242
transform 1 0 19320 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_88
timestamp 1701704242
transform 1 0 21436 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_89
timestamp 1701704242
transform 1 0 19504 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_90
timestamp 1701704242
transform 1 0 20884 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_91
timestamp 1701704242
transform 1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[6\].dly_stg3
timestamp 1701704242
transform -1 0 20700 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_92
timestamp 1701704242
transform 1 0 23092 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_93
timestamp 1701704242
transform -1 0 19504 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_94
timestamp 1701704242
transform -1 0 19964 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_95
timestamp 1701704242
transform 1 0 19504 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[7\].dly_stg3
timestamp 1701704242
transform -1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_96
timestamp 1701704242
transform 1 0 24932 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_97
timestamp 1701704242
transform 1 0 22172 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_98
timestamp 1701704242
transform -1 0 20792 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_99
timestamp 1701704242
transform 1 0 22356 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[8\].dly_stg3
timestamp 1701704242
transform 1 0 20792 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_100
timestamp 1701704242
transform -1 0 23460 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_101
timestamp 1701704242
transform -1 0 20608 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_102
timestamp 1701704242
transform -1 0 22172 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_103
timestamp 1701704242
transform -1 0 24380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[9\].dly_stg3
timestamp 1701704242
transform -1 0 23552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_104
timestamp 1701704242
transform -1 0 21344 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_105
timestamp 1701704242
transform 1 0 24380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_106
timestamp 1701704242
transform -1 0 23184 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_107
timestamp 1701704242
transform 1 0 25484 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[10\].dly_stg3
timestamp 1701704242
transform -1 0 24748 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_108
timestamp 1701704242
transform -1 0 22356 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_109
timestamp 1701704242
transform 1 0 23644 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_110
timestamp 1701704242
transform -1 0 21528 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_111
timestamp 1701704242
transform 1 0 26588 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[11\].dly_stg3
timestamp 1701704242
transform 1 0 23828 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_112
timestamp 1701704242
transform 1 0 21160 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_113
timestamp 1701704242
transform 1 0 26036 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_114
timestamp 1701704242
transform 1 0 20608 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_115
timestamp 1701704242
transform -1 0 24656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[12\].dly_stg3
timestamp 1701704242
transform -1 0 21160 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_116
timestamp 1701704242
transform 1 0 20792 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_117
timestamp 1701704242
transform 1 0 24656 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_118
timestamp 1701704242
transform 1 0 25208 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_119
timestamp 1701704242
transform -1 0 19504 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[13\].dly_stg3
timestamp 1701704242
transform 1 0 25760 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_120
timestamp 1701704242
transform -1 0 25760 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_121
timestamp 1701704242
transform -1 0 23644 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_122
timestamp 1701704242
transform 1 0 24104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_123
timestamp 1701704242
transform -1 0 26680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[14\].dly_stg3
timestamp 1701704242
transform -1 0 23276 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[14\].dly_stg4_124
timestamp 1701704242
transform 1 0 23828 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[14\].dly_stg4_125
timestamp 1701704242
transform -1 0 25484 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[14\].dly_stg4_126
timestamp 1701704242
transform 1 0 25484 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[14\].dly_stg4_127
timestamp 1701704242
transform 1 0 26312 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[15\].dly_stg3
timestamp 1701704242
transform -1 0 25392 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[15\].dly_stg4_128
timestamp 1701704242
transform 1 0 23828 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[15\].dly_stg4_129
timestamp 1701704242
transform 1 0 24380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[15\].dly_stg4_130
timestamp 1701704242
transform 1 0 21252 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[15\].dly_stg4_131
timestamp 1701704242
transform -1 0 25300 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[16\].dly_stg3
timestamp 1701704242
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[16\].dly_stg4_132
timestamp 1701704242
transform -1 0 21528 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[16\].dly_stg4_133
timestamp 1701704242
transform 1 0 23920 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[16\].dly_stg4_134
timestamp 1701704242
transform 1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[16\].dly_stg4_135
timestamp 1701704242
transform -1 0 25208 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[17\].dly_stg3
timestamp 1701704242
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[17\].dly_stg4_136
timestamp 1701704242
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[17\].dly_stg4_137
timestamp 1701704242
transform -1 0 21068 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[17\].dly_stg4_138
timestamp 1701704242
transform 1 0 20700 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[17\].dly_stg4_139
timestamp 1701704242
transform 1 0 19780 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[18\].dly_stg3
timestamp 1701704242
transform 1 0 20424 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[18\].dly_stg4_140
timestamp 1701704242
transform 1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[18\].dly_stg4_141
timestamp 1701704242
transform 1 0 24656 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[18\].dly_stg4_142
timestamp 1701704242
transform -1 0 24656 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[18\].dly_stg4_143
timestamp 1701704242
transform -1 0 25484 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[19\].dly_stg3
timestamp 1701704242
transform 1 0 19964 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[19\].dly_stg4_144
timestamp 1701704242
transform -1 0 22172 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[19\].dly_stg4_145
timestamp 1701704242
transform -1 0 21252 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[19\].dly_stg4_146
timestamp 1701704242
transform -1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[19\].dly_stg4_147
timestamp 1701704242
transform -1 0 19872 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[20\].dly_stg3
timestamp 1701704242
transform 1 0 20700 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[20\].dly_stg4_148
timestamp 1701704242
transform -1 0 26312 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[20\].dly_stg4_149
timestamp 1701704242
transform -1 0 20700 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[20\].dly_stg4_150
timestamp 1701704242
transform -1 0 25208 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[20\].dly_stg4_151
timestamp 1701704242
transform 1 0 26036 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[21\].dly_stg3
timestamp 1701704242
transform 1 0 24656 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[21\].dly_stg4_152
timestamp 1701704242
transform -1 0 24656 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[21\].dly_stg4_153
timestamp 1701704242
transform -1 0 21068 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[21\].dly_stg4_154
timestamp 1701704242
transform -1 0 22080 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[21\].dly_stg4_155
timestamp 1701704242
transform -1 0 20516 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[22\].dly_stg3
timestamp 1701704242
transform -1 0 24932 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[22\].dly_stg4_156
timestamp 1701704242
transform -1 0 24656 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[22\].dly_stg4_157
timestamp 1701704242
transform -1 0 25760 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[22\].dly_stg4_158
timestamp 1701704242
transform 1 0 24196 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[22\].dly_stg4_159
timestamp 1701704242
transform -1 0 26036 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[23\].dly_stg3
timestamp 1701704242
transform 1 0 22356 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[23\].dly_stg4_160
timestamp 1701704242
transform -1 0 24012 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[23\].dly_stg4_161
timestamp 1701704242
transform -1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[23\].dly_stg4_162
timestamp 1701704242
transform 1 0 24932 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[23\].dly_stg4_163
timestamp 1701704242
transform -1 0 26312 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[24\].dly_stg3
timestamp 1701704242
transform -1 0 24380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[24\].dly_stg4_164
timestamp 1701704242
transform 1 0 26312 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[24\].dly_stg4_165
timestamp 1701704242
transform -1 0 25024 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[24\].dly_stg4_166
timestamp 1701704242
transform -1 0 24748 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[24\].dly_stg4_167
timestamp 1701704242
transform 1 0 25852 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[25\].dly_stg3
timestamp 1701704242
transform -1 0 25576 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[25\].dly_stg4_168
timestamp 1701704242
transform -1 0 23092 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[25\].dly_stg4_169
timestamp 1701704242
transform -1 0 23368 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[25\].dly_stg4_170
timestamp 1701704242
transform -1 0 21528 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[25\].dly_stg4_171
timestamp 1701704242
transform 1 0 26588 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[26\].dly_stg3
timestamp 1701704242
transform -1 0 21160 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[26\].dly_stg4_172
timestamp 1701704242
transform -1 0 21804 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[26\].dly_stg4_173
timestamp 1701704242
transform 1 0 25208 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[26\].dly_stg4_174
timestamp 1701704242
transform -1 0 23460 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[26\].dly_stg4_175
timestamp 1701704242
transform -1 0 23736 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[27\].dly_stg3
timestamp 1701704242
transform -1 0 23644 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[27\].dly_stg4_176
timestamp 1701704242
transform 1 0 22632 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[27\].dly_stg4_177
timestamp 1701704242
transform -1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[27\].dly_stg4_178
timestamp 1701704242
transform -1 0 21528 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[27\].dly_stg4_179
timestamp 1701704242
transform -1 0 23184 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[28\].dly_stg3
timestamp 1701704242
transform -1 0 22264 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[28\].dly_stg4_180
timestamp 1701704242
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[28\].dly_stg4_181
timestamp 1701704242
transform -1 0 22080 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[28\].dly_stg4_182
timestamp 1701704242
transform -1 0 20148 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[28\].dly_stg4_183
timestamp 1701704242
transform 1 0 24656 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[29\].dly_stg3
timestamp 1701704242
transform -1 0 20056 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[29\].dly_stg4_184
timestamp 1701704242
transform 1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[29\].dly_stg4_185
timestamp 1701704242
transform -1 0 20424 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[29\].dly_stg4_186
timestamp 1701704242
transform -1 0 19504 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[29\].dly_stg4_187
timestamp 1701704242
transform 1 0 20608 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[30\].dly_stg3
timestamp 1701704242
transform -1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[30\].dly_stg4_188
timestamp 1701704242
transform 1 0 18308 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[30\].dly_stg4_189
timestamp 1701704242
transform -1 0 19780 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[30\].dly_stg4_190
timestamp 1701704242
transform -1 0 18860 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[30\].dly_stg4_191
timestamp 1701704242
transform -1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[31\].dly_stg3
timestamp 1701704242
transform 1 0 19136 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[31\].dly_stg4_192
timestamp 1701704242
transform -1 0 16928 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[31\].dly_stg4_193
timestamp 1701704242
transform -1 0 18308 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[31\].dly_stg4_194
timestamp 1701704242
transform -1 0 17480 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[31\].dly_stg4_195
timestamp 1701704242
transform -1 0 17296 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[32\].dly_stg3
timestamp 1701704242
transform 1 0 17480 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[32\].dly_stg4_196
timestamp 1701704242
transform -1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[32\].dly_stg4_197
timestamp 1701704242
transform 1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[32\].dly_stg4_198
timestamp 1701704242
transform 1 0 16652 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[32\].dly_stg4_199
timestamp 1701704242
transform -1 0 18032 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[33\].dly_stg3
timestamp 1701704242
transform 1 0 15732 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[33\].dly_stg4_200
timestamp 1701704242
transform 1 0 14260 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[33\].dly_stg4_201
timestamp 1701704242
transform -1 0 16376 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[33\].dly_stg4_202
timestamp 1701704242
transform 1 0 15548 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[33\].dly_stg4_203
timestamp 1701704242
transform -1 0 16008 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[34\].dly_stg3
timestamp 1701704242
transform -1 0 15548 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[34\].dly_stg4_204
timestamp 1701704242
transform 1 0 13892 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[34\].dly_stg4_205
timestamp 1701704242
transform 1 0 17204 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[34\].dly_stg4_206
timestamp 1701704242
transform -1 0 13064 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[34\].dly_stg4_207
timestamp 1701704242
transform -1 0 12604 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[35\].dly_stg3
timestamp 1701704242
transform -1 0 13984 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[35\].dly_stg4_208
timestamp 1701704242
transform -1 0 13432 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[35\].dly_stg4_209
timestamp 1701704242
transform 1 0 14720 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[35\].dly_stg4_210
timestamp 1701704242
transform -1 0 11868 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[35\].dly_stg4_211
timestamp 1701704242
transform -1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[36\].dly_stg3
timestamp 1701704242
transform 1 0 12604 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[36\].dly_stg4_212
timestamp 1701704242
transform 1 0 11776 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[36\].dly_stg4_213
timestamp 1701704242
transform -1 0 13156 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[36\].dly_stg4_214
timestamp 1701704242
transform -1 0 10028 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[36\].dly_stg4_215
timestamp 1701704242
transform 1 0 15180 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[37\].dly_stg3
timestamp 1701704242
transform 1 0 10304 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[37\].dly_stg4_216
timestamp 1701704242
transform -1 0 10580 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[37\].dly_stg4_217
timestamp 1701704242
transform -1 0 11316 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[37\].dly_stg4_218
timestamp 1701704242
transform -1 0 11500 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[37\].dly_stg4_219
timestamp 1701704242
transform -1 0 9752 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[38\].dly_stg3
timestamp 1701704242
transform -1 0 8924 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[38\].dly_stg4_220
timestamp 1701704242
transform 1 0 12328 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[38\].dly_stg4_221
timestamp 1701704242
transform 1 0 11224 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[38\].dly_stg4_222
timestamp 1701704242
transform 1 0 9752 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[38\].dly_stg4_223
timestamp 1701704242
transform 1 0 8004 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[39\].dly_stg3
timestamp 1701704242
transform -1 0 8096 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[39\].dly_stg4_224
timestamp 1701704242
transform 1 0 8096 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[39\].dly_stg4_225
timestamp 1701704242
transform 1 0 11500 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[39\].dly_stg4_226
timestamp 1701704242
transform 1 0 8924 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[39\].dly_stg4_227
timestamp 1701704242
transform -1 0 7544 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[40\].dly_stg3
timestamp 1701704242
transform 1 0 7176 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[40\].dly_stg4_228
timestamp 1701704242
transform 1 0 9752 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[40\].dly_stg4_229
timestamp 1701704242
transform 1 0 10304 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[40\].dly_stg4_230
timestamp 1701704242
transform 1 0 11132 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[40\].dly_stg4_231
timestamp 1701704242
transform 1 0 12236 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[41\].dly_stg3
timestamp 1701704242
transform 1 0 7544 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[41\].dly_stg4_232
timestamp 1701704242
transform 1 0 12696 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[41\].dly_stg4_233
timestamp 1701704242
transform 1 0 10028 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[41\].dly_stg4_234
timestamp 1701704242
transform 1 0 8372 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[41\].dly_stg4_235
timestamp 1701704242
transform 1 0 7820 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[42\].dly_stg3
timestamp 1701704242
transform 1 0 8004 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[42\].dly_stg4_236
timestamp 1701704242
transform 1 0 10948 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[42\].dly_stg4_237
timestamp 1701704242
transform -1 0 7728 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[42\].dly_stg4_238
timestamp 1701704242
transform 1 0 12420 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[42\].dly_stg4_239
timestamp 1701704242
transform 1 0 8924 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[43\].dly_stg3
timestamp 1701704242
transform -1 0 10028 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[43\].dly_stg4_240
timestamp 1701704242
transform 1 0 11040 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[43\].dly_stg4_241
timestamp 1701704242
transform -1 0 9200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[43\].dly_stg4_242
timestamp 1701704242
transform 1 0 13064 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[43\].dly_stg4_243
timestamp 1701704242
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[44\].dly_stg3
timestamp 1701704242
transform 1 0 10028 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[44\].dly_stg4_244
timestamp 1701704242
transform -1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[44\].dly_stg4_245
timestamp 1701704242
transform 1 0 13156 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[44\].dly_stg4_246
timestamp 1701704242
transform -1 0 13800 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[44\].dly_stg4_247
timestamp 1701704242
transform 1 0 11684 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[45\].dly_stg3
timestamp 1701704242
transform 1 0 11868 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[45\].dly_stg4_248
timestamp 1701704242
transform 1 0 13524 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[45\].dly_stg4_249
timestamp 1701704242
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[45\].dly_stg4_250
timestamp 1701704242
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[45\].dly_stg4_251
timestamp 1701704242
transform 1 0 11592 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[46\].dly_stg3
timestamp 1701704242
transform 1 0 13248 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[46\].dly_stg4_252
timestamp 1701704242
transform 1 0 14628 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[46\].dly_stg4_253
timestamp 1701704242
transform 1 0 12880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[46\].dly_stg4_254
timestamp 1701704242
transform -1 0 14352 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[46\].dly_stg4_255
timestamp 1701704242
transform -1 0 16376 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[47\].dly_stg3
timestamp 1701704242
transform -1 0 13892 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[47\].dly_stg4_256
timestamp 1701704242
transform -1 0 19320 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[47\].dly_stg4_257
timestamp 1701704242
transform 1 0 15916 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[47\].dly_stg4_258
timestamp 1701704242
transform 1 0 14444 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[47\].dly_stg4_259
timestamp 1701704242
transform -1 0 17204 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[48\].dly_stg3
timestamp 1701704242
transform -1 0 15456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[48\].dly_stg4_260
timestamp 1701704242
transform 1 0 18676 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[48\].dly_stg4_261
timestamp 1701704242
transform 1 0 16652 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[48\].dly_stg4_262
timestamp 1701704242
transform 1 0 16100 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[48\].dly_stg4_263
timestamp 1701704242
transform 1 0 19688 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[49\].dly_stg3
timestamp 1701704242
transform 1 0 15456 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[49\].dly_stg4_264
timestamp 1701704242
transform -1 0 16468 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[49\].dly_stg4_265
timestamp 1701704242
transform 1 0 16652 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[49\].dly_stg4_266
timestamp 1701704242
transform -1 0 14996 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[49\].dly_stg4_267
timestamp 1701704242
transform 1 0 18952 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[50\].dly_stg3
timestamp 1701704242
transform -1 0 18492 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[50\].dly_stg4_268
timestamp 1701704242
transform -1 0 15456 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[50\].dly_stg4_269
timestamp 1701704242
transform -1 0 16192 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[50\].dly_stg4_270
timestamp 1701704242
transform 1 0 16376 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[50\].dly_stg4_271
timestamp 1701704242
transform -1 0 18768 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[51\].dly_stg3
timestamp 1701704242
transform -1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[51\].dly_stg4_272
timestamp 1701704242
transform -1 0 13432 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[51\].dly_stg4_273
timestamp 1701704242
transform -1 0 15732 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[51\].dly_stg4_274
timestamp 1701704242
transform 1 0 14904 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[51\].dly_stg4_275
timestamp 1701704242
transform -1 0 17940 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[52\].dly_stg3
timestamp 1701704242
transform 1 0 13524 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[52\].dly_stg4_276
timestamp 1701704242
transform 1 0 13984 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[52\].dly_stg4_277
timestamp 1701704242
transform -1 0 15180 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[52\].dly_stg4_278
timestamp 1701704242
transform -1 0 12880 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[52\].dly_stg4_279
timestamp 1701704242
transform -1 0 15732 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[53\].dly_stg3
timestamp 1701704242
transform 1 0 12328 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[53\].dly_stg4_280
timestamp 1701704242
transform -1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[53\].dly_stg4_281
timestamp 1701704242
transform -1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[53\].dly_stg4_282
timestamp 1701704242
transform 1 0 13708 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[53\].dly_stg4_283
timestamp 1701704242
transform -1 0 11500 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[54\].dly_stg3
timestamp 1701704242
transform 1 0 11500 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[54\].dly_stg4_284
timestamp 1701704242
transform -1 0 10856 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[54\].dly_stg4_285
timestamp 1701704242
transform -1 0 13800 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[54\].dly_stg4_286
timestamp 1701704242
transform -1 0 11316 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[54\].dly_stg4_287
timestamp 1701704242
transform 1 0 13248 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[55\].dly_stg3
timestamp 1701704242
transform 1 0 10948 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[55\].dly_stg4_288
timestamp 1701704242
transform -1 0 10304 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[55\].dly_stg4_289
timestamp 1701704242
transform -1 0 12328 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[55\].dly_stg4_290
timestamp 1701704242
transform -1 0 9476 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[55\].dly_stg4_291
timestamp 1701704242
transform 1 0 10028 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[56\].dly_stg3
timestamp 1701704242
transform -1 0 9016 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[56\].dly_stg4_292
timestamp 1701704242
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[56\].dly_stg4_293
timestamp 1701704242
transform -1 0 10028 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[56\].dly_stg4_294
timestamp 1701704242
transform -1 0 9200 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[56\].dly_stg4_295
timestamp 1701704242
transform -1 0 9752 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[57\].dly_stg3
timestamp 1701704242
transform 1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[57\].dly_stg4_296
timestamp 1701704242
transform -1 0 7544 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[57\].dly_stg4_297
timestamp 1701704242
transform -1 0 8648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[57\].dly_stg4_298
timestamp 1701704242
transform -1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[57\].dly_stg4_299
timestamp 1701704242
transform -1 0 8004 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[58\].dly_stg3
timestamp 1701704242
transform -1 0 7636 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[58\].dly_stg4_300
timestamp 1701704242
transform -1 0 8372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[58\].dly_stg4_301
timestamp 1701704242
transform -1 0 8280 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[58\].dly_stg4_302
timestamp 1701704242
transform 1 0 6716 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[58\].dly_stg4_303
timestamp 1701704242
transform -1 0 6624 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[59\].dly_stg3
timestamp 1701704242
transform 1 0 6440 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[59\].dly_stg4_304
timestamp 1701704242
transform 1 0 8648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[59\].dly_stg4_305
timestamp 1701704242
transform 1 0 8464 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[59\].dly_stg4_306
timestamp 1701704242
transform 1 0 8372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[59\].dly_stg4_307
timestamp 1701704242
transform -1 0 10028 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[60\].dly_stg3
timestamp 1701704242
transform -1 0 8924 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[60\].dly_stg4_308
timestamp 1701704242
transform -1 0 7268 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[60\].dly_stg4_309
timestamp 1701704242
transform 1 0 8096 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[60\].dly_stg4_310
timestamp 1701704242
transform -1 0 9476 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[60\].dly_stg4_311
timestamp 1701704242
transform -1 0 6900 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[61\].dly_stg3
timestamp 1701704242
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[61\].dly_stg4_312
timestamp 1701704242
transform 1 0 8924 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[61\].dly_stg4_313
timestamp 1701704242
transform -1 0 7728 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[61\].dly_stg4_314
timestamp 1701704242
transform -1 0 8740 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[61\].dly_stg4_315
timestamp 1701704242
transform 1 0 10580 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[62\].dly_stg3
timestamp 1701704242
transform -1 0 10856 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[62\].dly_stg4_773
timestamp 1701704242
transform -1 0 8096 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_479
timestamp 1701704242
transform 1 0 11868 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_480
timestamp 1701704242
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_481
timestamp 1701704242
transform -1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_482
timestamp 1701704242
transform 1 0 12972 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_483
timestamp 1701704242
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_484
timestamp 1701704242
transform -1 0 12420 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg8_632
timestamp 1701704242
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_323
timestamp 1701704242
transform -1 0 15732 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_324
timestamp 1701704242
transform 1 0 16468 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_325
timestamp 1701704242
transform -1 0 13892 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_326
timestamp 1701704242
transform -1 0 15640 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_327
timestamp 1701704242
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_328
timestamp 1701704242
transform 1 0 13708 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg8_485
timestamp 1701704242
transform 1 0 15180 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_633
timestamp 1701704242
transform 1 0 17940 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_634
timestamp 1701704242
transform -1 0 17020 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_635
timestamp 1701704242
transform -1 0 16192 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_636
timestamp 1701704242
transform 1 0 20148 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_637
timestamp 1701704242
transform -1 0 19228 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_638
timestamp 1701704242
transform -1 0 18492 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg8_329
timestamp 1701704242
transform 1 0 15732 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_486
timestamp 1701704242
transform 1 0 19504 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_487
timestamp 1701704242
transform 1 0 20424 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_488
timestamp 1701704242
transform 1 0 18676 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_489
timestamp 1701704242
transform -1 0 20332 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_490
timestamp 1701704242
transform -1 0 19044 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_491
timestamp 1701704242
transform -1 0 16468 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg8_639
timestamp 1701704242
transform -1 0 17940 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_330
timestamp 1701704242
transform -1 0 15364 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_331
timestamp 1701704242
transform 1 0 20608 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_332
timestamp 1701704242
transform 1 0 18952 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_333
timestamp 1701704242
transform 1 0 21160 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_334
timestamp 1701704242
transform 1 0 18952 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_335
timestamp 1701704242
transform -1 0 20056 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg8_492
timestamp 1701704242
transform -1 0 18216 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_640
timestamp 1701704242
transform -1 0 18952 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_641
timestamp 1701704242
transform 1 0 21068 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_642
timestamp 1701704242
transform -1 0 19872 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_643
timestamp 1701704242
transform 1 0 20516 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_644
timestamp 1701704242
transform -1 0 21160 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_645
timestamp 1701704242
transform 1 0 20148 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg8_336
timestamp 1701704242
transform 1 0 20332 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_493
timestamp 1701704242
transform 1 0 19872 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_494
timestamp 1701704242
transform -1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_495
timestamp 1701704242
transform 1 0 19964 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_496
timestamp 1701704242
transform 1 0 23920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_497
timestamp 1701704242
transform -1 0 20332 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_498
timestamp 1701704242
transform -1 0 19688 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg8_646
timestamp 1701704242
transform -1 0 20516 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_337
timestamp 1701704242
transform -1 0 25484 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_338
timestamp 1701704242
transform -1 0 25760 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_339
timestamp 1701704242
transform -1 0 20976 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_340
timestamp 1701704242
transform 1 0 26036 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_341
timestamp 1701704242
transform -1 0 22080 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_342
timestamp 1701704242
transform -1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg8_499
timestamp 1701704242
transform -1 0 20056 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_647
timestamp 1701704242
transform 1 0 24748 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_648
timestamp 1701704242
transform 1 0 25760 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_649
timestamp 1701704242
transform 1 0 23828 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_650
timestamp 1701704242
transform -1 0 23092 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_651
timestamp 1701704242
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_652
timestamp 1701704242
transform 1 0 22632 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg8_343
timestamp 1701704242
transform -1 0 21068 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_500
timestamp 1701704242
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_501
timestamp 1701704242
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_502
timestamp 1701704242
transform 1 0 22724 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_503
timestamp 1701704242
transform -1 0 24380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_504
timestamp 1701704242
transform 1 0 24196 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_505
timestamp 1701704242
transform 1 0 22172 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg8_653
timestamp 1701704242
transform 1 0 24932 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_344
timestamp 1701704242
transform 1 0 26036 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_345
timestamp 1701704242
transform -1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_346
timestamp 1701704242
transform 1 0 25208 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_347
timestamp 1701704242
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_348
timestamp 1701704242
transform -1 0 25760 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_349
timestamp 1701704242
transform -1 0 25208 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg8_506
timestamp 1701704242
transform 1 0 25760 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_654
timestamp 1701704242
transform -1 0 20516 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_655
timestamp 1701704242
transform 1 0 24656 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_656
timestamp 1701704242
transform 1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_657
timestamp 1701704242
transform 1 0 20516 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_658
timestamp 1701704242
transform -1 0 22724 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_659
timestamp 1701704242
transform -1 0 20608 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg8_350
timestamp 1701704242
transform -1 0 22172 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_507
timestamp 1701704242
transform 1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_508
timestamp 1701704242
transform 1 0 21804 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_509
timestamp 1701704242
transform -1 0 23736 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_510
timestamp 1701704242
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_511
timestamp 1701704242
transform -1 0 25944 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_512
timestamp 1701704242
transform 1 0 24840 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg8_660
timestamp 1701704242
transform -1 0 21804 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg7_351
timestamp 1701704242
transform 1 0 25944 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg7_352
timestamp 1701704242
transform 1 0 24564 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg7_353
timestamp 1701704242
transform 1 0 26036 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg7_354
timestamp 1701704242
transform 1 0 21528 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg7_355
timestamp 1701704242
transform 1 0 23276 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg7_356
timestamp 1701704242
transform -1 0 21068 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg8_513
timestamp 1701704242
transform -1 0 25668 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[14\].dly_stg7_661
timestamp 1701704242
transform -1 0 25484 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[14\].dly_stg7_662
timestamp 1701704242
transform -1 0 21436 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[14\].dly_stg7_663
timestamp 1701704242
transform 1 0 24012 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[14\].dly_stg7_664
timestamp 1701704242
transform 1 0 23368 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[14\].dly_stg7_665
timestamp 1701704242
transform -1 0 24472 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[14\].dly_stg7_666
timestamp 1701704242
transform 1 0 24104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[14\].dly_stg8_357
timestamp 1701704242
transform 1 0 24288 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[15\].dly_stg7_514
timestamp 1701704242
transform 1 0 25300 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[15\].dly_stg7_515
timestamp 1701704242
transform 1 0 21344 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[15\].dly_stg7_516
timestamp 1701704242
transform 1 0 23644 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[15\].dly_stg7_517
timestamp 1701704242
transform -1 0 24104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[15\].dly_stg7_518
timestamp 1701704242
transform -1 0 20424 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[15\].dly_stg7_519
timestamp 1701704242
transform -1 0 21988 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[15\].dly_stg8_667
timestamp 1701704242
transform -1 0 24380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[16\].dly_stg7_358
timestamp 1701704242
transform -1 0 19780 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[16\].dly_stg7_359
timestamp 1701704242
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[16\].dly_stg7_360
timestamp 1701704242
transform -1 0 21804 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[16\].dly_stg7_361
timestamp 1701704242
transform 1 0 20240 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[16\].dly_stg7_362
timestamp 1701704242
transform 1 0 24380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[16\].dly_stg7_363
timestamp 1701704242
transform -1 0 22172 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[16\].dly_stg8_520
timestamp 1701704242
transform 1 0 21804 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[17\].dly_stg7_668
timestamp 1701704242
transform 1 0 25760 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[17\].dly_stg7_669
timestamp 1701704242
transform -1 0 25208 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[17\].dly_stg7_670
timestamp 1701704242
transform 1 0 24472 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[17\].dly_stg7_671
timestamp 1701704242
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[17\].dly_stg7_672
timestamp 1701704242
transform -1 0 21804 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[17\].dly_stg7_673
timestamp 1701704242
transform -1 0 21252 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[17\].dly_stg8_364
timestamp 1701704242
transform 1 0 24748 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[18\].dly_stg7_521
timestamp 1701704242
transform -1 0 20240 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[18\].dly_stg7_522
timestamp 1701704242
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[18\].dly_stg7_523
timestamp 1701704242
transform 1 0 21804 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[18\].dly_stg7_524
timestamp 1701704242
transform 1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[18\].dly_stg7_525
timestamp 1701704242
transform -1 0 20976 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[18\].dly_stg7_526
timestamp 1701704242
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[18\].dly_stg8_674
timestamp 1701704242
transform -1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[19\].dly_stg7_365
timestamp 1701704242
transform 1 0 25484 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[19\].dly_stg7_366
timestamp 1701704242
transform -1 0 25484 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[19\].dly_stg7_367
timestamp 1701704242
transform -1 0 21528 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[19\].dly_stg7_368
timestamp 1701704242
transform 1 0 26312 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[19\].dly_stg7_369
timestamp 1701704242
transform 1 0 21528 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[19\].dly_stg7_370
timestamp 1701704242
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[19\].dly_stg8_527
timestamp 1701704242
transform -1 0 20700 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[20\].dly_stg7_675
timestamp 1701704242
transform -1 0 20792 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[20\].dly_stg7_676
timestamp 1701704242
transform -1 0 24932 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[20\].dly_stg7_677
timestamp 1701704242
transform -1 0 22080 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[20\].dly_stg7_678
timestamp 1701704242
transform 1 0 25576 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[20\].dly_stg7_679
timestamp 1701704242
transform -1 0 24104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[20\].dly_stg7_680
timestamp 1701704242
transform 1 0 24656 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[20\].dly_stg8_371
timestamp 1701704242
transform 1 0 24380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[21\].dly_stg7_528
timestamp 1701704242
transform 1 0 26588 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[21\].dly_stg7_529
timestamp 1701704242
transform 1 0 22540 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[21\].dly_stg7_530
timestamp 1701704242
transform -1 0 26036 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[21\].dly_stg7_531
timestamp 1701704242
transform -1 0 25576 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[21\].dly_stg7_532
timestamp 1701704242
transform -1 0 20792 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[21\].dly_stg7_533
timestamp 1701704242
transform 1 0 21528 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[21\].dly_stg8_681
timestamp 1701704242
transform -1 0 22356 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[22\].dly_stg7_372
timestamp 1701704242
transform 1 0 26404 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[22\].dly_stg7_373
timestamp 1701704242
transform 1 0 24104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[22\].dly_stg7_374
timestamp 1701704242
transform -1 0 21528 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[22\].dly_stg7_375
timestamp 1701704242
transform -1 0 25852 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[22\].dly_stg7_376
timestamp 1701704242
transform 1 0 25024 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[22\].dly_stg7_377
timestamp 1701704242
transform -1 0 25484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[22\].dly_stg8_534
timestamp 1701704242
transform 1 0 23828 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[23\].dly_stg7_682
timestamp 1701704242
transform 1 0 25484 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[23\].dly_stg7_683
timestamp 1701704242
transform -1 0 25760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[23\].dly_stg7_684
timestamp 1701704242
transform 1 0 25760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[23\].dly_stg7_685
timestamp 1701704242
transform 1 0 24564 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[23\].dly_stg7_686
timestamp 1701704242
transform -1 0 23644 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[23\].dly_stg7_687
timestamp 1701704242
transform -1 0 25484 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[23\].dly_stg8_378
timestamp 1701704242
transform 1 0 26036 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[24\].dly_stg7_535
timestamp 1701704242
transform 1 0 24104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[24\].dly_stg7_536
timestamp 1701704242
transform -1 0 24380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[24\].dly_stg7_537
timestamp 1701704242
transform 1 0 24288 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[24\].dly_stg7_538
timestamp 1701704242
transform -1 0 24288 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[24\].dly_stg7_539
timestamp 1701704242
transform 1 0 22356 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[24\].dly_stg7_540
timestamp 1701704242
transform -1 0 21988 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[24\].dly_stg8_688
timestamp 1701704242
transform 1 0 24932 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[25\].dly_stg7_379
timestamp 1701704242
transform -1 0 24656 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[25\].dly_stg7_380
timestamp 1701704242
transform -1 0 23736 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[25\].dly_stg7_381
timestamp 1701704242
transform 1 0 23828 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[25\].dly_stg7_382
timestamp 1701704242
transform -1 0 22908 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[25\].dly_stg7_383
timestamp 1701704242
transform -1 0 24196 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[25\].dly_stg7_384
timestamp 1701704242
transform -1 0 20792 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[25\].dly_stg8_541
timestamp 1701704242
transform 1 0 22632 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[26\].dly_stg7_689
timestamp 1701704242
transform 1 0 24840 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[26\].dly_stg7_690
timestamp 1701704242
transform -1 0 22632 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[26\].dly_stg7_691
timestamp 1701704242
transform -1 0 21068 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[26\].dly_stg7_692
timestamp 1701704242
transform -1 0 20700 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[26\].dly_stg7_693
timestamp 1701704242
transform 1 0 22080 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[26\].dly_stg7_694
timestamp 1701704242
transform 1 0 22264 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[26\].dly_stg8_385
timestamp 1701704242
transform -1 0 23184 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[27\].dly_stg7_542
timestamp 1701704242
transform 1 0 20608 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[27\].dly_stg7_543
timestamp 1701704242
transform -1 0 21436 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[27\].dly_stg7_544
timestamp 1701704242
transform -1 0 23184 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[27\].dly_stg7_545
timestamp 1701704242
transform -1 0 19320 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[27\].dly_stg7_546
timestamp 1701704242
transform 1 0 23828 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[27\].dly_stg7_547
timestamp 1701704242
transform 1 0 20976 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[27\].dly_stg8_695
timestamp 1701704242
transform 1 0 23184 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[28\].dly_stg7_386
timestamp 1701704242
transform -1 0 19044 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[28\].dly_stg7_387
timestamp 1701704242
transform -1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[28\].dly_stg7_388
timestamp 1701704242
transform -1 0 22080 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[28\].dly_stg7_389
timestamp 1701704242
transform 1 0 19964 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[28\].dly_stg7_390
timestamp 1701704242
transform -1 0 22356 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[28\].dly_stg7_391
timestamp 1701704242
transform 1 0 19596 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[28\].dly_stg8_548
timestamp 1701704242
transform -1 0 22356 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[29\].dly_stg7_696
timestamp 1701704242
transform 1 0 20792 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[29\].dly_stg7_697
timestamp 1701704242
transform -1 0 19136 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[29\].dly_stg7_698
timestamp 1701704242
transform -1 0 20332 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[29\].dly_stg7_699
timestamp 1701704242
transform -1 0 18308 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[29\].dly_stg7_700
timestamp 1701704242
transform 1 0 18308 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[29\].dly_stg7_701
timestamp 1701704242
transform 1 0 18952 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[29\].dly_stg8_392
timestamp 1701704242
transform -1 0 20608 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[30\].dly_stg7_549
timestamp 1701704242
transform -1 0 17572 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[30\].dly_stg7_550
timestamp 1701704242
transform -1 0 17756 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[30\].dly_stg7_551
timestamp 1701704242
transform -1 0 18952 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[30\].dly_stg7_552
timestamp 1701704242
transform -1 0 18032 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[30\].dly_stg7_553
timestamp 1701704242
transform 1 0 17756 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[30\].dly_stg7_554
timestamp 1701704242
transform -1 0 20792 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[30\].dly_stg8_702
timestamp 1701704242
transform 1 0 19688 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[31\].dly_stg7_393
timestamp 1701704242
transform -1 0 18584 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[31\].dly_stg7_394
timestamp 1701704242
transform 1 0 16560 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[31\].dly_stg7_395
timestamp 1701704242
transform 1 0 18308 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[31\].dly_stg7_396
timestamp 1701704242
transform -1 0 15732 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[31\].dly_stg7_397
timestamp 1701704242
transform -1 0 18308 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[31\].dly_stg7_398
timestamp 1701704242
transform 1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[31\].dly_stg8_555
timestamp 1701704242
transform 1 0 19964 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[32\].dly_stg7_703
timestamp 1701704242
transform -1 0 16376 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[32\].dly_stg7_704
timestamp 1701704242
transform -1 0 13524 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[32\].dly_stg7_705
timestamp 1701704242
transform 1 0 16928 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[32\].dly_stg7_706
timestamp 1701704242
transform 1 0 13984 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[32\].dly_stg7_707
timestamp 1701704242
transform 1 0 16928 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[32\].dly_stg7_708
timestamp 1701704242
transform -1 0 16284 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[32\].dly_stg8_399
timestamp 1701704242
transform 1 0 18032 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[33\].dly_stg7_556
timestamp 1701704242
transform -1 0 15272 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[33\].dly_stg7_557
timestamp 1701704242
transform -1 0 14444 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[33\].dly_stg7_558
timestamp 1701704242
transform 1 0 16376 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[33\].dly_stg7_559
timestamp 1701704242
transform 1 0 13616 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[33\].dly_stg7_560
timestamp 1701704242
transform -1 0 14536 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[33\].dly_stg7_561
timestamp 1701704242
transform 1 0 14996 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[33\].dly_stg8_709
timestamp 1701704242
transform 1 0 18308 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[34\].dly_stg7_400
timestamp 1701704242
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[34\].dly_stg7_401
timestamp 1701704242
transform -1 0 13800 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[34\].dly_stg7_402
timestamp 1701704242
transform 1 0 14444 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[34\].dly_stg7_403
timestamp 1701704242
transform -1 0 13524 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[34\].dly_stg7_404
timestamp 1701704242
transform 1 0 13708 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[34\].dly_stg7_405
timestamp 1701704242
transform 1 0 13432 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[34\].dly_stg8_562
timestamp 1701704242
transform -1 0 14260 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[35\].dly_stg7_710
timestamp 1701704242
transform 1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[35\].dly_stg7_711
timestamp 1701704242
transform -1 0 12696 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[35\].dly_stg7_712
timestamp 1701704242
transform -1 0 13248 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[35\].dly_stg7_713
timestamp 1701704242
transform 1 0 10948 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[35\].dly_stg7_714
timestamp 1701704242
transform 1 0 11316 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[35\].dly_stg7_715
timestamp 1701704242
transform -1 0 10856 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[35\].dly_stg8_406
timestamp 1701704242
transform 1 0 13800 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[36\].dly_stg7_563
timestamp 1701704242
transform -1 0 11224 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[36\].dly_stg7_564
timestamp 1701704242
transform -1 0 11776 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[36\].dly_stg7_565
timestamp 1701704242
transform -1 0 12328 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[36\].dly_stg7_566
timestamp 1701704242
transform -1 0 11684 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[36\].dly_stg7_567
timestamp 1701704242
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[36\].dly_stg7_568
timestamp 1701704242
transform -1 0 9752 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[36\].dly_stg8_716
timestamp 1701704242
transform 1 0 12972 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[37\].dly_stg7_407
timestamp 1701704242
transform -1 0 8004 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[37\].dly_stg7_408
timestamp 1701704242
transform 1 0 8648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[37\].dly_stg7_409
timestamp 1701704242
transform 1 0 9752 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[37\].dly_stg7_410
timestamp 1701704242
transform 1 0 11684 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[37\].dly_stg7_411
timestamp 1701704242
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[37\].dly_stg7_412
timestamp 1701704242
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[37\].dly_stg8_569
timestamp 1701704242
transform 1 0 12696 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[38\].dly_stg7_717
timestamp 1701704242
transform -1 0 10212 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[38\].dly_stg7_718
timestamp 1701704242
transform -1 0 7820 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[38\].dly_stg7_719
timestamp 1701704242
transform 1 0 10028 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[38\].dly_stg7_720
timestamp 1701704242
transform -1 0 7728 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[38\].dly_stg7_721
timestamp 1701704242
transform 1 0 10580 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[38\].dly_stg7_722
timestamp 1701704242
transform 1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[38\].dly_stg8_413
timestamp 1701704242
transform 1 0 10856 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[39\].dly_stg7_570
timestamp 1701704242
transform 1 0 11960 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[39\].dly_stg7_571
timestamp 1701704242
transform -1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[39\].dly_stg7_572
timestamp 1701704242
transform 1 0 9476 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[39\].dly_stg7_573
timestamp 1701704242
transform 1 0 8556 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[39\].dly_stg7_574
timestamp 1701704242
transform -1 0 10856 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[39\].dly_stg7_575
timestamp 1701704242
transform -1 0 9476 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[39\].dly_stg8_723
timestamp 1701704242
transform -1 0 9200 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[40\].dly_stg7_414
timestamp 1701704242
transform -1 0 7544 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[40\].dly_stg7_415
timestamp 1701704242
transform 1 0 8096 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[40\].dly_stg7_416
timestamp 1701704242
transform 1 0 8648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[40\].dly_stg7_417
timestamp 1701704242
transform 1 0 9476 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[40\].dly_stg7_418
timestamp 1701704242
transform 1 0 8096 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[40\].dly_stg7_419
timestamp 1701704242
transform -1 0 9476 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[40\].dly_stg8_576
timestamp 1701704242
transform -1 0 9200 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[41\].dly_stg7_724
timestamp 1701704242
transform -1 0 9200 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[41\].dly_stg7_725
timestamp 1701704242
transform 1 0 9200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[41\].dly_stg7_726
timestamp 1701704242
transform -1 0 8096 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[41\].dly_stg7_727
timestamp 1701704242
transform 1 0 10028 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[41\].dly_stg7_728
timestamp 1701704242
transform 1 0 12144 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[41\].dly_stg7_729
timestamp 1701704242
transform -1 0 8648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[41\].dly_stg8_420
timestamp 1701704242
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[42\].dly_stg7_577
timestamp 1701704242
transform 1 0 10304 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[42\].dly_stg7_578
timestamp 1701704242
transform 1 0 10580 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[42\].dly_stg7_579
timestamp 1701704242
transform -1 0 12144 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[42\].dly_stg7_580
timestamp 1701704242
transform 1 0 10396 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[42\].dly_stg7_581
timestamp 1701704242
transform 1 0 10304 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[42\].dly_stg7_582
timestamp 1701704242
transform -1 0 9752 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[42\].dly_stg8_730
timestamp 1701704242
transform -1 0 8924 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[43\].dly_stg7_421
timestamp 1701704242
transform 1 0 11132 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[43\].dly_stg7_422
timestamp 1701704242
transform 1 0 14536 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[43\].dly_stg7_423
timestamp 1701704242
transform -1 0 10672 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[43\].dly_stg7_424
timestamp 1701704242
transform -1 0 14352 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[43\].dly_stg7_425
timestamp 1701704242
transform -1 0 11684 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[43\].dly_stg7_426
timestamp 1701704242
transform -1 0 11776 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[43\].dly_stg8_583
timestamp 1701704242
transform 1 0 10672 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[44\].dly_stg7_731
timestamp 1701704242
transform 1 0 11500 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[44\].dly_stg7_732
timestamp 1701704242
transform 1 0 12420 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[44\].dly_stg7_733
timestamp 1701704242
transform -1 0 10948 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[44\].dly_stg7_734
timestamp 1701704242
transform 1 0 12696 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[44\].dly_stg7_735
timestamp 1701704242
transform 1 0 13800 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[44\].dly_stg7_736
timestamp 1701704242
transform -1 0 13156 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[44\].dly_stg8_427
timestamp 1701704242
transform -1 0 11592 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[45\].dly_stg7_584
timestamp 1701704242
transform 1 0 16376 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[45\].dly_stg7_585
timestamp 1701704242
transform -1 0 15916 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[45\].dly_stg7_586
timestamp 1701704242
transform -1 0 12420 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[45\].dly_stg7_587
timestamp 1701704242
transform 1 0 14352 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[45\].dly_stg7_588
timestamp 1701704242
transform 1 0 16192 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[45\].dly_stg7_589
timestamp 1701704242
transform 1 0 12972 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[45\].dly_stg8_737
timestamp 1701704242
transform -1 0 13432 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[46\].dly_stg7_428
timestamp 1701704242
transform -1 0 17756 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[46\].dly_stg7_429
timestamp 1701704242
transform 1 0 13892 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[46\].dly_stg7_430
timestamp 1701704242
transform 1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[46\].dly_stg7_431
timestamp 1701704242
transform 1 0 19412 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[46\].dly_stg7_432
timestamp 1701704242
transform -1 0 16376 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[46\].dly_stg7_433
timestamp 1701704242
transform -1 0 14076 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[46\].dly_stg8_590
timestamp 1701704242
transform 1 0 16468 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[47\].dly_stg7_738
timestamp 1701704242
transform 1 0 17204 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[47\].dly_stg7_739
timestamp 1701704242
transform 1 0 14996 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[47\].dly_stg7_740
timestamp 1701704242
transform 1 0 15548 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[47\].dly_stg7_741
timestamp 1701704242
transform 1 0 17940 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[47\].dly_stg7_742
timestamp 1701704242
transform -1 0 16468 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[47\].dly_stg7_743
timestamp 1701704242
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[47\].dly_stg8_434
timestamp 1701704242
transform -1 0 15456 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[48\].dly_stg7_591
timestamp 1701704242
transform 1 0 18768 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[48\].dly_stg7_592
timestamp 1701704242
transform 1 0 19320 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[48\].dly_stg7_593
timestamp 1701704242
transform -1 0 15548 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[48\].dly_stg7_594
timestamp 1701704242
transform -1 0 16744 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[48\].dly_stg7_595
timestamp 1701704242
transform -1 0 17020 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[48\].dly_stg7_596
timestamp 1701704242
transform -1 0 17204 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[48\].dly_stg8_744
timestamp 1701704242
transform -1 0 15732 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[49\].dly_stg7_435
timestamp 1701704242
transform 1 0 19228 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[49\].dly_stg7_436
timestamp 1701704242
transform -1 0 15916 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[49\].dly_stg7_437
timestamp 1701704242
transform -1 0 16744 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[49\].dly_stg7_438
timestamp 1701704242
transform -1 0 16008 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[49\].dly_stg7_439
timestamp 1701704242
transform -1 0 18216 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[49\].dly_stg7_440
timestamp 1701704242
transform 1 0 15732 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[49\].dly_stg8_597
timestamp 1701704242
transform -1 0 16008 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[50\].dly_stg7_745
timestamp 1701704242
transform 1 0 18216 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[50\].dly_stg7_746
timestamp 1701704242
transform -1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[50\].dly_stg7_747
timestamp 1701704242
transform -1 0 17204 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[50\].dly_stg7_748
timestamp 1701704242
transform -1 0 15180 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[50\].dly_stg7_749
timestamp 1701704242
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[50\].dly_stg7_750
timestamp 1701704242
transform -1 0 16100 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[50\].dly_stg8_441
timestamp 1701704242
transform -1 0 18124 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[51\].dly_stg7_598
timestamp 1701704242
transform 1 0 18124 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[51\].dly_stg7_599
timestamp 1701704242
transform -1 0 13248 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[51\].dly_stg7_600
timestamp 1701704242
transform -1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[51\].dly_stg7_601
timestamp 1701704242
transform -1 0 12972 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[51\].dly_stg7_602
timestamp 1701704242
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[51\].dly_stg7_603
timestamp 1701704242
transform -1 0 14628 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[51\].dly_stg8_751
timestamp 1701704242
transform 1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[52\].dly_stg7_442
timestamp 1701704242
transform -1 0 12328 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[52\].dly_stg7_443
timestamp 1701704242
transform 1 0 12144 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[52\].dly_stg7_444
timestamp 1701704242
transform 1 0 14628 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[52\].dly_stg7_445
timestamp 1701704242
transform -1 0 12144 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[52\].dly_stg7_446
timestamp 1701704242
transform -1 0 14076 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[52\].dly_stg7_447
timestamp 1701704242
transform -1 0 13156 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[52\].dly_stg8_604
timestamp 1701704242
transform 1 0 14352 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[53\].dly_stg7_752
timestamp 1701704242
transform 1 0 12880 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[53\].dly_stg7_753
timestamp 1701704242
transform -1 0 12052 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[53\].dly_stg7_754
timestamp 1701704242
transform 1 0 14076 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[53\].dly_stg7_755
timestamp 1701704242
transform -1 0 11592 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[53\].dly_stg7_756
timestamp 1701704242
transform 1 0 12328 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[53\].dly_stg7_757
timestamp 1701704242
transform -1 0 13340 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[53\].dly_stg8_448
timestamp 1701704242
transform -1 0 13892 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[54\].dly_stg7_605
timestamp 1701704242
transform -1 0 10304 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[54\].dly_stg7_606
timestamp 1701704242
transform -1 0 10948 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[54\].dly_stg7_607
timestamp 1701704242
transform 1 0 12420 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[54\].dly_stg7_608
timestamp 1701704242
transform -1 0 10396 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[54\].dly_stg7_609
timestamp 1701704242
transform 1 0 10304 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[54\].dly_stg7_610
timestamp 1701704242
transform -1 0 11500 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[54\].dly_stg8_758
timestamp 1701704242
transform 1 0 12604 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[55\].dly_stg7_449
timestamp 1701704242
transform -1 0 10028 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[55\].dly_stg7_450
timestamp 1701704242
transform -1 0 9476 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[55\].dly_stg7_451
timestamp 1701704242
transform 1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[55\].dly_stg7_452
timestamp 1701704242
transform 1 0 10396 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[55\].dly_stg7_453
timestamp 1701704242
transform -1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[55\].dly_stg7_454
timestamp 1701704242
transform -1 0 9200 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[55\].dly_stg8_611
timestamp 1701704242
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[56\].dly_stg7_759
timestamp 1701704242
transform -1 0 8924 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[56\].dly_stg7_760
timestamp 1701704242
transform -1 0 9476 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[56\].dly_stg7_761
timestamp 1701704242
transform -1 0 9752 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[56\].dly_stg7_762
timestamp 1701704242
transform -1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[56\].dly_stg7_763
timestamp 1701704242
transform 1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[56\].dly_stg7_764
timestamp 1701704242
transform -1 0 8280 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[56\].dly_stg8_455
timestamp 1701704242
transform -1 0 10028 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[57\].dly_stg7_612
timestamp 1701704242
transform -1 0 7360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[57\].dly_stg7_613
timestamp 1701704242
transform -1 0 6900 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[57\].dly_stg7_614
timestamp 1701704242
transform -1 0 8464 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[57\].dly_stg7_615
timestamp 1701704242
transform -1 0 9016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[57\].dly_stg7_616
timestamp 1701704242
transform 1 0 7452 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[57\].dly_stg7_617
timestamp 1701704242
transform 1 0 7176 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[57\].dly_stg8_765
timestamp 1701704242
transform -1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[58\].dly_stg7_456
timestamp 1701704242
transform 1 0 10764 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[58\].dly_stg7_457
timestamp 1701704242
transform 1 0 7544 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[58\].dly_stg7_458
timestamp 1701704242
transform 1 0 8372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[58\].dly_stg7_459
timestamp 1701704242
transform 1 0 7820 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[58\].dly_stg7_460
timestamp 1701704242
transform -1 0 6348 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[58\].dly_stg7_461
timestamp 1701704242
transform -1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[58\].dly_stg8_618
timestamp 1701704242
transform 1 0 8924 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[59\].dly_stg7_766
timestamp 1701704242
transform -1 0 7176 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[59\].dly_stg7_767
timestamp 1701704242
transform 1 0 9476 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[59\].dly_stg7_768
timestamp 1701704242
transform 1 0 7452 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[59\].dly_stg7_769
timestamp 1701704242
transform -1 0 7544 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[59\].dly_stg7_770
timestamp 1701704242
transform 1 0 8004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[59\].dly_stg7_771
timestamp 1701704242
transform 1 0 7728 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[59\].dly_stg8_462
timestamp 1701704242
transform 1 0 8372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[60\].dly_stg7_619
timestamp 1701704242
transform 1 0 10488 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[60\].dly_stg7_620
timestamp 1701704242
transform 1 0 10764 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[60\].dly_stg7_621
timestamp 1701704242
transform -1 0 7820 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[60\].dly_stg7_622
timestamp 1701704242
transform 1 0 8096 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[60\].dly_stg7_623
timestamp 1701704242
transform -1 0 7452 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[60\].dly_stg7_624
timestamp 1701704242
transform -1 0 9752 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[60\].dly_stg8_772
timestamp 1701704242
transform 1 0 8648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[61\].dly_stg7_463
timestamp 1701704242
transform 1 0 8096 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[61\].dly_stg7_464
timestamp 1701704242
transform 1 0 7820 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[61\].dly_stg7_465
timestamp 1701704242
transform -1 0 7176 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[61\].dly_stg8_625
timestamp 1701704242
transform -1 0 8648 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[61\].dly_stg8_626
timestamp 1701704242
transform -1 0 8280 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[61\].dly_stg8_627
timestamp 1701704242
transform 1 0 11040 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[61\].dly_stg8_628
timestamp 1701704242
transform 1 0 11684 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[0\].dly_stp_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7728 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[1\].dly_stp_2
timestamp 1701704242
transform -1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[2\].dly_stp_3
timestamp 1701704242
transform 1 0 7452 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[3\].dly_stp_4
timestamp 1701704242
transform -1 0 8924 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[4\].dly_stp_5
timestamp 1701704242
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[5\].dly_stp_6
timestamp 1701704242
transform -1 0 9476 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[6\].dly_stp_7
timestamp 1701704242
transform 1 0 7728 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[7\].dly_stp_8
timestamp 1701704242
transform 1 0 9200 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[0\].dly_strt
timestamp 1701704242
transform -1 0 9016 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[1\].dly_strt
timestamp 1701704242
transform 1 0 6716 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[2\].dly_strt
timestamp 1701704242
transform -1 0 8188 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[3\].dly_strt
timestamp 1701704242
transform 1 0 6440 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[4\].dly_strt
timestamp 1701704242
transform 1 0 7636 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[5\].dly_strt
timestamp 1701704242
transform -1 0 8004 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[6\].dly_strt
timestamp 1701704242
transform 1 0 6164 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[7\].dly_strt
timestamp 1701704242
transform -1 0 7728 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[8\].dly_strt
timestamp 1701704242
transform -1 0 7452 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[9\].dly_strt
timestamp 1701704242
transform -1 0 6624 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[10\].dly_strt
timestamp 1701704242
transform 1 0 6072 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[11\].dly_strt
timestamp 1701704242
transform -1 0 8280 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[12\].dly_strt
timestamp 1701704242
transform -1 0 7544 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[13\].dly_strt
timestamp 1701704242
transform 1 0 6624 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[14\].dly_strt
timestamp 1701704242
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[15\].dly_strt
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7820 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_59
timestamp 1701704242
transform -1 0 21068 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_60
timestamp 1701704242
transform -1 0 12880 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_61
timestamp 1701704242
transform -1 0 24380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_62
timestamp 1701704242
transform -1 0 21528 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_63
timestamp 1701704242
transform -1 0 22448 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_64
timestamp 1701704242
transform -1 0 21712 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_65
timestamp 1701704242
transform 1 0 24932 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_66
timestamp 1701704242
transform 1 0 22080 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_67
timestamp 1701704242
transform 1 0 25760 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_68
timestamp 1701704242
transform -1 0 20332 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_69
timestamp 1701704242
transform -1 0 24932 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_70
timestamp 1701704242
transform 1 0 23828 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net59_71
timestamp 1701704242
transform -1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 31372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 31372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 31372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 31372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 31372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 31372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 31372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 31372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 31372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 31372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 31372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 31372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 31372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 31372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 31372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 31372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 31372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 31372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1701704242
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 31372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1701704242
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 31372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1701704242
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 31372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1701704242
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 31372 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1701704242
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 31372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1701704242
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 31372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1701704242
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 31372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1701704242
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 31372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1701704242
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 31372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1701704242
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 31372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1701704242
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 31372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1701704242
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 31372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1701704242
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 31372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1701704242
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1701704242
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1701704242
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1701704242
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1701704242
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1701704242
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1701704242
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1701704242
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1701704242
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_82
timestamp 1701704242
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp 1701704242
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 1701704242
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 1701704242
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 1701704242
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 1701704242
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 1701704242
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp 1701704242
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 1701704242
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_97
timestamp 1701704242
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 1701704242
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 1701704242
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 1701704242
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_101
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_103
timestamp 1701704242
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_104
timestamp 1701704242
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_105
timestamp 1701704242
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_108
timestamp 1701704242
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_109
timestamp 1701704242
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_110
timestamp 1701704242
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_111
timestamp 1701704242
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_112
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_113
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_114
timestamp 1701704242
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_115
timestamp 1701704242
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1701704242
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_117
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_118
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_119
timestamp 1701704242
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1701704242
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1701704242
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1701704242
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_123
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1701704242
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1701704242
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1701704242
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1701704242
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1701704242
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_132
timestamp 1701704242
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_133
timestamp 1701704242
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp 1701704242
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp 1701704242
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp 1701704242
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_140
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_141
timestamp 1701704242
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_142
timestamp 1701704242
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_143
timestamp 1701704242
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_144
timestamp 1701704242
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_145
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_146
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_147
timestamp 1701704242
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_148
timestamp 1701704242
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_149
timestamp 1701704242
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_150
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_152
timestamp 1701704242
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_153
timestamp 1701704242
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_154
timestamp 1701704242
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_155
timestamp 1701704242
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_156
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_157
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_158
timestamp 1701704242
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_159
timestamp 1701704242
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 1701704242
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_162
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_163
timestamp 1701704242
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 1701704242
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 1701704242
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 1701704242
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_167
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_168
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 1701704242
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_170
timestamp 1701704242
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 1701704242
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_172
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 1701704242
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 1701704242
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 1701704242
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 1701704242
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 1701704242
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 1701704242
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 1701704242
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_183
timestamp 1701704242
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_184
timestamp 1701704242
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_185
timestamp 1701704242
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 1701704242
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 1701704242
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 1701704242
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 1701704242
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_190
timestamp 1701704242
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_191
timestamp 1701704242
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_192
timestamp 1701704242
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 1701704242
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_194
timestamp 1701704242
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1701704242
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 1701704242
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 1701704242
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 1701704242
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 1701704242
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_200
timestamp 1701704242
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_201
timestamp 1701704242
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 1701704242
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 1701704242
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 1701704242
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_205
timestamp 1701704242
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 1701704242
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 1701704242
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 1701704242
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_209
timestamp 1701704242
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_210
timestamp 1701704242
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 1701704242
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 1701704242
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_213
timestamp 1701704242
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_214
timestamp 1701704242
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_215
timestamp 1701704242
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 1701704242
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 1701704242
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_218
timestamp 1701704242
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_219
timestamp 1701704242
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_220
timestamp 1701704242
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_221
timestamp 1701704242
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_222
timestamp 1701704242
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_223
timestamp 1701704242
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_224
timestamp 1701704242
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_225
timestamp 1701704242
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_226
timestamp 1701704242
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_227
timestamp 1701704242
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_228
timestamp 1701704242
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_229
timestamp 1701704242
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_230
timestamp 1701704242
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_231
timestamp 1701704242
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_232
timestamp 1701704242
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_233
timestamp 1701704242
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_234
timestamp 1701704242
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_235
timestamp 1701704242
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_236
timestamp 1701704242
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_237
timestamp 1701704242
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_238
timestamp 1701704242
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_239
timestamp 1701704242
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_240
timestamp 1701704242
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_241
timestamp 1701704242
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_242
timestamp 1701704242
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_243
timestamp 1701704242
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_244
timestamp 1701704242
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_245
timestamp 1701704242
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_246
timestamp 1701704242
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_247
timestamp 1701704242
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_248
timestamp 1701704242
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_249
timestamp 1701704242
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_250
timestamp 1701704242
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_251
timestamp 1701704242
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_252
timestamp 1701704242
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_253
timestamp 1701704242
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_254
timestamp 1701704242
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_255
timestamp 1701704242
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_256
timestamp 1701704242
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_257
timestamp 1701704242
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_258
timestamp 1701704242
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_259
timestamp 1701704242
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_260
timestamp 1701704242
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_261
timestamp 1701704242
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_262
timestamp 1701704242
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_263
timestamp 1701704242
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp 1701704242
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1701704242
transform 1 0 28888 0 -1 19040
box -38 -48 130 592
<< labels >>
flabel metal4 s 8096 496 8416 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15801 496 16121 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23506 496 23826 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 31211 496 31531 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4244 496 4564 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11949 496 12269 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19654 496 19974 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 27359 496 27679 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 7746 0 7802 400 0 FreeSans 224 90 0 0 i_start
port 2 nsew signal input
flabel metal2 s 8390 0 8446 400 0 FreeSans 224 90 0 0 i_stop
port 3 nsew signal input
flabel metal2 s 23202 0 23258 400 0 FreeSans 224 90 0 0 o_result_ctr[0]
port 4 nsew signal tristate
flabel metal2 s 21914 0 21970 400 0 FreeSans 224 90 0 0 o_result_ctr[1]
port 5 nsew signal tristate
flabel metal2 s 20626 0 20682 400 0 FreeSans 224 90 0 0 o_result_ctr[2]
port 6 nsew signal tristate
flabel metal2 s 16118 0 16174 400 0 FreeSans 224 90 0 0 o_result_ctr[3]
port 7 nsew signal tristate
flabel metal2 s 9034 0 9090 400 0 FreeSans 224 90 0 0 o_result_ctr[4]
port 8 nsew signal tristate
flabel metal2 s 10322 0 10378 400 0 FreeSans 224 90 0 0 o_result_ctr[5]
port 9 nsew signal tristate
flabel metal2 s 11610 0 11666 400 0 FreeSans 224 90 0 0 o_result_ctr[6]
port 10 nsew signal tristate
flabel metal2 s 10966 0 11022 400 0 FreeSans 224 90 0 0 o_result_ctr[7]
port 11 nsew signal tristate
flabel metal2 s 13542 0 13598 400 0 FreeSans 224 90 0 0 o_result_ring[0]
port 12 nsew signal tristate
flabel metal3 s 31600 4768 32000 4888 0 FreeSans 480 0 0 0 o_result_ring[10]
port 13 nsew signal tristate
flabel metal3 s 31600 6808 32000 6928 0 FreeSans 480 0 0 0 o_result_ring[11]
port 14 nsew signal tristate
flabel metal3 s 31600 7488 32000 7608 0 FreeSans 480 0 0 0 o_result_ring[12]
port 15 nsew signal tristate
flabel metal3 s 31600 5448 32000 5568 0 FreeSans 480 0 0 0 o_result_ring[13]
port 16 nsew signal tristate
flabel metal3 s 31600 8168 32000 8288 0 FreeSans 480 0 0 0 o_result_ring[14]
port 17 nsew signal tristate
flabel metal3 s 31600 8848 32000 8968 0 FreeSans 480 0 0 0 o_result_ring[15]
port 18 nsew signal tristate
flabel metal3 s 31600 9528 32000 9648 0 FreeSans 480 0 0 0 o_result_ring[16]
port 19 nsew signal tristate
flabel metal3 s 31600 10888 32000 11008 0 FreeSans 480 0 0 0 o_result_ring[17]
port 20 nsew signal tristate
flabel metal3 s 31600 10208 32000 10328 0 FreeSans 480 0 0 0 o_result_ring[18]
port 21 nsew signal tristate
flabel metal3 s 31600 15648 32000 15768 0 FreeSans 480 0 0 0 o_result_ring[19]
port 22 nsew signal tristate
flabel metal2 s 14186 0 14242 400 0 FreeSans 224 90 0 0 o_result_ring[1]
port 23 nsew signal tristate
flabel metal2 s 25134 19600 25190 20000 0 FreeSans 224 90 0 0 o_result_ring[20]
port 24 nsew signal tristate
flabel metal3 s 31600 11568 32000 11688 0 FreeSans 480 0 0 0 o_result_ring[21]
port 25 nsew signal tristate
flabel metal2 s 19982 19600 20038 20000 0 FreeSans 224 90 0 0 o_result_ring[22]
port 26 nsew signal tristate
flabel metal3 s 31600 12248 32000 12368 0 FreeSans 480 0 0 0 o_result_ring[23]
port 27 nsew signal tristate
flabel metal3 s 31600 12928 32000 13048 0 FreeSans 480 0 0 0 o_result_ring[24]
port 28 nsew signal tristate
flabel metal3 s 31600 13608 32000 13728 0 FreeSans 480 0 0 0 o_result_ring[25]
port 29 nsew signal tristate
flabel metal3 s 31600 14288 32000 14408 0 FreeSans 480 0 0 0 o_result_ring[26]
port 30 nsew signal tristate
flabel metal3 s 31600 14968 32000 15088 0 FreeSans 480 0 0 0 o_result_ring[27]
port 31 nsew signal tristate
flabel metal2 s 23202 19600 23258 20000 0 FreeSans 224 90 0 0 o_result_ring[28]
port 32 nsew signal tristate
flabel metal2 s 21914 19600 21970 20000 0 FreeSans 224 90 0 0 o_result_ring[29]
port 33 nsew signal tristate
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 o_result_ring[2]
port 34 nsew signal tristate
flabel metal2 s 21270 19600 21326 20000 0 FreeSans 224 90 0 0 o_result_ring[30]
port 35 nsew signal tristate
flabel metal2 s 20626 19600 20682 20000 0 FreeSans 224 90 0 0 o_result_ring[31]
port 36 nsew signal tristate
flabel metal2 s 24490 19600 24546 20000 0 FreeSans 224 90 0 0 o_result_ring[32]
port 37 nsew signal tristate
flabel metal2 s 22558 19600 22614 20000 0 FreeSans 224 90 0 0 o_result_ring[33]
port 38 nsew signal tristate
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 224 90 0 0 o_result_ring[34]
port 39 nsew signal tristate
flabel metal2 s 8390 19600 8446 20000 0 FreeSans 224 90 0 0 o_result_ring[35]
port 40 nsew signal tristate
flabel metal2 s 16118 19600 16174 20000 0 FreeSans 224 90 0 0 o_result_ring[36]
port 41 nsew signal tristate
flabel metal2 s 9034 19600 9090 20000 0 FreeSans 224 90 0 0 o_result_ring[37]
port 42 nsew signal tristate
flabel metal2 s 11610 19600 11666 20000 0 FreeSans 224 90 0 0 o_result_ring[38]
port 43 nsew signal tristate
flabel metal2 s 10322 19600 10378 20000 0 FreeSans 224 90 0 0 o_result_ring[39]
port 44 nsew signal tristate
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 o_result_ring[3]
port 45 nsew signal tristate
flabel metal2 s 9678 19600 9734 20000 0 FreeSans 224 90 0 0 o_result_ring[40]
port 46 nsew signal tristate
flabel metal2 s 12898 19600 12954 20000 0 FreeSans 224 90 0 0 o_result_ring[41]
port 47 nsew signal tristate
flabel metal3 s 0 12928 400 13048 0 FreeSans 480 0 0 0 o_result_ring[42]
port 48 nsew signal tristate
flabel metal2 s 10966 19600 11022 20000 0 FreeSans 224 90 0 0 o_result_ring[43]
port 49 nsew signal tristate
flabel metal2 s 12254 19600 12310 20000 0 FreeSans 224 90 0 0 o_result_ring[44]
port 50 nsew signal tristate
flabel metal2 s 15474 19600 15530 20000 0 FreeSans 224 90 0 0 o_result_ring[45]
port 51 nsew signal tristate
flabel metal2 s 14186 19600 14242 20000 0 FreeSans 224 90 0 0 o_result_ring[46]
port 52 nsew signal tristate
flabel metal2 s 16762 19600 16818 20000 0 FreeSans 224 90 0 0 o_result_ring[47]
port 53 nsew signal tristate
flabel metal2 s 18050 19600 18106 20000 0 FreeSans 224 90 0 0 o_result_ring[48]
port 54 nsew signal tristate
flabel metal2 s 23846 19600 23902 20000 0 FreeSans 224 90 0 0 o_result_ring[49]
port 55 nsew signal tristate
flabel metal2 s 18694 0 18750 400 0 FreeSans 224 90 0 0 o_result_ring[4]
port 56 nsew signal tristate
flabel metal2 s 19338 19600 19394 20000 0 FreeSans 224 90 0 0 o_result_ring[50]
port 57 nsew signal tristate
flabel metal2 s 18694 19600 18750 20000 0 FreeSans 224 90 0 0 o_result_ring[51]
port 58 nsew signal tristate
flabel metal2 s 19338 0 19394 400 0 FreeSans 224 90 0 0 o_result_ring[52]
port 59 nsew signal tristate
flabel metal2 s 17406 0 17462 400 0 FreeSans 224 90 0 0 o_result_ring[53]
port 60 nsew signal tristate
flabel metal2 s 14830 0 14886 400 0 FreeSans 224 90 0 0 o_result_ring[54]
port 61 nsew signal tristate
flabel metal2 s 14830 19600 14886 20000 0 FreeSans 224 90 0 0 o_result_ring[55]
port 62 nsew signal tristate
flabel metal2 s 13542 19600 13598 20000 0 FreeSans 224 90 0 0 o_result_ring[56]
port 63 nsew signal tristate
flabel metal3 s 0 10888 400 11008 0 FreeSans 480 0 0 0 o_result_ring[57]
port 64 nsew signal tristate
flabel metal3 s 0 10208 400 10328 0 FreeSans 480 0 0 0 o_result_ring[58]
port 65 nsew signal tristate
flabel metal3 s 0 9528 400 9648 0 FreeSans 480 0 0 0 o_result_ring[59]
port 66 nsew signal tristate
flabel metal2 s 19982 0 20038 400 0 FreeSans 224 90 0 0 o_result_ring[5]
port 67 nsew signal tristate
flabel metal2 s 12898 0 12954 400 0 FreeSans 224 90 0 0 o_result_ring[60]
port 68 nsew signal tristate
flabel metal3 s 0 8168 400 8288 0 FreeSans 480 0 0 0 o_result_ring[61]
port 69 nsew signal tristate
flabel metal2 s 9678 0 9734 400 0 FreeSans 224 90 0 0 o_result_ring[62]
port 70 nsew signal tristate
flabel metal2 s 12254 0 12310 400 0 FreeSans 224 90 0 0 o_result_ring[63]
port 71 nsew signal tristate
flabel metal2 s 18050 0 18106 400 0 FreeSans 224 90 0 0 o_result_ring[6]
port 72 nsew signal tristate
flabel metal2 s 22558 0 22614 400 0 FreeSans 224 90 0 0 o_result_ring[7]
port 73 nsew signal tristate
flabel metal2 s 21270 0 21326 400 0 FreeSans 224 90 0 0 o_result_ring[8]
port 74 nsew signal tristate
flabel metal3 s 31600 6128 32000 6248 0 FreeSans 480 0 0 0 o_result_ring[9]
port 75 nsew signal tristate
rlabel via1 16041 19040 16041 19040 0 VGND
rlabel metal1 15962 18496 15962 18496 0 VPWR
rlabel metal1 16284 3706 16284 3706 0 _000_
rlabel via1 14209 4046 14209 4046 0 _001_
rlabel metal1 15640 4522 15640 4522 0 _002_
rlabel metal1 13427 5746 13427 5746 0 _003_
rlabel metal1 11812 4046 11812 4046 0 _004_
rlabel metal2 8786 3774 8786 3774 0 _005_
rlabel metal1 8448 5066 8448 5066 0 _006_
rlabel via1 9701 5746 9701 5746 0 _007_
rlabel metal1 7590 6800 7590 6800 0 _008_
rlabel metal1 9246 5814 9246 5814 0 _009_
rlabel metal1 16238 3570 16238 3570 0 _010_
rlabel metal1 14398 3706 14398 3706 0 _011_
rlabel metal1 16514 5338 16514 5338 0 _012_
rlabel metal1 16330 4522 16330 4522 0 _013_
rlabel metal1 15410 4624 15410 4624 0 _014_
rlabel metal1 13202 5134 13202 5134 0 _015_
rlabel metal1 13340 5066 13340 5066 0 _016_
rlabel metal1 13478 4658 13478 4658 0 _017_
rlabel metal1 11362 4046 11362 4046 0 _018_
rlabel metal1 9798 4182 9798 4182 0 _019_
rlabel metal1 9936 3910 9936 3910 0 _020_
rlabel metal1 9246 3910 9246 3910 0 _021_
rlabel metal1 9798 6290 9798 6290 0 _022_
rlabel metal1 10028 4794 10028 4794 0 _023_
rlabel metal1 8050 5168 8050 5168 0 _024_
rlabel metal1 10028 6154 10028 6154 0 _025_
rlabel metal1 14352 13430 14352 13430 0 clknet_0_i_stop
rlabel metal2 15226 13634 15226 13634 0 clknet_0_net9
rlabel metal1 10258 8534 10258 8534 0 clknet_3_0__leaf_i_stop
rlabel metal1 8694 10608 8694 10608 0 clknet_3_0__leaf_net9
rlabel metal1 14490 5780 14490 5780 0 clknet_3_1__leaf_i_stop
rlabel metal1 13984 7310 13984 7310 0 clknet_3_1__leaf_net9
rlabel metal2 7774 11492 7774 11492 0 clknet_3_2__leaf_i_stop
rlabel metal1 7130 14314 7130 14314 0 clknet_3_2__leaf_net9
rlabel metal1 13846 12750 13846 12750 0 clknet_3_3__leaf_i_stop
rlabel metal1 15594 16048 15594 16048 0 clknet_3_3__leaf_net9
rlabel metal1 18078 6698 18078 6698 0 clknet_3_4__leaf_i_stop
rlabel metal1 24150 7480 24150 7480 0 clknet_3_4__leaf_net9
rlabel metal1 18929 9010 18929 9010 0 clknet_3_5__leaf_i_stop
rlabel metal1 21758 10132 21758 10132 0 clknet_3_5__leaf_net9
rlabel metal1 18308 14994 18308 14994 0 clknet_3_6__leaf_i_stop
rlabel metal1 19458 16626 19458 16626 0 clknet_3_6__leaf_net9
rlabel metal1 21850 15062 21850 15062 0 clknet_3_7__leaf_i_stop
rlabel metal1 24426 11662 24426 11662 0 clknet_3_7__leaf_net9
rlabel metal2 7774 415 7774 415 0 i_start
rlabel via3 15203 8364 15203 8364 0 i_stop
rlabel metal1 8798 5746 8798 5746 0 net1
rlabel metal1 21896 5338 21896 5338 0 net10
rlabel metal2 22494 5831 22494 5831 0 net100
rlabel metal1 24288 7310 24288 7310 0 net101
rlabel metal1 22724 5066 22724 5066 0 net103
rlabel metal1 21850 6392 21850 6392 0 net104
rlabel metal1 20516 9010 20516 9010 0 net106
rlabel metal1 23598 5814 23598 5814 0 net107
rlabel metal1 22903 7310 22903 7310 0 net108
rlabel metal2 21022 5083 21022 5083 0 net11
rlabel metal1 21666 6256 21666 6256 0 net110
rlabel metal2 21390 6528 21390 6528 0 net111
rlabel metal2 25530 8177 25530 8177 0 net112
rlabel metal1 23736 7310 23736 7310 0 net113
rlabel metal1 21114 8330 21114 8330 0 net115
rlabel via2 21942 8347 21942 8347 0 net116
rlabel metal1 24702 10098 24702 10098 0 net117
rlabel metal1 25576 9010 25576 9010 0 net119
rlabel metal2 19274 5474 19274 5474 0 net12
rlabel metal1 19090 8602 19090 8602 0 net120
rlabel metal1 23506 11186 23506 11186 0 net121
rlabel metal1 23230 8500 23230 8500 0 net123
rlabel metal1 25254 8976 25254 8976 0 net124
rlabel metal2 21390 9996 21390 9996 0 net125
rlabel metal1 25484 9690 25484 9690 0 net127
rlabel metal1 23041 9486 23041 9486 0 net128
rlabel metal1 24196 10642 24196 10642 0 net129
rlabel metal1 19918 5882 19918 5882 0 net13
rlabel metal1 20976 9010 20976 9010 0 net131
rlabel metal1 23363 10098 23363 10098 0 net132
rlabel metal2 21712 13124 21712 13124 0 net133
rlabel metal1 20562 10030 20562 10030 0 net135
rlabel metal1 23777 10506 23777 10506 0 net136
rlabel metal1 21528 13362 21528 13362 0 net137
rlabel metal1 20470 10506 20470 10506 0 net139
rlabel metal2 9338 7412 9338 7412 0 net14
rlabel metal1 19499 10166 19499 10166 0 net140
rlabel metal1 21666 13498 21666 13498 0 net141
rlabel metal1 21206 11798 21206 11798 0 net143
rlabel metal2 25162 11322 25162 11322 0 net144
rlabel metal1 21390 13226 21390 13226 0 net145
rlabel metal1 21022 12682 21022 12682 0 net147
rlabel metal2 19734 11492 19734 11492 0 net148
rlabel metal1 22540 16014 22540 16014 0 net149
rlabel metal2 9890 7548 9890 7548 0 net15
rlabel metal2 24702 11900 24702 11900 0 net151
rlabel metal1 23225 11662 23225 11662 0 net152
rlabel metal1 24242 13838 24242 13838 0 net153
rlabel via2 21942 15555 21942 15555 0 net155
rlabel metal1 19683 12682 19683 12682 0 net156
rlabel metal2 24610 15980 24610 15980 0 net157
rlabel metal1 23869 14314 23869 14314 0 net159
rlabel metal1 8694 6863 8694 6863 0 net16
rlabel metal1 24651 12342 24651 12342 0 net160
rlabel metal1 21942 15980 21942 15980 0 net161
rlabel metal2 24380 12750 24380 12750 0 net163
rlabel metal2 23690 13039 23690 13039 0 net164
rlabel metal1 23782 15538 23782 15538 0 net165
rlabel metal2 24610 13889 24610 13889 0 net167
rlabel metal1 24283 13362 24283 13362 0 net168
rlabel metal1 22954 15946 22954 15946 0 net169
rlabel metal1 19550 6800 19550 6800 0 net17
rlabel metal1 21160 16014 21160 16014 0 net171
rlabel metal1 22903 13838 22903 13838 0 net172
rlabel metal1 19274 17102 19274 17102 0 net173
rlabel metal1 23598 14960 23598 14960 0 net175
rlabel metal1 22903 14518 22903 14518 0 net176
rlabel metal1 19090 16626 19090 16626 0 net177
rlabel metal1 21620 17306 21620 17306 0 net179
rlabel metal1 6670 8976 6670 8976 0 net18
rlabel metal1 22581 14858 22581 14858 0 net180
rlabel metal1 20516 15334 20516 15334 0 net181
rlabel metal2 20010 16218 20010 16218 0 net183
rlabel metal1 23322 14994 23322 14994 0 net184
rlabel metal1 20746 13872 20746 13872 0 net185
rlabel metal1 19412 15538 19412 15538 0 net187
rlabel metal1 19637 14926 19637 14926 0 net188
rlabel metal1 16556 16014 16556 16014 0 net189
rlabel metal1 7222 9622 7222 9622 0 net19
rlabel metal1 19136 14450 19136 14450 0 net191
rlabel metal1 19959 13430 19959 13430 0 net192
rlabel metal1 14030 16592 14030 16592 0 net193
rlabel metal1 17434 14450 17434 14450 0 net195
rlabel metal1 17107 14858 17107 14858 0 net196
rlabel metal1 13662 15946 13662 15946 0 net197
rlabel metal1 16238 15674 16238 15674 0 net199
rlabel viali 8522 11662 8522 11662 0 net2
rlabel metal1 8142 10064 8142 10064 0 net20
rlabel via1 17981 13362 17981 13362 0 net200
rlabel metal1 13432 16626 13432 16626 0 net201
rlabel metal1 15502 15504 15502 15504 0 net203
rlabel metal1 15543 14858 15543 14858 0 net204
rlabel metal2 14030 16660 14030 16660 0 net205
rlabel metal1 13432 14994 13432 14994 0 net207
rlabel metal1 14770 13770 14770 13770 0 net208
rlabel metal1 11454 16014 11454 16014 0 net209
rlabel metal1 8786 10166 8786 10166 0 net21
rlabel metal2 12650 15844 12650 15844 0 net211
rlabel via1 14669 14450 14669 14450 0 net212
rlabel metal1 7958 14960 7958 14960 0 net213
rlabel metal1 9890 14824 9890 14824 0 net215
rlabel metal1 15011 14858 15011 14858 0 net216
rlabel metal1 7682 14450 7682 14450 0 net217
rlabel metal1 8878 14960 8878 14960 0 net219
rlabel metal1 11178 9520 11178 9520 0 net22
rlabel metal1 10083 15980 10083 15980 0 net220
rlabel metal2 7958 13668 7958 13668 0 net221
rlabel metal2 8050 15164 8050 15164 0 net223
rlabel metal1 9430 14824 9430 14824 0 net224
rlabel metal2 8096 13362 8096 13362 0 net225
rlabel metal1 7222 13906 7222 13906 0 net227
rlabel metal1 8632 13770 8632 13770 0 net228
rlabel metal1 8004 13362 8004 13362 0 net229
rlabel metal2 11914 9282 11914 9282 0 net23
rlabel metal1 7636 13362 7636 13362 0 net231
rlabel via1 12277 13430 12277 13430 0 net232
rlabel metal1 12098 15572 12098 15572 0 net233
rlabel metal1 8096 12750 8096 12750 0 net235
rlabel metal1 9618 12682 9618 12682 0 net236
rlabel metal2 14306 14620 14306 14620 0 net237
rlabel metal1 9982 13328 9982 13328 0 net239
rlabel metal1 13524 8602 13524 8602 0 net24
rlabel metal1 9966 11594 9966 11594 0 net240
rlabel metal1 13110 13804 13110 13804 0 net241
rlabel metal2 13156 13668 13156 13668 0 net243
rlabel metal1 11086 11730 11086 11730 0 net244
rlabel metal1 16238 13804 16238 13804 0 net245
rlabel metal1 13248 14382 13248 14382 0 net247
rlabel metal2 13018 12920 13018 12920 0 net248
rlabel metal1 17296 12954 17296 12954 0 net249
rlabel metal1 15272 9010 15272 9010 0 net25
rlabel metal2 13294 12444 13294 12444 0 net251
rlabel metal1 13018 12104 13018 12104 0 net252
rlabel metal1 16422 11764 16422 11764 0 net253
rlabel metal2 13846 11900 13846 11900 0 net255
rlabel metal1 16320 13362 16320 13362 0 net256
rlabel metal1 19366 11152 19366 11152 0 net257
rlabel metal1 14766 11798 14766 11798 0 net259
rlabel metal1 15778 9044 15778 9044 0 net26
rlabel metal1 17234 12682 17234 12682 0 net260
rlabel metal1 16422 9486 16422 9486 0 net261
rlabel metal1 15548 11186 15548 11186 0 net263
rlabel metal1 18032 11662 18032 11662 0 net264
rlabel metal1 17664 9146 17664 9146 0 net265
rlabel metal1 18446 11152 18446 11152 0 net267
rlabel metal1 18211 10506 18211 10506 0 net268
rlabel metal1 16560 9622 16560 9622 0 net269
rlabel metal1 18170 11186 18170 11186 0 net27
rlabel metal1 16238 9010 16238 9010 0 net271
rlabel metal1 18073 10098 18073 10098 0 net272
rlabel metal1 14030 10132 14030 10132 0 net273
rlabel metal1 13570 9418 13570 9418 0 net275
rlabel metal1 18032 8602 18032 8602 0 net276
rlabel metal1 13294 8942 13294 8942 0 net277
rlabel metal1 12374 9520 12374 9520 0 net279
rlabel metal1 15640 6970 15640 6970 0 net28
rlabel metal1 15992 8330 15992 8330 0 net280
rlabel metal1 12466 10132 12466 10132 0 net281
rlabel metal1 13524 8534 13524 8534 0 net283
rlabel metal1 13606 9010 13606 9010 0 net284
rlabel metal1 10442 9452 10442 9452 0 net285
rlabel metal1 11040 9486 11040 9486 0 net287
rlabel metal2 13386 10370 13386 10370 0 net288
rlabel metal1 10258 8806 10258 8806 0 net289
rlabel metal1 15686 11220 15686 11220 0 net29
rlabel metal1 9154 10098 9154 10098 0 net291
rlabel metal1 11944 10506 11944 10506 0 net292
rlabel metal1 8464 10098 8464 10098 0 net293
rlabel metal1 8004 10098 8004 10098 0 net295
rlabel via1 11550 10506 11550 10506 0 net296
rlabel metal1 7038 10064 7038 10064 0 net297
rlabel metal1 7728 9690 7728 9690 0 net299
rlabel metal1 7623 11662 7623 11662 0 net3
rlabel metal1 14766 11866 14766 11866 0 net30
rlabel metal1 9848 10098 9848 10098 0 net300
rlabel metal1 7728 8398 7728 8398 0 net301
rlabel metal1 6532 9010 6532 9010 0 net303
rlabel via1 9802 9418 9802 9418 0 net304
rlabel metal1 7774 7990 7774 7990 0 net305
rlabel metal2 8878 7310 8878 7310 0 net307
rlabel metal1 11883 8296 11883 8296 0 net308
rlabel metal2 7176 7310 7176 7310 0 net309
rlabel metal1 13478 11662 13478 11662 0 net31
rlabel metal1 9062 7344 9062 7344 0 net311
rlabel metal1 9894 8330 9894 8330 0 net312
rlabel metal2 10396 6426 10396 6426 0 net314
rlabel metal1 9292 6834 9292 6834 0 net315
rlabel metal2 12650 7514 12650 7514 0 net316
rlabel metal1 10396 6426 10396 6426 0 net317
rlabel metal1 8878 6970 8878 6970 0 net318
rlabel metal1 11224 6834 11224 6834 0 net319
rlabel metal1 14812 14042 14812 14042 0 net32
rlabel metal2 13754 7786 13754 7786 0 net320
rlabel metal1 12719 6358 12719 6358 0 net321
rlabel metal1 10856 6902 10856 6902 0 net322
rlabel metal1 12558 8568 12558 8568 0 net323
rlabel metal1 15460 7920 15460 7920 0 net324
rlabel via1 16694 7310 16694 7310 0 net325
rlabel metal1 13478 6154 13478 6154 0 net326
rlabel metal1 15088 7310 15088 7310 0 net327
rlabel metal1 15778 7820 15778 7820 0 net328
rlabel metal1 14260 7242 14260 7242 0 net329
rlabel metal1 12558 13906 12558 13906 0 net33
rlabel metal1 15824 7514 15824 7514 0 net330
rlabel metal1 15870 6188 15870 6188 0 net331
rlabel metal1 20838 7310 20838 7310 0 net332
rlabel metal1 19504 7310 19504 7310 0 net333
rlabel metal1 21390 7310 21390 7310 0 net334
rlabel metal2 19090 6630 19090 6630 0 net335
rlabel metal1 19734 6970 19734 6970 0 net336
rlabel metal1 19872 6086 19872 6086 0 net337
rlabel metal2 25346 6698 25346 6698 0 net338
rlabel metal2 22126 5202 22126 5202 0 net339
rlabel metal1 11086 13974 11086 13974 0 net34
rlabel metal1 20562 5780 20562 5780 0 net340
rlabel metal2 26174 6732 26174 6732 0 net341
rlabel metal1 21114 5134 21114 5134 0 net342
rlabel metal1 20654 4522 20654 4522 0 net343
rlabel metal1 21068 4998 21068 4998 0 net344
rlabel metal1 24564 7310 24564 7310 0 net345
rlabel metal1 20704 8398 20704 8398 0 net346
rlabel metal1 25484 7854 25484 7854 0 net347
rlabel metal2 21206 8602 21206 8602 0 net348
rlabel metal2 22126 7038 22126 7038 0 net349
rlabel metal1 9798 13396 9798 13396 0 net35
rlabel metal1 25070 7276 25070 7276 0 net350
rlabel metal1 22034 6154 22034 6154 0 net351
rlabel metal1 26312 9486 26312 9486 0 net352
rlabel metal2 24702 9792 24702 9792 0 net353
rlabel metal2 25438 8636 25438 8636 0 net354
rlabel metal1 21988 9078 21988 9078 0 net355
rlabel metal2 23414 9350 23414 9350 0 net356
rlabel metal2 23046 8160 23046 8160 0 net357
rlabel metal1 24472 9690 24472 9690 0 net358
rlabel metal1 19826 10608 19826 10608 0 net359
rlabel metal1 8510 12682 8510 12682 0 net36
rlabel metal2 20746 10846 20746 10846 0 net360
rlabel metal1 21160 10098 21160 10098 0 net361
rlabel metal1 20930 11220 20930 11220 0 net362
rlabel metal1 24610 10778 24610 10778 0 net363
rlabel metal1 21390 10234 21390 10234 0 net364
rlabel metal2 24886 10880 24886 10880 0 net365
rlabel metal1 26082 11764 26082 11764 0 net366
rlabel metal1 25254 12274 25254 12274 0 net367
rlabel metal1 20654 11628 20654 11628 0 net368
rlabel metal1 26266 12784 26266 12784 0 net369
rlabel metal1 7774 13396 7774 13396 0 net37
rlabel metal1 24426 12716 24426 12716 0 net370
rlabel metal1 21574 12614 21574 12614 0 net371
rlabel metal2 24518 13039 24518 13039 0 net372
rlabel metal1 26266 12308 26266 12308 0 net373
rlabel metal2 24794 13362 24794 13362 0 net374
rlabel metal1 21298 13872 21298 13872 0 net375
rlabel metal1 24518 15538 24518 15538 0 net376
rlabel metal1 26082 13872 26082 13872 0 net377
rlabel metal2 25346 14722 25346 14722 0 net378
rlabel metal2 26174 14127 26174 14127 0 net379
rlabel metal2 10166 15385 10166 15385 0 net38
rlabel metal1 24104 16218 24104 16218 0 net380
rlabel metal1 23506 15538 23506 15538 0 net381
rlabel metal1 24242 16014 24242 16014 0 net382
rlabel metal1 21758 17136 21758 17136 0 net383
rlabel metal2 24058 15096 24058 15096 0 net384
rlabel metal1 20976 16218 20976 16218 0 net385
rlabel metal2 20378 16677 20378 16677 0 net386
rlabel metal1 20654 16048 20654 16048 0 net387
rlabel metal1 19964 15674 19964 15674 0 net388
rlabel metal1 21850 16626 21850 16626 0 net389
rlabel metal1 16238 7344 16238 7344 0 net39
rlabel metal1 21390 13804 21390 13804 0 net390
rlabel metal2 21758 14450 21758 14450 0 net391
rlabel metal1 19734 16218 19734 16218 0 net392
rlabel metal1 20056 15946 20056 15946 0 net393
rlabel metal1 18032 13838 18032 13838 0 net394
rlabel via1 16698 15537 16698 15537 0 net395
rlabel metal2 19458 14892 19458 14892 0 net396
rlabel metal1 12006 13804 12006 13804 0 net397
rlabel metal1 18124 14042 18124 14042 0 net398
rlabel metal1 18354 14586 18354 14586 0 net399
rlabel metal1 8860 11662 8860 11662 0 net4
rlabel metal1 7452 14042 7452 14042 0 net40
rlabel metal1 17848 14246 17848 14246 0 net400
rlabel metal1 14858 16660 14858 16660 0 net401
rlabel metal1 11914 17068 11914 17068 0 net402
rlabel metal1 14674 16014 14674 16014 0 net403
rlabel metal2 13386 16218 13386 16218 0 net404
rlabel metal2 13846 16932 13846 16932 0 net405
rlabel metal1 13662 15674 13662 15674 0 net406
rlabel metal1 13478 16218 13478 16218 0 net407
rlabel metal1 8050 14892 8050 14892 0 net408
rlabel metal1 9292 15674 9292 15674 0 net409
rlabel metal1 8740 14926 8740 14926 0 net41
rlabel metal1 9936 15674 9936 15674 0 net410
rlabel metal1 12098 16218 12098 16218 0 net411
rlabel metal1 8050 14042 8050 14042 0 net412
rlabel metal1 8602 14790 8602 14790 0 net413
rlabel metal2 10994 16354 10994 16354 0 net414
rlabel metal1 7636 12274 7636 12274 0 net415
rlabel metal1 8326 13362 8326 13362 0 net416
rlabel metal1 9154 14246 9154 14246 0 net417
rlabel metal2 12926 14603 12926 14603 0 net418
rlabel metal1 8510 13838 8510 13838 0 net419
rlabel metal1 10580 15538 10580 15538 0 net42
rlabel metal1 8188 13294 8188 13294 0 net420
rlabel metal2 7590 13362 7590 13362 0 net421
rlabel metal1 11730 13396 11730 13396 0 net422
rlabel metal1 13754 14416 13754 14416 0 net423
rlabel metal2 10534 14178 10534 14178 0 net424
rlabel metal2 13846 13838 13846 13838 0 net425
rlabel metal2 11546 12716 11546 12716 0 net426
rlabel metal1 10948 14042 10948 14042 0 net427
rlabel metal2 11592 13260 11592 13260 0 net428
rlabel metal1 17158 13872 17158 13872 0 net429
rlabel metal2 12834 16218 12834 16218 0 net43
rlabel metal1 14490 11730 14490 11730 0 net430
rlabel metal1 14858 13498 14858 13498 0 net431
rlabel metal1 19274 11220 19274 11220 0 net432
rlabel metal1 15824 9894 15824 9894 0 net433
rlabel metal1 13846 11866 13846 11866 0 net434
rlabel metal2 16790 10608 16790 10608 0 net435
rlabel metal2 19366 10914 19366 10914 0 net436
rlabel metal1 16422 10132 16422 10132 0 net437
rlabel metal1 16146 10608 16146 10608 0 net438
rlabel metal1 15410 9554 15410 9554 0 net439
rlabel metal1 13202 15062 13202 15062 0 net44
rlabel metal2 18078 9316 18078 9316 0 net440
rlabel metal2 18262 11543 18262 11543 0 net441
rlabel via2 17986 9605 17986 9605 0 net442
rlabel metal1 11454 9452 11454 9452 0 net443
rlabel metal2 12926 9622 12926 9622 0 net444
rlabel metal1 14030 9520 14030 9520 0 net445
rlabel metal1 12006 9520 12006 9520 0 net446
rlabel metal1 13892 10234 13892 10234 0 net447
rlabel metal1 12742 9418 12742 9418 0 net448
rlabel metal1 13708 10234 13708 10234 0 net449
rlabel metal1 15318 15572 15318 15572 0 net45
rlabel metal1 9798 10574 9798 10574 0 net450
rlabel metal1 9246 11186 9246 11186 0 net451
rlabel metal1 9982 10642 9982 10642 0 net452
rlabel metal1 10626 9044 10626 9044 0 net453
rlabel metal2 10442 10132 10442 10132 0 net454
rlabel metal1 8970 10234 8970 10234 0 net455
rlabel metal1 8740 10778 8740 10778 0 net456
rlabel metal2 10902 8772 10902 8772 0 net457
rlabel metal1 8464 7922 8464 7922 0 net458
rlabel metal2 8510 8602 8510 8602 0 net459
rlabel metal1 15962 15980 15962 15980 0 net46
rlabel metal1 8648 7922 8648 7922 0 net460
rlabel metal2 6210 10370 6210 10370 0 net461
rlabel metal2 6670 9520 6670 9520 0 net462
rlabel metal1 8372 11050 8372 11050 0 net463
rlabel metal1 8142 6970 8142 6970 0 net464
rlabel metal1 8786 6698 8786 6698 0 net465
rlabel metal2 7038 7463 7038 7463 0 net466
rlabel metal1 13018 7820 13018 7820 0 net467
rlabel metal1 10120 6086 10120 6086 0 net469
rlabel metal1 17710 14484 17710 14484 0 net47
rlabel metal1 12640 6834 12640 6834 0 net470
rlabel metal1 10534 4794 10534 4794 0 net471
rlabel metal1 9568 5542 9568 5542 0 net472
rlabel metal1 9522 4250 9522 4250 0 net473
rlabel metal1 12604 4590 12604 4590 0 net474
rlabel metal1 13156 4794 13156 4794 0 net475
rlabel metal1 16836 5066 16836 5066 0 net476
rlabel metal1 14720 3502 14720 3502 0 net477
rlabel metal1 16146 3434 16146 3434 0 net478
rlabel metal1 8786 5882 8786 5882 0 net479
rlabel metal1 19366 14484 19366 14484 0 net48
rlabel metal2 12374 6290 12374 6290 0 net480
rlabel metal1 15502 5134 15502 5134 0 net481
rlabel metal1 11362 6863 11362 6863 0 net482
rlabel metal2 14996 6460 14996 6460 0 net483
rlabel metal1 15272 5134 15272 5134 0 net484
rlabel metal1 11684 6970 11684 6970 0 net485
rlabel metal1 15410 5338 15410 5338 0 net486
rlabel metal1 19734 8398 19734 8398 0 net487
rlabel metal2 19458 6477 19458 6477 0 net488
rlabel metal1 19274 7344 19274 7344 0 net489
rlabel metal1 19182 15504 19182 15504 0 net49
rlabel metal1 20102 6868 20102 6868 0 net490
rlabel metal1 18170 6256 18170 6256 0 net491
rlabel metal1 15916 6766 15916 6766 0 net492
rlabel metal1 18032 6222 18032 6222 0 net493
rlabel metal1 20700 4454 20700 4454 0 net494
rlabel metal1 20746 4692 20746 4692 0 net495
rlabel metal2 20102 4896 20102 4896 0 net496
rlabel metal2 24978 7004 24978 7004 0 net497
rlabel metal1 20102 5746 20102 5746 0 net498
rlabel metal1 20056 5338 20056 5338 0 net499
rlabel metal1 8267 11662 8267 11662 0 net5
rlabel metal1 16146 4692 16146 4692 0 net50
rlabel metal1 20194 5542 20194 5542 0 net500
rlabel metal1 26542 8398 26542 8398 0 net501
rlabel metal2 21482 5916 21482 5916 0 net502
rlabel metal1 23276 6426 23276 6426 0 net503
rlabel metal1 22310 5780 22310 5780 0 net504
rlabel metal1 24380 6834 24380 6834 0 net505
rlabel metal1 23460 5338 23460 5338 0 net506
rlabel metal1 26036 8262 26036 8262 0 net507
rlabel metal1 26818 9010 26818 9010 0 net508
rlabel metal1 22080 9146 22080 9146 0 net509
rlabel metal1 19826 16048 19826 16048 0 net51
rlabel metal2 23598 6902 23598 6902 0 net510
rlabel metal1 26220 9690 26220 9690 0 net511
rlabel metal1 25714 10098 25714 10098 0 net512
rlabel metal2 25990 9554 25990 9554 0 net513
rlabel metal1 25438 8602 25438 8602 0 net514
rlabel metal1 25392 10982 25392 10982 0 net515
rlabel metal1 21574 10098 21574 10098 0 net516
rlabel metal1 23874 11186 23874 11186 0 net517
rlabel metal1 21574 11560 21574 11560 0 net518
rlabel metal1 21896 10574 21896 10574 0 net519
rlabel metal1 22034 16048 22034 16048 0 net52
rlabel metal2 21114 9282 21114 9282 0 net520
rlabel metal2 20930 10472 20930 10472 0 net521
rlabel metal1 19826 11220 19826 11220 0 net522
rlabel metal1 21298 12716 21298 12716 0 net523
rlabel metal1 21298 11662 21298 11662 0 net524
rlabel metal2 22034 13600 22034 13600 0 net525
rlabel metal1 20746 11866 20746 11866 0 net526
rlabel metal1 20792 11050 20792 11050 0 net527
rlabel metal2 20562 11968 20562 11968 0 net528
rlabel metal1 26036 12274 26036 12274 0 net529
rlabel metal2 22494 16320 22494 16320 0 net53
rlabel metal1 24242 14416 24242 14416 0 net530
rlabel metal1 25806 12750 25806 12750 0 net531
rlabel metal2 24610 14756 24610 14756 0 net532
rlabel metal2 20470 14025 20470 14025 0 net533
rlabel metal1 24748 12954 24748 12954 0 net534
rlabel metal1 21643 13974 21643 13974 0 net535
rlabel metal2 26634 14858 26634 14858 0 net536
rlabel metal2 21574 16847 21574 16847 0 net537
rlabel metal1 23874 15674 23874 15674 0 net538
rlabel metal2 24150 15742 24150 15742 0 net539
rlabel metal2 20930 15657 20930 15657 0 net54
rlabel metal1 22586 17102 22586 17102 0 net540
rlabel metal4 21988 14552 21988 14552 0 net541
rlabel metal1 22954 17000 22954 17000 0 net542
rlabel metal2 21482 15844 21482 15844 0 net543
rlabel metal1 21344 16218 21344 16218 0 net544
rlabel metal1 22954 16762 22954 16762 0 net545
rlabel metal1 20562 15504 20562 15504 0 net546
rlabel metal2 23966 16184 23966 16184 0 net547
rlabel metal2 22126 16728 22126 16728 0 net548
rlabel metal1 21758 16694 21758 16694 0 net549
rlabel metal1 24794 13464 24794 13464 0 net55
rlabel metal1 17342 16014 17342 16014 0 net550
rlabel metal1 17526 15538 17526 15538 0 net551
rlabel metal1 18262 15981 18262 15981 0 net552
rlabel metal1 16882 14416 16882 14416 0 net553
rlabel metal1 20010 14518 20010 14518 0 net554
rlabel metal1 19964 14042 19964 14042 0 net555
rlabel metal1 19826 14246 19826 14246 0 net556
rlabel metal1 12650 13838 12650 13838 0 net557
rlabel metal1 13018 14892 13018 14892 0 net558
rlabel metal1 17250 14484 17250 14484 0 net559
rlabel metal1 24150 12784 24150 12784 0 net56
rlabel metal1 13846 16014 13846 16014 0 net560
rlabel metal1 14306 15538 14306 15538 0 net561
rlabel metal1 15226 15674 15226 15674 0 net562
rlabel metal1 14490 15674 14490 15674 0 net563
rlabel metal1 9706 16048 9706 16048 0 net564
rlabel metal1 11362 17102 11362 17102 0 net565
rlabel metal1 11270 15606 11270 15606 0 net566
rlabel metal1 10534 14892 10534 14892 0 net567
rlabel metal1 12742 17136 12742 17136 0 net568
rlabel metal2 9614 15198 9614 15198 0 net569
rlabel metal2 23322 14773 23322 14773 0 net57
rlabel metal2 11362 16966 11362 16966 0 net570
rlabel metal1 12190 16014 12190 16014 0 net571
rlabel metal1 7682 13702 7682 13702 0 net572
rlabel metal1 9890 15606 9890 15606 0 net573
rlabel metal1 9798 12308 9798 12308 0 net574
rlabel metal2 9154 14892 9154 14892 0 net575
rlabel metal1 7958 13974 7958 13974 0 net576
rlabel metal1 9660 14586 9660 14586 0 net577
rlabel metal1 10534 12274 10534 12274 0 net578
rlabel metal1 10994 13226 10994 13226 0 net579
rlabel metal1 24748 12750 24748 12750 0 net58
rlabel metal1 9154 13391 9154 13391 0 net580
rlabel metal1 10810 12886 10810 12886 0 net581
rlabel metal1 10580 13498 10580 13498 0 net582
rlabel metal1 9752 12410 9752 12410 0 net583
rlabel metal2 13294 14892 13294 14892 0 net584
rlabel metal1 16330 14416 16330 14416 0 net585
rlabel metal1 14306 12303 14306 12303 0 net586
rlabel metal2 12926 12444 12926 12444 0 net587
rlabel metal1 14582 12274 14582 12274 0 net588
rlabel metal1 16422 13838 16422 13838 0 net589
rlabel metal1 24886 11628 24886 11628 0 net59
rlabel metal1 13248 12070 13248 12070 0 net590
rlabel metal1 16330 13906 16330 13906 0 net591
rlabel metal1 18952 10574 18952 10574 0 net592
rlabel metal2 19458 11475 19458 11475 0 net593
rlabel metal1 15456 11866 15456 11866 0 net594
rlabel metal1 16514 10574 16514 10574 0 net595
rlabel metal2 16882 10948 16882 10948 0 net596
rlabel metal1 16008 11322 16008 11322 0 net597
rlabel metal1 15962 10778 15962 10778 0 net598
rlabel metal1 15640 9010 15640 9010 0 net599
rlabel metal1 8487 11526 8487 11526 0 net6
rlabel metal2 20930 12716 20930 12716 0 net60
rlabel metal1 12926 9486 12926 9486 0 net600
rlabel metal1 15456 10234 15456 10234 0 net601
rlabel metal1 13938 8398 13938 8398 0 net602
rlabel metal1 14306 9690 14306 9690 0 net603
rlabel metal1 14076 9418 14076 9418 0 net604
rlabel metal2 13938 9792 13938 9792 0 net605
rlabel metal1 10120 10574 10120 10574 0 net606
rlabel metal1 10810 9656 10810 9656 0 net607
rlabel metal2 12558 10676 12558 10676 0 net608
rlabel metal1 10258 9078 10258 9078 0 net609
rlabel metal2 12742 6834 12742 6834 0 net61
rlabel metal1 10994 11220 10994 11220 0 net610
rlabel metal1 11224 9622 11224 9622 0 net611
rlabel metal2 9890 10336 9890 10336 0 net612
rlabel metal1 6670 9486 6670 9486 0 net613
rlabel metal1 6762 9078 6762 9078 0 net614
rlabel metal1 8326 9559 8326 9559 0 net615
rlabel metal1 8602 7514 8602 7514 0 net616
rlabel metal1 8878 9010 8878 9010 0 net617
rlabel metal1 7406 9690 7406 9690 0 net618
rlabel metal1 8832 8602 8832 8602 0 net619
rlabel metal1 20194 11254 20194 11254 0 net62
rlabel metal1 10626 7990 10626 7990 0 net620
rlabel metal1 10672 6154 10672 6154 0 net621
rlabel via1 7678 7310 7678 7310 0 net622
rlabel metal1 9016 7922 9016 7922 0 net623
rlabel metal1 8188 7310 8188 7310 0 net624
rlabel metal1 9384 7514 9384 7514 0 net625
rlabel metal1 7774 7242 7774 7242 0 net627
rlabel metal1 11316 5678 11316 5678 0 net628
rlabel metal1 11587 6154 11587 6154 0 net629
rlabel metal1 20654 10608 20654 10608 0 net63
rlabel metal1 11040 7514 11040 7514 0 net630
rlabel metal1 10120 6970 10120 6970 0 net631
rlabel metal1 10994 4454 10994 4454 0 net632
rlabel metal2 11454 7582 11454 7582 0 net633
rlabel metal1 18722 8432 18722 8432 0 net634
rlabel metal1 16698 6868 16698 6868 0 net635
rlabel metal1 15962 7310 15962 7310 0 net636
rlabel metal1 18446 6154 18446 6154 0 net637
rlabel metal1 17894 6188 17894 6188 0 net638
rlabel metal1 16744 7242 16744 7242 0 net639
rlabel metal1 20746 10064 20746 10064 0 net64
rlabel metal1 18216 6426 18216 6426 0 net640
rlabel metal1 19090 5270 19090 5270 0 net641
rlabel metal1 19918 5168 19918 5168 0 net642
rlabel metal1 19458 6256 19458 6256 0 net643
rlabel metal1 20746 4998 20746 4998 0 net644
rlabel metal1 20470 5100 20470 5100 0 net645
rlabel metal1 20424 6630 20424 6630 0 net646
rlabel metal2 20562 5117 20562 5117 0 net647
rlabel metal1 25208 6970 25208 6970 0 net648
rlabel metal1 23230 5746 23230 5746 0 net649
rlabel viali 21118 9010 21118 9010 0 net65
rlabel metal1 24426 8432 24426 8432 0 net650
rlabel metal1 21666 5032 21666 5032 0 net651
rlabel via2 21482 5355 21482 5355 0 net652
rlabel metal1 23046 5882 23046 5882 0 net653
rlabel metal2 24886 6630 24886 6630 0 net654
rlabel metal2 19458 8942 19458 8942 0 net655
rlabel metal1 24794 9588 24794 9588 0 net656
rlabel metal2 21758 7072 21758 7072 0 net657
rlabel metal1 20746 9486 20746 9486 0 net658
rlabel metal2 21942 6375 21942 6375 0 net659
rlabel metal1 25116 9690 25116 9690 0 net66
rlabel metal1 20746 8330 20746 8330 0 net660
rlabel metal2 21666 6035 21666 6035 0 net661
rlabel metal1 25300 10778 25300 10778 0 net662
rlabel metal2 21298 9180 21298 9180 0 net663
rlabel metal1 24380 9486 24380 9486 0 net664
rlabel metal1 23690 10574 23690 10574 0 net665
rlabel metal2 24334 10778 24334 10778 0 net666
rlabel metal2 25254 9248 25254 9248 0 net667
rlabel metal1 24150 10778 24150 10778 0 net668
rlabel metal1 25438 11730 25438 11730 0 net669
rlabel metal2 23046 8602 23046 8602 0 net67
rlabel metal1 24610 11594 24610 11594 0 net670
rlabel metal1 24656 10574 24656 10574 0 net671
rlabel metal1 21712 13362 21712 13362 0 net672
rlabel metal1 21482 11798 21482 11798 0 net673
rlabel metal1 20838 10506 20838 10506 0 net674
rlabel metal1 21022 12614 21022 12614 0 net675
rlabel metal1 20562 12750 20562 12750 0 net676
rlabel metal2 22034 14943 22034 14943 0 net677
rlabel metal1 21022 14484 21022 14484 0 net678
rlabel metal1 24794 13804 24794 13804 0 net679
rlabel metal1 25944 9010 25944 9010 0 net68
rlabel metal1 23184 13770 23184 13770 0 net680
rlabel metal2 24794 12070 24794 12070 0 net681
rlabel metal4 23276 14144 23276 14144 0 net682
rlabel metal1 25898 14484 25898 14484 0 net683
rlabel metal1 24702 14416 24702 14416 0 net684
rlabel metal1 25576 13974 25576 13974 0 net685
rlabel metal2 26358 14654 26358 14654 0 net686
rlabel via2 24794 14909 24794 14909 0 net687
rlabel metal1 24426 12818 24426 12818 0 net688
rlabel via2 23322 16235 23322 16235 0 net689
rlabel metal1 20884 8398 20884 8398 0 net69
rlabel metal2 24978 16388 24978 16388 0 net690
rlabel metal2 21482 16932 21482 16932 0 net691
rlabel metal1 20516 16626 20516 16626 0 net692
rlabel metal1 22678 15606 22678 15606 0 net693
rlabel metal1 23230 16660 23230 16660 0 net694
rlabel metal1 23046 15130 23046 15130 0 net695
rlabel metal2 23322 17000 23322 17000 0 net696
rlabel metal1 20838 14042 20838 14042 0 net697
rlabel metal1 18906 15538 18906 15538 0 net698
rlabel metal1 19642 16014 19642 16014 0 net699
rlabel metal1 8372 12818 8372 12818 0 net7
rlabel metal1 24104 7310 24104 7310 0 net70
rlabel metal1 18262 14926 18262 14926 0 net700
rlabel metal1 19734 15572 19734 15572 0 net701
rlabel metal1 19136 15674 19136 15674 0 net702
rlabel metal2 19826 15878 19826 15878 0 net703
rlabel metal1 16100 16626 16100 16626 0 net704
rlabel metal1 14444 14586 14444 14586 0 net705
rlabel metal1 16330 15504 16330 15504 0 net706
rlabel metal1 14214 16626 14214 16626 0 net707
rlabel metal2 18354 14076 18354 14076 0 net708
rlabel metal1 16054 15878 16054 15878 0 net709
rlabel metal1 24242 6426 24242 6426 0 net71
rlabel metal1 18446 13940 18446 13940 0 net710
rlabel metal1 15226 16694 15226 16694 0 net711
rlabel metal2 9982 14977 9982 14977 0 net712
rlabel metal2 13110 16218 13110 16218 0 net713
rlabel metal2 11086 16898 11086 16898 0 net714
rlabel metal2 11408 15538 11408 15538 0 net715
rlabel metal2 12742 15504 12742 15504 0 net716
rlabel metal1 12466 16592 12466 16592 0 net717
rlabel metal1 7498 14518 7498 14518 0 net718
rlabel metal1 8004 14518 8004 14518 0 net719
rlabel metal1 9522 6868 9522 6868 0 net72
rlabel metal1 10216 15538 10216 15538 0 net720
rlabel metal1 7866 13906 7866 13906 0 net721
rlabel metal1 9154 14994 9154 14994 0 net722
rlabel metal2 7958 15674 7958 15674 0 net723
rlabel metal2 9844 15130 9844 15130 0 net724
rlabel metal1 8970 11764 8970 11764 0 net725
rlabel metal2 12466 14535 12466 14535 0 net726
rlabel metal1 7682 12784 7682 12784 0 net727
rlabel metal2 10166 13634 10166 13634 0 net728
rlabel metal1 8878 13294 8878 13294 0 net729
rlabel metal1 16146 7276 16146 7276 0 net73
rlabel metal1 8372 12614 8372 12614 0 net730
rlabel metal1 8924 13158 8924 13158 0 net731
rlabel metal2 11638 11798 11638 11798 0 net732
rlabel metal1 12650 12410 12650 12410 0 net733
rlabel metal1 10902 12954 10902 12954 0 net734
rlabel metal1 13570 12240 13570 12240 0 net735
rlabel metal1 13570 13838 13570 13838 0 net736
rlabel metal1 12420 13974 12420 13974 0 net737
rlabel metal1 13248 12954 13248 12954 0 net738
rlabel metal1 18354 13702 18354 13702 0 net739
rlabel metal1 9338 7344 9338 7344 0 net74
rlabel metal2 15134 11832 15134 11832 0 net740
rlabel metal1 16698 10064 16698 10064 0 net741
rlabel metal1 18400 10574 18400 10574 0 net742
rlabel metal1 16008 11866 16008 11866 0 net743
rlabel metal1 15134 12410 15134 12410 0 net744
rlabel metal1 16192 12410 16192 12410 0 net745
rlabel metal1 17894 8466 17894 8466 0 net746
rlabel metal1 14858 9486 14858 9486 0 net747
rlabel metal1 15732 9486 15732 9486 0 net748
rlabel metal1 14490 9146 14490 9146 0 net749
rlabel metal1 16284 4658 16284 4658 0 net75
rlabel metal1 15778 10064 15778 10064 0 net750
rlabel metal1 15732 9146 15732 9146 0 net751
rlabel via2 15870 10013 15870 10013 0 net752
rlabel metal1 13294 10132 13294 10132 0 net753
rlabel metal2 11270 10540 11270 10540 0 net754
rlabel metal1 13754 10064 13754 10064 0 net755
rlabel metal1 10810 10132 10810 10132 0 net756
rlabel metal1 12558 11186 12558 11186 0 net757
rlabel metal2 11730 9248 11730 9248 0 net758
rlabel metal1 12466 11050 12466 11050 0 net759
rlabel metal1 14669 6834 14669 6834 0 net76
rlabel metal1 7958 10540 7958 10540 0 net760
rlabel metal1 9000 9146 9000 9146 0 net761
rlabel metal1 8602 10642 8602 10642 0 net762
rlabel metal1 7498 9044 7498 9044 0 net763
rlabel metal1 10166 8058 10166 8058 0 net764
rlabel metal2 8050 10336 8050 10336 0 net765
rlabel metal1 8372 9418 8372 9418 0 net766
rlabel metal1 6946 8398 6946 8398 0 net767
rlabel metal1 9522 7922 9522 7922 0 net768
rlabel metal1 7866 10778 7866 10778 0 net769
rlabel metal1 16422 6766 16422 6766 0 net77
rlabel metal1 7314 7922 7314 7922 0 net770
rlabel metal1 8234 8602 8234 8602 0 net771
rlabel via1 8786 6749 8786 6749 0 net772
rlabel metal1 8924 8058 8924 8058 0 net773
rlabel metal2 8556 6834 8556 6834 0 net774
rlabel metal1 9476 7310 9476 7310 0 net775
rlabel metal1 16422 7344 16422 7344 0 net79
rlabel metal1 8487 12886 8487 12886 0 net8
rlabel metal2 15318 8160 15318 8160 0 net80
rlabel metal1 20010 7378 20010 7378 0 net81
rlabel metal1 16284 6970 16284 6970 0 net83
rlabel metal1 17797 7922 17797 7922 0 net84
rlabel metal1 20562 5168 20562 5168 0 net85
rlabel metal1 19090 6154 19090 6154 0 net87
rlabel metal1 18119 7242 18119 7242 0 net88
rlabel metal2 23230 6494 23230 6494 0 net89
rlabel metal2 9522 11373 9522 11373 0 net9
rlabel metal1 20746 6834 20746 6834 0 net91
rlabel metal1 16176 6154 16176 6154 0 net92
rlabel metal1 20930 6800 20930 6800 0 net93
rlabel metal1 20240 5270 20240 5270 0 net95
rlabel metal1 18349 5746 18349 5746 0 net96
rlabel metal1 22678 5678 22678 5678 0 net97
rlabel metal1 20838 4624 20838 4624 0 net99
rlabel metal1 20792 3366 20792 3366 0 o_result_ctr[0]
rlabel metal1 20148 4250 20148 4250 0 o_result_ctr[1]
rlabel metal1 20102 4182 20102 4182 0 o_result_ctr[2]
rlabel metal1 16100 5542 16100 5542 0 o_result_ctr[3]
rlabel metal2 9062 1962 9062 1962 0 o_result_ctr[4]
rlabel metal2 10350 1860 10350 1860 0 o_result_ctr[5]
rlabel metal2 11638 2676 11638 2676 0 o_result_ctr[6]
rlabel metal1 11224 5610 11224 5610 0 o_result_ctr[7]
rlabel metal1 13800 6630 13800 6630 0 o_result_ring[0]
rlabel metal3 23230 7208 23230 7208 0 o_result_ring[10]
rlabel metal1 24794 7752 24794 7752 0 o_result_ring[11]
rlabel via2 22862 8517 22862 8517 0 o_result_ring[12]
rlabel metal4 20700 6460 20700 6460 0 o_result_ring[13]
rlabel via2 31702 8228 31702 8228 0 o_result_ring[14]
rlabel metal2 23322 9265 23322 9265 0 o_result_ring[15]
rlabel metal2 28290 9911 28290 9911 0 o_result_ring[16]
rlabel metal2 28290 10829 28290 10829 0 o_result_ring[17]
rlabel metal2 20194 9792 20194 9792 0 o_result_ring[18]
rlabel metal2 23322 11509 23322 11509 0 o_result_ring[19]
rlabel metal1 14536 7718 14536 7718 0 o_result_ring[1]
rlabel metal1 20332 11866 20332 11866 0 o_result_ring[20]
rlabel metal2 24150 11390 24150 11390 0 o_result_ring[21]
rlabel metal1 20148 12954 20148 12954 0 o_result_ring[22]
rlabel metal2 28290 12359 28290 12359 0 o_result_ring[23]
rlabel metal1 24219 13158 24219 13158 0 o_result_ring[24]
rlabel metal1 25806 13158 25806 13158 0 o_result_ring[25]
rlabel metal1 23552 13974 23552 13974 0 o_result_ring[26]
rlabel metal1 24012 14246 24012 14246 0 o_result_ring[27]
rlabel metal2 23230 17350 23230 17350 0 o_result_ring[28]
rlabel metal1 20378 14824 20378 14824 0 o_result_ring[29]
rlabel metal2 15502 1557 15502 1557 0 o_result_ring[2]
rlabel metal1 20470 15130 20470 15130 0 o_result_ring[30]
rlabel metal1 20608 13498 20608 13498 0 o_result_ring[31]
rlabel via2 18630 15045 18630 15045 0 o_result_ring[32]
rlabel metal2 19090 13583 19090 13583 0 o_result_ring[33]
rlabel metal1 17020 15130 17020 15130 0 o_result_ring[34]
rlabel metal1 13892 13974 13892 13974 0 o_result_ring[35]
rlabel metal1 16008 14586 16008 14586 0 o_result_ring[36]
rlabel metal2 13662 15487 13662 15487 0 o_result_ring[37]
rlabel metal1 11960 14790 11960 14790 0 o_result_ring[38]
rlabel metal1 10672 14586 10672 14586 0 o_result_ring[39]
rlabel metal2 16790 1557 16790 1557 0 o_result_ring[3]
rlabel metal1 9982 14042 9982 14042 0 o_result_ring[40]
rlabel metal2 13386 14688 13386 14688 0 o_result_ring[41]
rlabel metal3 1533 12988 1533 12988 0 o_result_ring[42]
rlabel metal1 11408 11866 11408 11866 0 o_result_ring[43]
rlabel metal2 11730 12427 11730 12427 0 o_result_ring[44]
rlabel metal1 15226 12954 15226 12954 0 o_result_ring[45]
rlabel metal2 14306 16014 14306 16014 0 o_result_ring[46]
rlabel metal1 17158 13498 17158 13498 0 o_result_ring[47]
rlabel metal1 18308 12954 18308 12954 0 o_result_ring[48]
rlabel metal1 18492 11866 18492 11866 0 o_result_ring[49]
rlabel metal2 18722 415 18722 415 0 o_result_ring[4]
rlabel metal2 19458 10948 19458 10948 0 o_result_ring[50]
rlabel metal1 18676 10234 18676 10234 0 o_result_ring[51]
rlabel metal1 19780 4590 19780 4590 0 o_result_ring[52]
rlabel metal2 17434 1557 17434 1557 0 o_result_ring[53]
rlabel metal2 14858 1571 14858 1571 0 o_result_ring[54]
rlabel metal1 15594 16150 15594 16150 0 o_result_ring[55]
rlabel metal3 13455 15980 13455 15980 0 o_result_ring[56]
rlabel metal3 1533 10948 1533 10948 0 o_result_ring[57]
rlabel metal3 1533 10268 1533 10268 0 o_result_ring[58]
rlabel via2 8694 9605 8694 9605 0 o_result_ring[59]
rlabel metal2 20010 1557 20010 1557 0 o_result_ring[5]
rlabel metal2 13018 6891 13018 6891 0 o_result_ring[60]
rlabel metal3 1533 8228 1533 8228 0 o_result_ring[61]
rlabel metal2 11776 6324 11776 6324 0 o_result_ring[62]
rlabel metal2 12328 5644 12328 5644 0 o_result_ring[63]
rlabel metal1 17802 6358 17802 6358 0 o_result_ring[6]
rlabel metal2 22586 415 22586 415 0 o_result_ring[7]
rlabel metal1 21114 6154 21114 6154 0 o_result_ring[8]
rlabel metal2 22678 6409 22678 6409 0 o_result_ring[9]
rlabel metal2 17066 3774 17066 3774 0 r_ring_ctr\[0\]
rlabel metal2 15870 4556 15870 4556 0 r_ring_ctr\[1\]
rlabel via1 17337 5134 17337 5134 0 r_ring_ctr\[2\]
rlabel via1 14490 5882 14490 5882 0 r_ring_ctr\[3\]
rlabel metal2 13018 3740 13018 3740 0 r_ring_ctr\[4\]
rlabel metal1 10442 4658 10442 4658 0 r_ring_ctr\[5\]
rlabel metal1 10580 4726 10580 4726 0 r_ring_ctr\[6\]
rlabel metal1 10810 5848 10810 5848 0 r_ring_ctr\[7\]
rlabel metal1 6312 7310 6312 7310 0 w_dly_strt\[10\]
rlabel metal1 8108 6222 8108 6222 0 w_dly_strt\[11\]
rlabel metal1 7797 6426 7797 6426 0 w_dly_strt\[12\]
rlabel metal1 7199 6970 7199 6970 0 w_dly_strt\[13\]
rlabel metal1 7009 6834 7009 6834 0 w_dly_strt\[14\]
rlabel metal1 8389 6222 8389 6222 0 w_dly_strt\[15\]
rlabel metal1 9361 6426 9361 6426 0 w_dly_strt\[16\]
rlabel metal1 8487 5542 8487 5542 0 w_dly_strt\[1\]
rlabel metal1 7958 5746 7958 5746 0 w_dly_strt\[2\]
rlabel metal1 7291 5610 7291 5610 0 w_dly_strt\[3\]
rlabel metal1 7239 5746 7239 5746 0 w_dly_strt\[4\]
rlabel via1 7843 5882 7843 5882 0 w_dly_strt\[5\]
rlabel metal1 7613 6086 7613 6086 0 w_dly_strt\[6\]
rlabel metal1 7664 6222 7664 6222 0 w_dly_strt\[7\]
rlabel metal1 7457 6222 7457 6222 0 w_dly_strt\[8\]
rlabel metal1 7199 6086 7199 6086 0 w_dly_strt\[9\]
rlabel metal1 15318 5746 15318 5746 0 w_ring_ctr_clk
rlabel metal1 8694 6256 8694 6256 0 w_strt_pulse
<< properties >>
string FIXED_BBOX 0 0 32000 20000
<< end >>
