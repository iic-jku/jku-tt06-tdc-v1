magic
tech sky130A
magscale 1 2
timestamp 1710546466
<< viali >>
rect 14289 14569 14323 14603
rect 15853 14569 15887 14603
rect 12909 14433 12943 14467
rect 13176 14433 13210 14467
rect 14473 14433 14507 14467
rect 14740 14433 14774 14467
rect 18337 14433 18371 14467
rect 18429 14229 18463 14263
rect 12909 14025 12943 14059
rect 14841 14025 14875 14059
rect 17601 14025 17635 14059
rect 20085 14025 20119 14059
rect 11529 13889 11563 13923
rect 17877 13889 17911 13923
rect 18429 13889 18463 13923
rect 10977 13821 11011 13855
rect 11437 13821 11471 13855
rect 11785 13821 11819 13855
rect 13921 13821 13955 13855
rect 14565 13821 14599 13855
rect 14749 13821 14783 13855
rect 15117 13821 15151 13855
rect 16221 13821 16255 13855
rect 17785 13821 17819 13855
rect 18061 13821 18095 13855
rect 18153 13821 18187 13855
rect 18521 13821 18555 13855
rect 18705 13821 18739 13855
rect 18961 13821 18995 13855
rect 20545 13821 20579 13855
rect 20637 13821 20671 13855
rect 16466 13753 16500 13787
rect 11069 13685 11103 13719
rect 11345 13685 11379 13719
rect 14013 13685 14047 13719
rect 14473 13685 14507 13719
rect 15209 13685 15243 13719
rect 20453 13685 20487 13719
rect 20729 13685 20763 13719
rect 11529 13481 11563 13515
rect 12541 13481 12575 13515
rect 14013 13481 14047 13515
rect 14473 13481 14507 13515
rect 15577 13481 15611 13515
rect 16221 13481 16255 13515
rect 17325 13481 17359 13515
rect 18981 13481 19015 13515
rect 21005 13481 21039 13515
rect 13093 13413 13127 13447
rect 15301 13413 15335 13447
rect 19441 13413 19475 13447
rect 10793 13345 10827 13379
rect 10977 13345 11011 13379
rect 11621 13345 11655 13379
rect 11713 13345 11747 13379
rect 12173 13345 12207 13379
rect 12265 13345 12299 13379
rect 12633 13345 12667 13379
rect 12817 13345 12851 13379
rect 12909 13345 12943 13379
rect 13001 13345 13035 13379
rect 13369 13345 13403 13379
rect 13829 13345 13863 13379
rect 13921 13345 13955 13379
rect 14381 13345 14415 13379
rect 14657 13345 14691 13379
rect 14933 13345 14967 13379
rect 15209 13345 15243 13379
rect 15485 13345 15519 13379
rect 15761 13345 15795 13379
rect 15853 13345 15887 13379
rect 16129 13345 16163 13379
rect 16589 13345 16623 13379
rect 16681 13345 16715 13379
rect 17141 13345 17175 13379
rect 17417 13345 17451 13379
rect 17601 13345 17635 13379
rect 17857 13345 17891 13379
rect 19533 13345 19567 13379
rect 19625 13345 19659 13379
rect 19881 13345 19915 13379
rect 13737 13277 13771 13311
rect 14749 13277 14783 13311
rect 15025 13277 15059 13311
rect 13461 13209 13495 13243
rect 10701 13141 10735 13175
rect 11069 13141 11103 13175
rect 11805 13141 11839 13175
rect 17049 13141 17083 13175
rect 10057 12937 10091 12971
rect 12909 12937 12943 12971
rect 17969 12937 18003 12971
rect 18797 12937 18831 12971
rect 19349 12937 19383 12971
rect 20453 12937 20487 12971
rect 22017 12937 22051 12971
rect 19625 12869 19659 12903
rect 23581 12869 23615 12903
rect 14749 12801 14783 12835
rect 20637 12801 20671 12835
rect 11170 12733 11204 12767
rect 11437 12733 11471 12767
rect 11713 12733 11747 12767
rect 11989 12733 12023 12767
rect 12265 12733 12299 12767
rect 12725 12733 12759 12767
rect 12817 12733 12851 12767
rect 16589 12733 16623 12767
rect 18153 12733 18187 12767
rect 18705 12733 18739 12767
rect 19165 12733 19199 12767
rect 19441 12733 19475 12767
rect 19533 12733 19567 12767
rect 19809 12733 19843 12767
rect 20085 12733 20119 12767
rect 20361 12733 20395 12767
rect 22201 12733 22235 12767
rect 12081 12665 12115 12699
rect 16497 12665 16531 12699
rect 16856 12665 16890 12699
rect 18245 12665 18279 12699
rect 19073 12665 19107 12699
rect 20882 12665 20916 12699
rect 22446 12665 22480 12699
rect 11621 12597 11655 12631
rect 12357 12597 12391 12631
rect 12633 12597 12667 12631
rect 19901 12597 19935 12631
rect 20177 12597 20211 12631
rect 9045 12393 9079 12427
rect 11345 12393 11379 12427
rect 11621 12393 11655 12427
rect 11989 12393 12023 12427
rect 13553 12393 13587 12427
rect 15117 12393 15151 12427
rect 15669 12393 15703 12427
rect 16313 12393 16347 12427
rect 18429 12393 18463 12427
rect 19257 12393 19291 12427
rect 22845 12393 22879 12427
rect 24777 12393 24811 12427
rect 10158 12257 10192 12291
rect 10793 12257 10827 12291
rect 10977 12257 11011 12291
rect 11437 12257 11471 12291
rect 11713 12257 11747 12291
rect 12081 12257 12115 12291
rect 12173 12257 12207 12291
rect 12429 12257 12463 12291
rect 13737 12257 13771 12291
rect 14004 12257 14038 12291
rect 15577 12257 15611 12291
rect 16221 12257 16255 12291
rect 16957 12257 16991 12291
rect 19165 12257 19199 12291
rect 19809 12257 19843 12291
rect 19901 12257 19935 12291
rect 20177 12257 20211 12291
rect 20637 12257 20671 12291
rect 20729 12257 20763 12291
rect 21557 12257 21591 12291
rect 23397 12257 23431 12291
rect 23653 12257 23687 12291
rect 10425 12189 10459 12223
rect 20821 12189 20855 12223
rect 11069 12121 11103 12155
rect 19993 12121 20027 12155
rect 20545 12121 20579 12155
rect 10701 12053 10735 12087
rect 19717 12053 19751 12087
rect 20269 12053 20303 12087
rect 9413 11849 9447 11883
rect 12725 11849 12759 11883
rect 15393 11849 15427 11883
rect 18429 11849 18463 11883
rect 21925 11849 21959 11883
rect 23581 11849 23615 11883
rect 12449 11781 12483 11815
rect 20821 11781 20855 11815
rect 21649 11781 21683 11815
rect 22201 11713 22235 11747
rect 9045 11645 9079 11679
rect 9481 11639 9515 11673
rect 9605 11639 9639 11673
rect 11805 11645 11839 11679
rect 12265 11645 12299 11679
rect 12541 11645 12575 11679
rect 12633 11645 12667 11679
rect 14013 11645 14047 11679
rect 17049 11645 17083 11679
rect 19809 11645 19843 11679
rect 20085 11645 20119 11679
rect 20361 11645 20395 11679
rect 20637 11645 20671 11679
rect 20729 11645 20763 11679
rect 21189 11645 21223 11679
rect 21465 11645 21499 11679
rect 21557 11645 21591 11679
rect 21833 11645 21867 11679
rect 9137 11577 9171 11611
rect 9873 11577 9907 11611
rect 14258 11577 14292 11611
rect 17316 11577 17350 11611
rect 19993 11577 20027 11611
rect 20545 11577 20579 11611
rect 22446 11577 22480 11611
rect 9689 11509 9723 11543
rect 11161 11509 11195 11543
rect 11897 11509 11931 11543
rect 12173 11509 12207 11543
rect 19717 11509 19751 11543
rect 20269 11509 20303 11543
rect 21097 11509 21131 11543
rect 21373 11509 21407 11543
rect 8125 11305 8159 11339
rect 10333 11305 10367 11339
rect 10609 11305 10643 11339
rect 11069 11305 11103 11339
rect 11345 11305 11379 11339
rect 14197 11305 14231 11339
rect 15761 11305 15795 11339
rect 17509 11305 17543 11339
rect 20913 11305 20947 11339
rect 21925 11305 21959 11339
rect 22477 11305 22511 11339
rect 24317 11305 24351 11339
rect 9238 11237 9272 11271
rect 20729 11237 20763 11271
rect 21649 11237 21683 11271
rect 9689 11169 9723 11203
rect 10057 11169 10091 11203
rect 10149 11169 10183 11203
rect 10425 11169 10459 11203
rect 10701 11169 10735 11203
rect 11161 11169 11195 11203
rect 12458 11169 12492 11203
rect 12725 11169 12759 11203
rect 12817 11169 12851 11203
rect 13073 11169 13107 11203
rect 14381 11169 14415 11203
rect 14648 11169 14682 11203
rect 16129 11169 16163 11203
rect 16385 11169 16419 11203
rect 19073 11169 19107 11203
rect 21005 11169 21039 11203
rect 21281 11169 21315 11203
rect 21557 11169 21591 11203
rect 21833 11169 21867 11203
rect 22293 11169 22327 11203
rect 22569 11169 22603 11203
rect 22661 11169 22695 11203
rect 23193 11169 23227 11203
rect 9505 11101 9539 11135
rect 19349 11101 19383 11135
rect 22937 11101 22971 11135
rect 9781 11033 9815 11067
rect 21373 11033 21407 11067
rect 22201 11033 22235 11067
rect 22753 10965 22787 10999
rect 9781 10761 9815 10795
rect 10057 10761 10091 10795
rect 10333 10761 10367 10795
rect 11897 10761 11931 10795
rect 18429 10761 18463 10795
rect 15945 10693 15979 10727
rect 22017 10693 22051 10727
rect 10517 10625 10551 10659
rect 10793 10625 10827 10659
rect 22293 10625 22327 10659
rect 9137 10557 9171 10591
rect 9597 10557 9631 10591
rect 9689 10557 9723 10591
rect 10149 10557 10183 10591
rect 10241 10557 10275 10591
rect 14473 10557 14507 10591
rect 15209 10557 15243 10591
rect 15761 10557 15795 10591
rect 15853 10557 15887 10591
rect 17049 10557 17083 10591
rect 21649 10557 21683 10591
rect 22109 10557 22143 10591
rect 22385 10557 22419 10591
rect 22661 10557 22695 10591
rect 22753 10557 22787 10591
rect 9229 10489 9263 10523
rect 9505 10489 9539 10523
rect 17294 10489 17328 10523
rect 21741 10489 21775 10523
rect 22569 10489 22603 10523
rect 14381 10421 14415 10455
rect 15301 10421 15335 10455
rect 15669 10421 15703 10455
rect 22845 10421 22879 10455
rect 7113 10217 7147 10251
rect 9873 10217 9907 10251
rect 10149 10217 10183 10251
rect 15301 10217 15335 10251
rect 22753 10217 22787 10251
rect 24317 10217 24351 10251
rect 8769 10149 8803 10183
rect 9597 10149 9631 10183
rect 23182 10149 23216 10183
rect 8237 10081 8271 10115
rect 8493 10081 8527 10115
rect 8861 10081 8895 10115
rect 9137 10081 9171 10115
rect 9689 10081 9723 10115
rect 9781 10081 9815 10115
rect 10241 10081 10275 10115
rect 14565 10081 14599 10115
rect 14657 10081 14691 10115
rect 15117 10081 15151 10115
rect 15393 10081 15427 10115
rect 15669 10081 15703 10115
rect 15945 10081 15979 10115
rect 16129 10081 16163 10115
rect 18153 10081 18187 10115
rect 18593 10081 18627 10115
rect 21465 10081 21499 10115
rect 21741 10081 21775 10115
rect 22025 10081 22059 10115
rect 22293 10087 22327 10121
rect 22385 10081 22419 10115
rect 22845 10081 22879 10115
rect 22937 10081 22971 10115
rect 9045 10013 9079 10047
rect 13921 10013 13955 10047
rect 14197 10013 14231 10047
rect 18337 10013 18371 10047
rect 21373 10013 21407 10047
rect 15577 9945 15611 9979
rect 21649 9945 21683 9979
rect 22477 9945 22511 9979
rect 12633 9877 12667 9911
rect 14473 9877 14507 9911
rect 14749 9877 14783 9911
rect 15025 9877 15059 9911
rect 15853 9877 15887 9911
rect 17601 9877 17635 9911
rect 18061 9877 18095 9911
rect 19717 9877 19751 9911
rect 21925 9877 21959 9911
rect 22201 9877 22235 9911
rect 8493 9673 8527 9707
rect 8861 9673 8895 9707
rect 9137 9673 9171 9707
rect 14565 9673 14599 9707
rect 16129 9673 16163 9707
rect 16405 9673 16439 9707
rect 16681 9673 16715 9707
rect 17693 9673 17727 9707
rect 9781 9605 9815 9639
rect 17233 9605 17267 9639
rect 13001 9537 13035 9571
rect 8217 9469 8251 9503
rect 8585 9469 8619 9503
rect 8953 9469 8987 9503
rect 9229 9469 9263 9503
rect 9321 9469 9355 9503
rect 10894 9469 10928 9503
rect 11161 9469 11195 9503
rect 13277 9469 13311 9503
rect 13553 9469 13587 9503
rect 14381 9469 14415 9503
rect 14657 9469 14691 9503
rect 14933 9469 14967 9503
rect 15025 9469 15059 9503
rect 16221 9469 16255 9503
rect 16497 9469 16531 9503
rect 16773 9469 16807 9503
rect 17049 9469 17083 9503
rect 17325 9469 17359 9503
rect 17785 9469 17819 9503
rect 18061 9469 18095 9503
rect 18337 9469 18371 9503
rect 18889 9469 18923 9503
rect 18981 9469 19015 9503
rect 19349 9469 19383 9503
rect 22017 9469 22051 9503
rect 8125 9401 8159 9435
rect 12756 9401 12790 9435
rect 13185 9401 13219 9435
rect 15117 9401 15151 9435
rect 17969 9401 18003 9435
rect 18245 9401 18279 9435
rect 18797 9401 18831 9435
rect 19594 9401 19628 9435
rect 22284 9401 22318 9435
rect 9413 9333 9447 9367
rect 11621 9333 11655 9367
rect 13645 9333 13679 9367
rect 14289 9333 14323 9367
rect 14841 9333 14875 9367
rect 16957 9333 16991 9367
rect 19073 9333 19107 9367
rect 20729 9333 20763 9367
rect 23397 9333 23431 9367
rect 8309 9129 8343 9163
rect 8861 9129 8895 9163
rect 9137 9129 9171 9163
rect 13001 9129 13035 9163
rect 17969 9129 18003 9163
rect 18797 9129 18831 9163
rect 19073 9129 19107 9163
rect 19349 9129 19383 9163
rect 19901 9129 19935 9163
rect 7880 9061 7914 9095
rect 10526 9061 10560 9095
rect 16488 9061 16522 9095
rect 18245 9061 18279 9095
rect 18521 9061 18555 9095
rect 8125 8993 8159 9027
rect 8401 8993 8435 9027
rect 8493 8993 8527 9027
rect 8953 8993 8987 9027
rect 9045 8993 9079 9027
rect 12817 8993 12851 9027
rect 13101 8993 13135 9027
rect 13553 8993 13587 9027
rect 13829 8993 13863 9027
rect 14105 8993 14139 9027
rect 14381 8993 14415 9027
rect 14729 8993 14763 9027
rect 18061 8993 18095 9027
rect 18337 8993 18371 9027
rect 18613 8993 18647 9027
rect 18889 8993 18923 9027
rect 19165 8993 19199 9027
rect 19441 8993 19475 9027
rect 19625 8993 19659 9027
rect 19717 8993 19751 9027
rect 19993 8993 20027 9027
rect 20085 8993 20119 9027
rect 20545 8993 20579 9027
rect 20729 8993 20763 9027
rect 20821 8993 20855 9027
rect 10793 8925 10827 8959
rect 14473 8925 14507 8959
rect 16221 8925 16255 8959
rect 21465 8925 21499 8959
rect 21741 8925 21775 8959
rect 6745 8857 6779 8891
rect 12725 8857 12759 8891
rect 13461 8857 13495 8891
rect 20453 8857 20487 8891
rect 8585 8789 8619 8823
rect 9413 8789 9447 8823
rect 13737 8789 13771 8823
rect 14013 8789 14047 8823
rect 14289 8789 14323 8823
rect 15853 8789 15887 8823
rect 17601 8789 17635 8823
rect 20177 8789 20211 8823
rect 23029 8789 23063 8823
rect 8677 8585 8711 8619
rect 8953 8585 8987 8619
rect 22661 8585 22695 8619
rect 13645 8517 13679 8551
rect 21189 8517 21223 8551
rect 8125 8449 8159 8483
rect 12817 8449 12851 8483
rect 19798 8449 19832 8483
rect 7941 8381 7975 8415
rect 8217 8381 8251 8415
rect 8769 8381 8803 8415
rect 9045 8381 9079 8415
rect 10701 8381 10735 8415
rect 12561 8381 12595 8415
rect 13185 8381 13219 8415
rect 13553 8381 13587 8415
rect 14013 8381 14047 8415
rect 14289 8381 14323 8415
rect 14381 8381 14415 8415
rect 14657 8381 14691 8415
rect 19441 8381 19475 8415
rect 19717 8381 19751 8415
rect 21373 8381 21407 8415
rect 23213 8381 23247 8415
rect 7849 8313 7883 8347
rect 10434 8313 10468 8347
rect 13921 8313 13955 8347
rect 14197 8313 14231 8347
rect 14902 8313 14936 8347
rect 20076 8313 20110 8347
rect 9321 8245 9355 8279
rect 11437 8245 11471 8279
rect 13277 8245 13311 8279
rect 14473 8245 14507 8279
rect 16037 8245 16071 8279
rect 19349 8245 19383 8279
rect 19625 8245 19659 8279
rect 23305 8245 23339 8279
rect 8309 8041 8343 8075
rect 13461 8041 13495 8075
rect 19901 8041 19935 8075
rect 10793 7973 10827 8007
rect 15945 7973 15979 8007
rect 18052 7973 18086 8007
rect 20453 7973 20487 8007
rect 21373 7973 21407 8007
rect 21649 7973 21683 8007
rect 7766 7905 7800 7939
rect 8401 7905 8435 7939
rect 8677 7905 8711 7939
rect 8953 7905 8987 7939
rect 12182 7905 12216 7939
rect 13001 7905 13035 7939
rect 13093 7905 13127 7939
rect 13553 7905 13587 7939
rect 13829 7905 13863 7939
rect 14105 7905 14139 7939
rect 16129 7905 16163 7939
rect 16385 7905 16419 7939
rect 19993 7905 20027 7939
rect 20269 7903 20303 7937
rect 20361 7905 20395 7939
rect 20821 7905 20855 7939
rect 21005 7905 21039 7939
rect 21097 7905 21131 7939
rect 21281 7905 21315 7939
rect 21741 7905 21775 7939
rect 21925 7905 21959 7939
rect 22181 7905 22215 7939
rect 8033 7837 8067 7871
rect 8861 7837 8895 7871
rect 12449 7837 12483 7871
rect 17785 7837 17819 7871
rect 8585 7769 8619 7803
rect 13185 7769 13219 7803
rect 13737 7769 13771 7803
rect 20177 7769 20211 7803
rect 6653 7701 6687 7735
rect 9505 7701 9539 7735
rect 11069 7701 11103 7735
rect 12909 7701 12943 7735
rect 14013 7701 14047 7735
rect 14657 7701 14691 7735
rect 17509 7701 17543 7735
rect 19165 7701 19199 7735
rect 20729 7701 20763 7735
rect 23305 7701 23339 7735
rect 7849 7497 7883 7531
rect 9137 7497 9171 7531
rect 10333 7497 10367 7531
rect 12725 7497 12759 7531
rect 14381 7497 14415 7531
rect 20269 7497 20303 7531
rect 21649 7497 21683 7531
rect 7573 7429 7607 7463
rect 8861 7429 8895 7463
rect 11897 7429 11931 7463
rect 19993 7429 20027 7463
rect 9505 7361 9539 7395
rect 10057 7361 10091 7395
rect 13829 7361 13863 7395
rect 22017 7361 22051 7395
rect 7665 7293 7699 7327
rect 7941 7293 7975 7327
rect 8033 7293 8067 7327
rect 8125 7293 8159 7327
rect 8585 7293 8619 7327
rect 8945 7295 8979 7329
rect 9045 7293 9079 7327
rect 9597 7293 9631 7327
rect 9873 7293 9907 7327
rect 9965 7293 9999 7327
rect 10425 7293 10459 7327
rect 11989 7293 12023 7327
rect 12173 7293 12207 7327
rect 12265 7293 12299 7327
rect 12541 7293 12575 7327
rect 12633 7303 12667 7337
rect 13093 7293 13127 7327
rect 13185 7293 13219 7327
rect 13921 7293 13955 7327
rect 14013 7293 14047 7327
rect 14289 7293 14323 7327
rect 15770 7293 15804 7327
rect 16037 7293 16071 7327
rect 18521 7293 18555 7327
rect 19349 7293 19383 7327
rect 19809 7293 19843 7327
rect 19901 7293 19935 7327
rect 20361 7293 20395 7327
rect 20453 7293 20487 7327
rect 20737 7293 20771 7327
rect 21189 7293 21223 7327
rect 21281 7293 21315 7327
rect 21373 7293 21407 7327
rect 21741 7293 21775 7327
rect 8493 7225 8527 7259
rect 9781 7225 9815 7259
rect 13001 7225 13035 7259
rect 19441 7225 19475 7259
rect 19717 7225 19751 7259
rect 20545 7225 20579 7259
rect 20821 7225 20855 7259
rect 22284 7225 22318 7259
rect 12449 7157 12483 7191
rect 13277 7157 13311 7191
rect 14105 7157 14139 7191
rect 14657 7157 14691 7191
rect 17049 7157 17083 7191
rect 21097 7157 21131 7191
rect 23397 7157 23431 7191
rect 9413 6953 9447 6987
rect 10425 6953 10459 6987
rect 19809 6953 19843 6987
rect 20361 6953 20395 6987
rect 20637 6953 20671 6987
rect 20913 6953 20947 6987
rect 10149 6885 10183 6919
rect 13912 6885 13946 6919
rect 19257 6885 19291 6919
rect 19533 6885 19567 6919
rect 8962 6817 8996 6851
rect 9505 6817 9539 6851
rect 9781 6817 9815 6851
rect 9873 6817 9907 6851
rect 10057 6817 10091 6851
rect 10517 6817 10551 6851
rect 10793 6817 10827 6851
rect 11161 6817 11195 6851
rect 11437 6817 11471 6851
rect 11713 6817 11747 6851
rect 11989 6807 12023 6841
rect 12265 6817 12299 6851
rect 12357 6817 12391 6851
rect 17049 6817 17083 6851
rect 17316 6817 17350 6851
rect 18613 6817 18647 6851
rect 18889 6817 18923 6851
rect 19341 6817 19375 6851
rect 19441 6823 19475 6857
rect 19717 6817 19751 6851
rect 19993 6817 20027 6851
rect 20453 6817 20487 6851
rect 20545 6817 20579 6851
rect 20821 6817 20855 6851
rect 21281 6817 21315 6851
rect 21537 6817 21571 6851
rect 9229 6749 9263 6783
rect 13645 6749 13679 6783
rect 18705 6749 18739 6783
rect 11897 6681 11931 6715
rect 12173 6681 12207 6715
rect 20085 6681 20119 6715
rect 7849 6613 7883 6647
rect 10701 6613 10735 6647
rect 11069 6613 11103 6647
rect 11345 6613 11379 6647
rect 11621 6613 11655 6647
rect 12449 6613 12483 6647
rect 15025 6613 15059 6647
rect 18429 6613 18463 6647
rect 18981 6613 19015 6647
rect 22661 6613 22695 6647
rect 10609 6409 10643 6443
rect 10977 6409 11011 6443
rect 17509 6341 17543 6375
rect 18797 6273 18831 6307
rect 10425 6205 10459 6239
rect 10701 6205 10735 6239
rect 11069 6205 11103 6239
rect 11897 6205 11931 6239
rect 14565 6205 14599 6239
rect 16129 6205 16163 6239
rect 16396 6205 16430 6239
rect 17693 6205 17727 6239
rect 17969 6205 18003 6239
rect 18061 6205 18095 6239
rect 18245 6205 18279 6239
rect 19064 6205 19098 6239
rect 20361 6205 20395 6239
rect 10180 6137 10214 6171
rect 12164 6137 12198 6171
rect 14832 6137 14866 6171
rect 17785 6137 17819 6171
rect 20628 6137 20662 6171
rect 9045 6069 9079 6103
rect 13277 6069 13311 6103
rect 15945 6069 15979 6103
rect 18337 6069 18371 6103
rect 20177 6069 20211 6103
rect 21741 6069 21775 6103
rect 16221 5865 16255 5899
rect 17141 5865 17175 5899
rect 17785 5865 17819 5899
rect 19165 5865 19199 5899
rect 11336 5797 11370 5831
rect 18889 5797 18923 5831
rect 11069 5729 11103 5763
rect 15045 5729 15079 5763
rect 15301 5729 15335 5763
rect 16313 5729 16347 5763
rect 16405 5729 16439 5763
rect 16957 5729 16991 5763
rect 17233 5729 17267 5763
rect 17509 5729 17543 5763
rect 17869 5735 17903 5769
rect 17969 5727 18003 5761
rect 18245 5729 18279 5763
rect 18521 5729 18555 5763
rect 18797 5729 18831 5763
rect 19257 5729 19291 5763
rect 16497 5593 16531 5627
rect 16865 5593 16899 5627
rect 18061 5593 18095 5627
rect 18337 5593 18371 5627
rect 12449 5525 12483 5559
rect 13921 5525 13955 5559
rect 17417 5525 17451 5559
rect 18613 5525 18647 5559
rect 15853 5321 15887 5355
rect 16497 5321 16531 5355
rect 17049 5185 17083 5219
rect 15669 5117 15703 5151
rect 15761 5117 15795 5151
rect 16313 5117 16347 5151
rect 16589 5117 16623 5151
rect 16681 5117 16715 5151
rect 16773 5117 16807 5151
rect 17316 5117 17350 5151
rect 15577 5049 15611 5083
rect 18429 4981 18463 5015
rect 16405 4777 16439 4811
rect 16497 4641 16531 4675
rect 22937 833 22971 867
rect 22661 765 22695 799
<< metal1 >>
rect 552 19066 31531 19088
rect 552 19014 8102 19066
rect 8154 19014 8166 19066
rect 8218 19014 8230 19066
rect 8282 19014 8294 19066
rect 8346 19014 8358 19066
rect 8410 19014 15807 19066
rect 15859 19014 15871 19066
rect 15923 19014 15935 19066
rect 15987 19014 15999 19066
rect 16051 19014 16063 19066
rect 16115 19014 23512 19066
rect 23564 19014 23576 19066
rect 23628 19014 23640 19066
rect 23692 19014 23704 19066
rect 23756 19014 23768 19066
rect 23820 19014 31217 19066
rect 31269 19014 31281 19066
rect 31333 19014 31345 19066
rect 31397 19014 31409 19066
rect 31461 19014 31473 19066
rect 31525 19014 31531 19066
rect 552 18992 31531 19014
rect 552 18522 31372 18544
rect 552 18470 4250 18522
rect 4302 18470 4314 18522
rect 4366 18470 4378 18522
rect 4430 18470 4442 18522
rect 4494 18470 4506 18522
rect 4558 18470 11955 18522
rect 12007 18470 12019 18522
rect 12071 18470 12083 18522
rect 12135 18470 12147 18522
rect 12199 18470 12211 18522
rect 12263 18470 19660 18522
rect 19712 18470 19724 18522
rect 19776 18470 19788 18522
rect 19840 18470 19852 18522
rect 19904 18470 19916 18522
rect 19968 18470 27365 18522
rect 27417 18470 27429 18522
rect 27481 18470 27493 18522
rect 27545 18470 27557 18522
rect 27609 18470 27621 18522
rect 27673 18470 31372 18522
rect 552 18448 31372 18470
rect 552 17978 31531 18000
rect 552 17926 8102 17978
rect 8154 17926 8166 17978
rect 8218 17926 8230 17978
rect 8282 17926 8294 17978
rect 8346 17926 8358 17978
rect 8410 17926 15807 17978
rect 15859 17926 15871 17978
rect 15923 17926 15935 17978
rect 15987 17926 15999 17978
rect 16051 17926 16063 17978
rect 16115 17926 23512 17978
rect 23564 17926 23576 17978
rect 23628 17926 23640 17978
rect 23692 17926 23704 17978
rect 23756 17926 23768 17978
rect 23820 17926 31217 17978
rect 31269 17926 31281 17978
rect 31333 17926 31345 17978
rect 31397 17926 31409 17978
rect 31461 17926 31473 17978
rect 31525 17926 31531 17978
rect 552 17904 31531 17926
rect 552 17434 31372 17456
rect 552 17382 4250 17434
rect 4302 17382 4314 17434
rect 4366 17382 4378 17434
rect 4430 17382 4442 17434
rect 4494 17382 4506 17434
rect 4558 17382 11955 17434
rect 12007 17382 12019 17434
rect 12071 17382 12083 17434
rect 12135 17382 12147 17434
rect 12199 17382 12211 17434
rect 12263 17382 19660 17434
rect 19712 17382 19724 17434
rect 19776 17382 19788 17434
rect 19840 17382 19852 17434
rect 19904 17382 19916 17434
rect 19968 17382 27365 17434
rect 27417 17382 27429 17434
rect 27481 17382 27493 17434
rect 27545 17382 27557 17434
rect 27609 17382 27621 17434
rect 27673 17382 31372 17434
rect 552 17360 31372 17382
rect 552 16890 31531 16912
rect 552 16838 8102 16890
rect 8154 16838 8166 16890
rect 8218 16838 8230 16890
rect 8282 16838 8294 16890
rect 8346 16838 8358 16890
rect 8410 16838 15807 16890
rect 15859 16838 15871 16890
rect 15923 16838 15935 16890
rect 15987 16838 15999 16890
rect 16051 16838 16063 16890
rect 16115 16838 23512 16890
rect 23564 16838 23576 16890
rect 23628 16838 23640 16890
rect 23692 16838 23704 16890
rect 23756 16838 23768 16890
rect 23820 16838 31217 16890
rect 31269 16838 31281 16890
rect 31333 16838 31345 16890
rect 31397 16838 31409 16890
rect 31461 16838 31473 16890
rect 31525 16838 31531 16890
rect 552 16816 31531 16838
rect 552 16346 31372 16368
rect 552 16294 4250 16346
rect 4302 16294 4314 16346
rect 4366 16294 4378 16346
rect 4430 16294 4442 16346
rect 4494 16294 4506 16346
rect 4558 16294 11955 16346
rect 12007 16294 12019 16346
rect 12071 16294 12083 16346
rect 12135 16294 12147 16346
rect 12199 16294 12211 16346
rect 12263 16294 19660 16346
rect 19712 16294 19724 16346
rect 19776 16294 19788 16346
rect 19840 16294 19852 16346
rect 19904 16294 19916 16346
rect 19968 16294 27365 16346
rect 27417 16294 27429 16346
rect 27481 16294 27493 16346
rect 27545 16294 27557 16346
rect 27609 16294 27621 16346
rect 27673 16294 31372 16346
rect 552 16272 31372 16294
rect 552 15802 31531 15824
rect 552 15750 8102 15802
rect 8154 15750 8166 15802
rect 8218 15750 8230 15802
rect 8282 15750 8294 15802
rect 8346 15750 8358 15802
rect 8410 15750 15807 15802
rect 15859 15750 15871 15802
rect 15923 15750 15935 15802
rect 15987 15750 15999 15802
rect 16051 15750 16063 15802
rect 16115 15750 23512 15802
rect 23564 15750 23576 15802
rect 23628 15750 23640 15802
rect 23692 15750 23704 15802
rect 23756 15750 23768 15802
rect 23820 15750 31217 15802
rect 31269 15750 31281 15802
rect 31333 15750 31345 15802
rect 31397 15750 31409 15802
rect 31461 15750 31473 15802
rect 31525 15750 31531 15802
rect 552 15728 31531 15750
rect 552 15258 31372 15280
rect 552 15206 4250 15258
rect 4302 15206 4314 15258
rect 4366 15206 4378 15258
rect 4430 15206 4442 15258
rect 4494 15206 4506 15258
rect 4558 15206 11955 15258
rect 12007 15206 12019 15258
rect 12071 15206 12083 15258
rect 12135 15206 12147 15258
rect 12199 15206 12211 15258
rect 12263 15206 19660 15258
rect 19712 15206 19724 15258
rect 19776 15206 19788 15258
rect 19840 15206 19852 15258
rect 19904 15206 19916 15258
rect 19968 15206 27365 15258
rect 27417 15206 27429 15258
rect 27481 15206 27493 15258
rect 27545 15206 27557 15258
rect 27609 15206 27621 15258
rect 27673 15206 31372 15258
rect 552 15184 31372 15206
rect 552 14714 31531 14736
rect 552 14662 8102 14714
rect 8154 14662 8166 14714
rect 8218 14662 8230 14714
rect 8282 14662 8294 14714
rect 8346 14662 8358 14714
rect 8410 14662 15807 14714
rect 15859 14662 15871 14714
rect 15923 14662 15935 14714
rect 15987 14662 15999 14714
rect 16051 14662 16063 14714
rect 16115 14662 23512 14714
rect 23564 14662 23576 14714
rect 23628 14662 23640 14714
rect 23692 14662 23704 14714
rect 23756 14662 23768 14714
rect 23820 14662 31217 14714
rect 31269 14662 31281 14714
rect 31333 14662 31345 14714
rect 31397 14662 31409 14714
rect 31461 14662 31473 14714
rect 31525 14662 31531 14714
rect 552 14640 31531 14662
rect 14182 14560 14188 14612
rect 14240 14600 14246 14612
rect 14277 14603 14335 14609
rect 14277 14600 14289 14603
rect 14240 14572 14289 14600
rect 14240 14560 14246 14572
rect 14277 14569 14289 14572
rect 14323 14569 14335 14603
rect 14277 14563 14335 14569
rect 15841 14603 15899 14609
rect 15841 14569 15853 14603
rect 15887 14600 15899 14603
rect 16758 14600 16764 14612
rect 15887 14572 16764 14600
rect 15887 14569 15899 14572
rect 15841 14563 15899 14569
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 12912 14504 14504 14532
rect 12912 14473 12940 14504
rect 14476 14476 14504 14504
rect 13170 14473 13176 14476
rect 12897 14467 12955 14473
rect 12897 14433 12909 14467
rect 12943 14433 12955 14467
rect 12897 14427 12955 14433
rect 13164 14427 13176 14473
rect 13170 14424 13176 14427
rect 13228 14424 13234 14476
rect 14458 14424 14464 14476
rect 14516 14424 14522 14476
rect 14734 14473 14740 14476
rect 14728 14427 14740 14473
rect 14734 14424 14740 14427
rect 14792 14424 14798 14476
rect 18325 14467 18383 14473
rect 18325 14433 18337 14467
rect 18371 14464 18383 14467
rect 18598 14464 18604 14476
rect 18371 14436 18604 14464
rect 18371 14433 18383 14436
rect 18325 14427 18383 14433
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 18417 14263 18475 14269
rect 18417 14229 18429 14263
rect 18463 14260 18475 14263
rect 19426 14260 19432 14272
rect 18463 14232 19432 14260
rect 18463 14229 18475 14232
rect 18417 14223 18475 14229
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 552 14170 31372 14192
rect 552 14118 4250 14170
rect 4302 14118 4314 14170
rect 4366 14118 4378 14170
rect 4430 14118 4442 14170
rect 4494 14118 4506 14170
rect 4558 14118 11955 14170
rect 12007 14118 12019 14170
rect 12071 14118 12083 14170
rect 12135 14118 12147 14170
rect 12199 14118 12211 14170
rect 12263 14118 19660 14170
rect 19712 14118 19724 14170
rect 19776 14118 19788 14170
rect 19840 14118 19852 14170
rect 19904 14118 19916 14170
rect 19968 14118 27365 14170
rect 27417 14118 27429 14170
rect 27481 14118 27493 14170
rect 27545 14118 27557 14170
rect 27609 14118 27621 14170
rect 27673 14118 31372 14170
rect 552 14096 31372 14118
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12492 14028 12909 14056
rect 12492 14016 12498 14028
rect 12897 14025 12909 14028
rect 12943 14025 12955 14059
rect 12897 14019 12955 14025
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 14829 14059 14887 14065
rect 14829 14056 14841 14059
rect 14792 14028 14841 14056
rect 14792 14016 14798 14028
rect 14829 14025 14841 14028
rect 14875 14025 14887 14059
rect 14829 14019 14887 14025
rect 17589 14059 17647 14065
rect 17589 14025 17601 14059
rect 17635 14056 17647 14059
rect 18046 14056 18052 14068
rect 17635 14028 18052 14056
rect 17635 14025 17647 14028
rect 17589 14019 17647 14025
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14056 20131 14059
rect 20622 14056 20628 14068
rect 20119 14028 20628 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 20622 14016 20628 14028
rect 20680 14016 20686 14068
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 11348 13892 11529 13920
rect 11348 13864 11376 13892
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 13170 13880 13176 13932
rect 13228 13920 13234 13932
rect 17865 13923 17923 13929
rect 13228 13892 14596 13920
rect 13228 13880 13234 13892
rect 10965 13855 11023 13861
rect 10965 13852 10977 13855
rect 10704 13824 10977 13852
rect 10704 13728 10732 13824
rect 10965 13821 10977 13824
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 11330 13812 11336 13864
rect 11388 13812 11394 13864
rect 11422 13812 11428 13864
rect 11480 13812 11486 13864
rect 11773 13855 11831 13861
rect 11773 13852 11785 13855
rect 11532 13824 11785 13852
rect 11532 13784 11560 13824
rect 11773 13821 11785 13824
rect 11819 13852 11831 13855
rect 13446 13852 13452 13864
rect 11819 13824 13452 13852
rect 11819 13821 11831 13824
rect 11773 13815 11831 13821
rect 13446 13812 13452 13824
rect 13504 13852 13510 13864
rect 14568 13861 14596 13892
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 18417 13923 18475 13929
rect 18417 13920 18429 13923
rect 17911 13892 18429 13920
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 18417 13889 18429 13892
rect 18463 13920 18475 13923
rect 18463 13892 18828 13920
rect 18463 13889 18475 13892
rect 18417 13883 18475 13889
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13504 13824 13921 13852
rect 13504 13812 13510 13824
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 13909 13815 13967 13821
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 14737 13855 14795 13861
rect 14737 13821 14749 13855
rect 14783 13852 14795 13855
rect 15105 13855 15163 13861
rect 15105 13852 15117 13855
rect 14783 13824 15117 13852
rect 14783 13821 14795 13824
rect 14737 13815 14795 13821
rect 15105 13821 15117 13824
rect 15151 13821 15163 13855
rect 15105 13815 15163 13821
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13852 16267 13855
rect 16255 13824 17632 13852
rect 16255 13821 16267 13824
rect 16209 13815 16267 13821
rect 14752 13784 14780 13815
rect 16482 13793 16488 13796
rect 16454 13787 16488 13793
rect 16454 13784 16466 13787
rect 11348 13756 11560 13784
rect 14476 13756 14780 13784
rect 15672 13756 16466 13784
rect 10686 13676 10692 13728
rect 10744 13676 10750 13728
rect 11057 13719 11115 13725
rect 11057 13685 11069 13719
rect 11103 13716 11115 13719
rect 11146 13716 11152 13728
rect 11103 13688 11152 13716
rect 11103 13685 11115 13688
rect 11057 13679 11115 13685
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11348 13725 11376 13756
rect 11333 13719 11391 13725
rect 11333 13685 11345 13719
rect 11379 13685 11391 13719
rect 11333 13679 11391 13685
rect 13998 13676 14004 13728
rect 14056 13676 14062 13728
rect 14366 13676 14372 13728
rect 14424 13716 14430 13728
rect 14476 13725 14504 13756
rect 15672 13728 15700 13756
rect 16454 13753 16466 13756
rect 16454 13747 16488 13753
rect 16482 13744 16488 13747
rect 16540 13744 16546 13796
rect 17604 13784 17632 13824
rect 17770 13812 17776 13864
rect 17828 13812 17834 13864
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 18012 13824 18061 13852
rect 18012 13812 18018 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18141 13855 18199 13861
rect 18141 13821 18153 13855
rect 18187 13852 18199 13855
rect 18509 13855 18567 13861
rect 18509 13852 18521 13855
rect 18187 13824 18521 13852
rect 18187 13821 18199 13824
rect 18141 13815 18199 13821
rect 18509 13821 18521 13824
rect 18555 13852 18567 13855
rect 18598 13852 18604 13864
rect 18555 13824 18604 13852
rect 18555 13821 18567 13824
rect 18509 13815 18567 13821
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 18690 13812 18696 13864
rect 18748 13812 18754 13864
rect 18800 13852 18828 13892
rect 20456 13892 20668 13920
rect 18966 13861 18972 13864
rect 18949 13855 18972 13861
rect 18949 13852 18961 13855
rect 18800 13824 18961 13852
rect 18949 13821 18961 13824
rect 18949 13815 18972 13821
rect 18966 13812 18972 13815
rect 19024 13812 19030 13864
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 20456 13852 20484 13892
rect 20640 13861 20668 13892
rect 19484 13824 20484 13852
rect 20533 13855 20591 13861
rect 19484 13812 19490 13824
rect 20533 13821 20545 13855
rect 20579 13821 20591 13855
rect 20533 13815 20591 13821
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 18708 13784 18736 13812
rect 17604 13756 18736 13784
rect 20548 13784 20576 13815
rect 20548 13756 20668 13784
rect 20640 13728 20668 13756
rect 14461 13719 14519 13725
rect 14461 13716 14473 13719
rect 14424 13688 14473 13716
rect 14424 13676 14430 13688
rect 14461 13685 14473 13688
rect 14507 13685 14519 13719
rect 14461 13679 14519 13685
rect 15197 13719 15255 13725
rect 15197 13685 15209 13719
rect 15243 13716 15255 13719
rect 15654 13716 15660 13728
rect 15243 13688 15660 13716
rect 15243 13685 15255 13688
rect 15197 13679 15255 13685
rect 15654 13676 15660 13688
rect 15712 13676 15718 13728
rect 20438 13676 20444 13728
rect 20496 13676 20502 13728
rect 20622 13676 20628 13728
rect 20680 13716 20686 13728
rect 20717 13719 20775 13725
rect 20717 13716 20729 13719
rect 20680 13688 20729 13716
rect 20680 13676 20686 13688
rect 20717 13685 20729 13688
rect 20763 13685 20775 13719
rect 20717 13679 20775 13685
rect 552 13626 31531 13648
rect 552 13574 8102 13626
rect 8154 13574 8166 13626
rect 8218 13574 8230 13626
rect 8282 13574 8294 13626
rect 8346 13574 8358 13626
rect 8410 13574 15807 13626
rect 15859 13574 15871 13626
rect 15923 13574 15935 13626
rect 15987 13574 15999 13626
rect 16051 13574 16063 13626
rect 16115 13574 23512 13626
rect 23564 13574 23576 13626
rect 23628 13574 23640 13626
rect 23692 13574 23704 13626
rect 23756 13574 23768 13626
rect 23820 13574 31217 13626
rect 31269 13574 31281 13626
rect 31333 13574 31345 13626
rect 31397 13574 31409 13626
rect 31461 13574 31473 13626
rect 31525 13574 31531 13626
rect 552 13552 31531 13574
rect 11422 13472 11428 13524
rect 11480 13512 11486 13524
rect 11517 13515 11575 13521
rect 11517 13512 11529 13515
rect 11480 13484 11529 13512
rect 11480 13472 11486 13484
rect 11517 13481 11529 13484
rect 11563 13481 11575 13515
rect 11517 13475 11575 13481
rect 12529 13515 12587 13521
rect 12529 13481 12541 13515
rect 12575 13512 12587 13515
rect 13446 13512 13452 13524
rect 12575 13484 13452 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 13998 13472 14004 13524
rect 14056 13472 14062 13524
rect 14461 13515 14519 13521
rect 14461 13481 14473 13515
rect 14507 13512 14519 13515
rect 14734 13512 14740 13524
rect 14507 13484 14740 13512
rect 14507 13481 14519 13484
rect 14461 13475 14519 13481
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 15565 13515 15623 13521
rect 15565 13481 15577 13515
rect 15611 13512 15623 13515
rect 16209 13515 16267 13521
rect 16209 13512 16221 13515
rect 15611 13484 16221 13512
rect 15611 13481 15623 13484
rect 15565 13475 15623 13481
rect 16209 13481 16221 13484
rect 16255 13481 16267 13515
rect 16209 13475 16267 13481
rect 11146 13404 11152 13456
rect 11204 13444 11210 13456
rect 13081 13447 13139 13453
rect 11204 13416 12204 13444
rect 11204 13404 11210 13416
rect 12176 13385 12204 13416
rect 12820 13416 13032 13444
rect 12820 13385 12848 13416
rect 13004 13385 13032 13416
rect 13081 13413 13093 13447
rect 13127 13444 13139 13447
rect 13170 13444 13176 13456
rect 13127 13416 13176 13444
rect 13127 13413 13139 13416
rect 13081 13407 13139 13413
rect 13170 13404 13176 13416
rect 13228 13404 13234 13456
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 10827 13348 10977 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 10965 13345 10977 13348
rect 11011 13376 11023 13379
rect 11609 13379 11667 13385
rect 11609 13376 11621 13379
rect 11011 13348 11284 13376
rect 11011 13345 11023 13348
rect 10965 13339 11023 13345
rect 11256 13252 11284 13348
rect 11348 13348 11621 13376
rect 10704 13212 11192 13240
rect 10134 13132 10140 13184
rect 10192 13172 10198 13184
rect 10704 13181 10732 13212
rect 10689 13175 10747 13181
rect 10689 13172 10701 13175
rect 10192 13144 10701 13172
rect 10192 13132 10198 13144
rect 10689 13141 10701 13144
rect 10735 13141 10747 13175
rect 10689 13135 10747 13141
rect 11054 13132 11060 13184
rect 11112 13132 11118 13184
rect 11164 13172 11192 13212
rect 11238 13200 11244 13252
rect 11296 13200 11302 13252
rect 11348 13172 11376 13348
rect 11609 13345 11621 13348
rect 11655 13376 11667 13379
rect 11701 13379 11759 13385
rect 11701 13376 11713 13379
rect 11655 13348 11713 13376
rect 11655 13345 11667 13348
rect 11609 13339 11667 13345
rect 11701 13345 11713 13348
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 12161 13379 12219 13385
rect 12161 13345 12173 13379
rect 12207 13345 12219 13379
rect 12161 13339 12219 13345
rect 12253 13379 12311 13385
rect 12253 13345 12265 13379
rect 12299 13376 12311 13379
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 12299 13348 12633 13376
rect 12299 13345 12311 13348
rect 12253 13339 12311 13345
rect 12621 13345 12633 13348
rect 12667 13376 12679 13379
rect 12805 13379 12863 13385
rect 12805 13376 12817 13379
rect 12667 13348 12817 13376
rect 12667 13345 12679 13348
rect 12621 13339 12679 13345
rect 12805 13345 12817 13348
rect 12851 13345 12863 13379
rect 12805 13339 12863 13345
rect 12897 13379 12955 13385
rect 12897 13345 12909 13379
rect 12943 13345 12955 13379
rect 12897 13339 12955 13345
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13345 13047 13379
rect 12989 13339 13047 13345
rect 11164 13144 11376 13172
rect 11790 13132 11796 13184
rect 11848 13132 11854 13184
rect 12912 13172 12940 13339
rect 13188 13308 13216 13404
rect 13357 13379 13415 13385
rect 13357 13345 13369 13379
rect 13403 13376 13415 13379
rect 13464 13376 13492 13472
rect 14016 13444 14044 13472
rect 13832 13416 14412 13444
rect 13832 13385 13860 13416
rect 13403 13348 13492 13376
rect 13817 13379 13875 13385
rect 13403 13345 13415 13348
rect 13357 13339 13415 13345
rect 13817 13345 13829 13379
rect 13863 13345 13875 13379
rect 13817 13339 13875 13345
rect 13909 13379 13967 13385
rect 13909 13345 13921 13379
rect 13955 13376 13967 13379
rect 13998 13376 14004 13388
rect 13955 13348 14004 13376
rect 13955 13345 13967 13348
rect 13909 13339 13967 13345
rect 13998 13336 14004 13348
rect 14056 13336 14062 13388
rect 14384 13385 14412 13416
rect 14369 13379 14427 13385
rect 14369 13345 14381 13379
rect 14415 13345 14427 13379
rect 14369 13339 14427 13345
rect 14645 13379 14703 13385
rect 14645 13345 14657 13379
rect 14691 13345 14703 13379
rect 14752 13376 14780 13472
rect 15289 13447 15347 13453
rect 15289 13413 15301 13447
rect 15335 13444 15347 13447
rect 16224 13444 16252 13475
rect 16482 13472 16488 13524
rect 16540 13512 16546 13524
rect 17313 13515 17371 13521
rect 16540 13484 16620 13512
rect 16540 13472 16546 13484
rect 15335 13416 15884 13444
rect 16224 13416 16528 13444
rect 15335 13413 15347 13416
rect 15289 13407 15347 13413
rect 15856 13385 15884 13416
rect 14921 13379 14979 13385
rect 14921 13376 14933 13379
rect 14752 13348 14933 13376
rect 14645 13339 14703 13345
rect 14921 13345 14933 13348
rect 14967 13376 14979 13379
rect 15197 13379 15255 13385
rect 15197 13376 15209 13379
rect 14967 13348 15209 13376
rect 14967 13345 14979 13348
rect 14921 13339 14979 13345
rect 15197 13345 15209 13348
rect 15243 13345 15255 13379
rect 15197 13339 15255 13345
rect 15473 13379 15531 13385
rect 15473 13345 15485 13379
rect 15519 13345 15531 13379
rect 15749 13379 15807 13385
rect 15749 13376 15761 13379
rect 15473 13339 15531 13345
rect 15672 13348 15761 13376
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13188 13280 13737 13308
rect 13725 13277 13737 13280
rect 13771 13308 13783 13311
rect 14660 13308 14688 13339
rect 13771 13280 14688 13308
rect 14737 13311 14795 13317
rect 13771 13277 13783 13280
rect 13725 13271 13783 13277
rect 14737 13277 14749 13311
rect 14783 13308 14795 13311
rect 15013 13311 15071 13317
rect 15013 13308 15025 13311
rect 14783 13280 15025 13308
rect 14783 13277 14795 13280
rect 14737 13271 14795 13277
rect 15013 13277 15025 13280
rect 15059 13308 15071 13311
rect 15488 13308 15516 13339
rect 15672 13320 15700 13348
rect 15749 13345 15761 13348
rect 15795 13345 15807 13379
rect 15749 13339 15807 13345
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13376 15899 13379
rect 16117 13379 16175 13385
rect 16117 13376 16129 13379
rect 15887 13348 16129 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 16117 13345 16129 13348
rect 16163 13376 16175 13379
rect 16298 13376 16304 13388
rect 16163 13348 16304 13376
rect 16163 13345 16175 13348
rect 16117 13339 16175 13345
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 15562 13308 15568 13320
rect 15059 13280 15568 13308
rect 15059 13277 15071 13280
rect 15013 13271 15071 13277
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 15654 13268 15660 13320
rect 15712 13268 15718 13320
rect 16500 13308 16528 13416
rect 16592 13385 16620 13484
rect 17313 13481 17325 13515
rect 17359 13512 17371 13515
rect 17770 13512 17776 13524
rect 17359 13484 17776 13512
rect 17359 13481 17371 13484
rect 17313 13475 17371 13481
rect 16577 13379 16635 13385
rect 16577 13345 16589 13379
rect 16623 13345 16635 13379
rect 16577 13339 16635 13345
rect 16669 13379 16727 13385
rect 16669 13345 16681 13379
rect 16715 13376 16727 13379
rect 17129 13379 17187 13385
rect 17129 13376 17141 13379
rect 16715 13348 17141 13376
rect 16715 13345 16727 13348
rect 16669 13339 16727 13345
rect 17129 13345 17141 13348
rect 17175 13376 17187 13379
rect 17328 13376 17356 13475
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 18969 13515 19027 13521
rect 18969 13481 18981 13515
rect 19015 13512 19027 13515
rect 19978 13512 19984 13524
rect 19015 13484 19984 13512
rect 19015 13481 19027 13484
rect 18969 13475 19027 13481
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 20993 13515 21051 13521
rect 20993 13481 21005 13515
rect 21039 13512 21051 13515
rect 21910 13512 21916 13524
rect 21039 13484 21916 13512
rect 21039 13481 21051 13484
rect 20993 13475 21051 13481
rect 21910 13472 21916 13484
rect 21968 13472 21974 13524
rect 18690 13444 18696 13456
rect 17604 13416 18696 13444
rect 17604 13385 17632 13416
rect 18690 13404 18696 13416
rect 18748 13404 18754 13456
rect 19429 13447 19487 13453
rect 19429 13413 19441 13447
rect 19475 13444 19487 13447
rect 20622 13444 20628 13456
rect 19475 13416 20628 13444
rect 19475 13413 19487 13416
rect 19429 13407 19487 13413
rect 20622 13404 20628 13416
rect 20680 13404 20686 13456
rect 17862 13385 17868 13388
rect 17175 13348 17356 13376
rect 17405 13379 17463 13385
rect 17175 13345 17187 13348
rect 17129 13339 17187 13345
rect 17405 13345 17417 13379
rect 17451 13345 17463 13379
rect 17405 13339 17463 13345
rect 17589 13379 17647 13385
rect 17589 13345 17601 13379
rect 17635 13345 17647 13379
rect 17845 13379 17868 13385
rect 17845 13376 17857 13379
rect 17589 13339 17647 13345
rect 17696 13348 17857 13376
rect 17420 13308 17448 13339
rect 17696 13308 17724 13348
rect 17845 13345 17857 13348
rect 17845 13339 17868 13345
rect 17862 13336 17868 13339
rect 17920 13336 17926 13388
rect 19518 13336 19524 13388
rect 19576 13336 19582 13388
rect 19610 13336 19616 13388
rect 19668 13336 19674 13388
rect 19869 13379 19927 13385
rect 19869 13376 19881 13379
rect 19720 13348 19881 13376
rect 16500 13280 17724 13308
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19720 13308 19748 13348
rect 19869 13345 19881 13348
rect 19915 13345 19927 13379
rect 19869 13339 19927 13345
rect 19484 13280 19748 13308
rect 19484 13268 19490 13280
rect 13449 13243 13507 13249
rect 13449 13209 13461 13243
rect 13495 13240 13507 13243
rect 14366 13240 14372 13252
rect 13495 13212 14372 13240
rect 13495 13209 13507 13212
rect 13449 13203 13507 13209
rect 14366 13200 14372 13212
rect 14424 13200 14430 13252
rect 13998 13172 14004 13184
rect 12912 13144 14004 13172
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 17037 13175 17095 13181
rect 17037 13172 17049 13175
rect 16816 13144 17049 13172
rect 16816 13132 16822 13144
rect 17037 13141 17049 13144
rect 17083 13141 17095 13175
rect 17037 13135 17095 13141
rect 552 13082 31372 13104
rect 552 13030 4250 13082
rect 4302 13030 4314 13082
rect 4366 13030 4378 13082
rect 4430 13030 4442 13082
rect 4494 13030 4506 13082
rect 4558 13030 11955 13082
rect 12007 13030 12019 13082
rect 12071 13030 12083 13082
rect 12135 13030 12147 13082
rect 12199 13030 12211 13082
rect 12263 13030 19660 13082
rect 19712 13030 19724 13082
rect 19776 13030 19788 13082
rect 19840 13030 19852 13082
rect 19904 13030 19916 13082
rect 19968 13030 27365 13082
rect 27417 13030 27429 13082
rect 27481 13030 27493 13082
rect 27545 13030 27557 13082
rect 27609 13030 27621 13082
rect 27673 13030 31372 13082
rect 552 13008 31372 13030
rect 10045 12971 10103 12977
rect 10045 12937 10057 12971
rect 10091 12968 10103 12971
rect 10778 12968 10784 12980
rect 10091 12940 10784 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11112 12940 11468 12968
rect 11112 12928 11118 12940
rect 11440 12832 11468 12940
rect 11514 12928 11520 12980
rect 11572 12968 11578 12980
rect 12897 12971 12955 12977
rect 12897 12968 12909 12971
rect 11572 12940 12909 12968
rect 11572 12928 11578 12940
rect 11440 12804 11744 12832
rect 11146 12724 11152 12776
rect 11204 12773 11210 12776
rect 11204 12764 11216 12773
rect 11204 12736 11284 12764
rect 11204 12727 11216 12736
rect 11204 12724 11210 12727
rect 11256 12696 11284 12736
rect 11330 12724 11336 12776
rect 11388 12764 11394 12776
rect 11716 12773 11744 12804
rect 11790 12792 11796 12844
rect 11848 12832 11854 12844
rect 11848 12804 12020 12832
rect 11848 12792 11854 12804
rect 11425 12767 11483 12773
rect 11425 12764 11437 12767
rect 11388 12736 11437 12764
rect 11388 12724 11394 12736
rect 11425 12733 11437 12736
rect 11471 12733 11483 12767
rect 11425 12727 11483 12733
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12764 11759 12767
rect 11882 12764 11888 12776
rect 11747 12736 11888 12764
rect 11747 12733 11759 12736
rect 11701 12727 11759 12733
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 11992 12773 12020 12804
rect 12728 12773 12756 12940
rect 12897 12937 12909 12940
rect 12943 12937 12955 12971
rect 12897 12931 12955 12937
rect 17957 12971 18015 12977
rect 17957 12937 17969 12971
rect 18003 12968 18015 12971
rect 18506 12968 18512 12980
rect 18003 12940 18512 12968
rect 18003 12937 18015 12940
rect 17957 12931 18015 12937
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 18598 12928 18604 12980
rect 18656 12968 18662 12980
rect 18785 12971 18843 12977
rect 18785 12968 18797 12971
rect 18656 12940 18797 12968
rect 18656 12928 18662 12940
rect 18785 12937 18797 12940
rect 18831 12937 18843 12971
rect 18785 12931 18843 12937
rect 19337 12971 19395 12977
rect 19337 12937 19349 12971
rect 19383 12968 19395 12971
rect 19426 12968 19432 12980
rect 19383 12940 19432 12968
rect 19383 12937 19395 12940
rect 19337 12931 19395 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 20438 12928 20444 12980
rect 20496 12928 20502 12980
rect 22005 12971 22063 12977
rect 22005 12937 22017 12971
rect 22051 12968 22063 12971
rect 28258 12968 28264 12980
rect 22051 12940 28264 12968
rect 22051 12937 22063 12940
rect 22005 12931 22063 12937
rect 28258 12928 28264 12940
rect 28316 12928 28322 12980
rect 28534 12928 28540 12980
rect 28592 12968 28598 12980
rect 31662 12968 31668 12980
rect 28592 12940 31668 12968
rect 28592 12928 28598 12940
rect 31662 12928 31668 12940
rect 31720 12928 31726 12980
rect 18690 12860 18696 12912
rect 18748 12860 18754 12912
rect 19518 12860 19524 12912
rect 19576 12900 19582 12912
rect 19613 12903 19671 12909
rect 19613 12900 19625 12903
rect 19576 12872 19625 12900
rect 19576 12860 19582 12872
rect 19613 12869 19625 12872
rect 19659 12900 19671 12903
rect 20162 12900 20168 12912
rect 19659 12872 20168 12900
rect 19659 12869 19671 12872
rect 19613 12863 19671 12869
rect 20162 12860 20168 12872
rect 20220 12860 20226 12912
rect 23569 12903 23627 12909
rect 23569 12869 23581 12903
rect 23615 12900 23627 12903
rect 27982 12900 27988 12912
rect 23615 12872 27988 12900
rect 23615 12869 23627 12872
rect 23569 12863 23627 12869
rect 27982 12860 27988 12872
rect 28040 12860 28046 12912
rect 14458 12792 14464 12844
rect 14516 12832 14522 12844
rect 14737 12835 14795 12841
rect 14737 12832 14749 12835
rect 14516 12804 14749 12832
rect 14516 12792 14522 12804
rect 14737 12801 14749 12804
rect 14783 12801 14795 12835
rect 18708 12832 18736 12860
rect 14737 12795 14795 12801
rect 17604 12804 18736 12832
rect 19168 12804 19840 12832
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12764 12035 12767
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 12023 12736 12265 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 12253 12733 12265 12736
rect 12299 12733 12311 12767
rect 12253 12727 12311 12733
rect 12713 12767 12771 12773
rect 12713 12733 12725 12767
rect 12759 12733 12771 12767
rect 12713 12727 12771 12733
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 16577 12767 16635 12773
rect 16577 12733 16589 12767
rect 16623 12764 16635 12767
rect 17604 12764 17632 12804
rect 18141 12767 18199 12773
rect 18141 12764 18153 12767
rect 16623 12736 17632 12764
rect 17972 12736 18153 12764
rect 16623 12733 16635 12736
rect 16577 12727 16635 12733
rect 12069 12699 12127 12705
rect 12069 12696 12081 12699
rect 11256 12668 12081 12696
rect 12069 12665 12081 12668
rect 12115 12696 12127 12699
rect 12820 12696 12848 12727
rect 12115 12668 12848 12696
rect 12115 12665 12127 12668
rect 12069 12659 12127 12665
rect 16482 12656 16488 12708
rect 16540 12656 16546 12708
rect 16844 12699 16902 12705
rect 16844 12665 16856 12699
rect 16890 12665 16902 12699
rect 16844 12659 16902 12665
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 11609 12631 11667 12637
rect 11609 12628 11621 12631
rect 10744 12600 11621 12628
rect 10744 12588 10750 12600
rect 11609 12597 11621 12600
rect 11655 12597 11667 12631
rect 11609 12591 11667 12597
rect 12345 12631 12403 12637
rect 12345 12597 12357 12631
rect 12391 12628 12403 12631
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 12391 12600 12633 12628
rect 12391 12597 12403 12600
rect 12345 12591 12403 12597
rect 12621 12597 12633 12600
rect 12667 12628 12679 12631
rect 13998 12628 14004 12640
rect 12667 12600 14004 12628
rect 12667 12597 12679 12600
rect 12621 12591 12679 12597
rect 13998 12588 14004 12600
rect 14056 12588 14062 12640
rect 16758 12588 16764 12640
rect 16816 12628 16822 12640
rect 16868 12628 16896 12659
rect 17972 12628 18000 12736
rect 18141 12733 18153 12736
rect 18187 12764 18199 12767
rect 18693 12767 18751 12773
rect 18693 12764 18705 12767
rect 18187 12736 18705 12764
rect 18187 12733 18199 12736
rect 18141 12727 18199 12733
rect 18693 12733 18705 12736
rect 18739 12733 18751 12767
rect 18693 12727 18751 12733
rect 18966 12724 18972 12776
rect 19024 12764 19030 12776
rect 19168 12773 19196 12804
rect 19812 12773 19840 12804
rect 19978 12792 19984 12844
rect 20036 12832 20042 12844
rect 20530 12832 20536 12844
rect 20036 12804 20536 12832
rect 20036 12792 20042 12804
rect 20530 12792 20536 12804
rect 20588 12832 20594 12844
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20588 12804 20637 12832
rect 20588 12792 20594 12804
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 19153 12767 19211 12773
rect 19153 12764 19165 12767
rect 19024 12736 19165 12764
rect 19024 12724 19030 12736
rect 19153 12733 19165 12736
rect 19199 12733 19211 12767
rect 19153 12727 19211 12733
rect 19429 12767 19487 12773
rect 19429 12733 19441 12767
rect 19475 12764 19487 12767
rect 19521 12767 19579 12773
rect 19521 12764 19533 12767
rect 19475 12736 19533 12764
rect 19475 12733 19487 12736
rect 19429 12727 19487 12733
rect 19521 12733 19533 12736
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12733 19855 12767
rect 20073 12767 20131 12773
rect 20073 12764 20085 12767
rect 19797 12727 19855 12733
rect 19904 12736 20085 12764
rect 18233 12699 18291 12705
rect 18233 12665 18245 12699
rect 18279 12696 18291 12699
rect 19061 12699 19119 12705
rect 19061 12696 19073 12699
rect 18279 12668 19073 12696
rect 18279 12665 18291 12668
rect 18233 12659 18291 12665
rect 19061 12665 19073 12668
rect 19107 12696 19119 12699
rect 19444 12696 19472 12727
rect 19107 12668 19472 12696
rect 19107 12665 19119 12668
rect 19061 12659 19119 12665
rect 19904 12640 19932 12736
rect 20073 12733 20085 12736
rect 20119 12764 20131 12767
rect 20349 12767 20407 12773
rect 20349 12764 20361 12767
rect 20119 12736 20361 12764
rect 20119 12733 20131 12736
rect 20073 12727 20131 12733
rect 20349 12733 20361 12736
rect 20395 12733 20407 12767
rect 20640 12764 20668 12795
rect 22186 12764 22192 12776
rect 20640 12736 22192 12764
rect 20349 12727 20407 12733
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 20438 12656 20444 12708
rect 20496 12696 20502 12708
rect 20870 12699 20928 12705
rect 20870 12696 20882 12699
rect 20496 12668 20882 12696
rect 20496 12656 20502 12668
rect 20870 12665 20882 12668
rect 20916 12665 20928 12699
rect 22434 12699 22492 12705
rect 22434 12696 22446 12699
rect 20870 12659 20928 12665
rect 22066 12668 22446 12696
rect 16816 12600 18000 12628
rect 16816 12588 16822 12600
rect 19886 12588 19892 12640
rect 19944 12588 19950 12640
rect 20162 12588 20168 12640
rect 20220 12628 20226 12640
rect 20622 12628 20628 12640
rect 20220 12600 20628 12628
rect 20220 12588 20226 12600
rect 20622 12588 20628 12600
rect 20680 12628 20686 12640
rect 22066 12628 22094 12668
rect 22434 12665 22446 12668
rect 22480 12665 22492 12699
rect 22434 12659 22492 12665
rect 20680 12600 22094 12628
rect 20680 12588 20686 12600
rect 552 12538 31531 12560
rect 552 12486 8102 12538
rect 8154 12486 8166 12538
rect 8218 12486 8230 12538
rect 8282 12486 8294 12538
rect 8346 12486 8358 12538
rect 8410 12486 15807 12538
rect 15859 12486 15871 12538
rect 15923 12486 15935 12538
rect 15987 12486 15999 12538
rect 16051 12486 16063 12538
rect 16115 12486 23512 12538
rect 23564 12486 23576 12538
rect 23628 12486 23640 12538
rect 23692 12486 23704 12538
rect 23756 12486 23768 12538
rect 23820 12486 31217 12538
rect 31269 12486 31281 12538
rect 31333 12486 31345 12538
rect 31397 12486 31409 12538
rect 31461 12486 31473 12538
rect 31525 12486 31531 12538
rect 552 12464 31531 12486
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 6972 12396 9045 12424
rect 6972 12384 6978 12396
rect 9033 12393 9045 12396
rect 9079 12393 9091 12427
rect 9033 12387 9091 12393
rect 11238 12384 11244 12436
rect 11296 12424 11302 12436
rect 11333 12427 11391 12433
rect 11333 12424 11345 12427
rect 11296 12396 11345 12424
rect 11296 12384 11302 12396
rect 11333 12393 11345 12396
rect 11379 12424 11391 12427
rect 11609 12427 11667 12433
rect 11609 12424 11621 12427
rect 11379 12396 11621 12424
rect 11379 12393 11391 12396
rect 11333 12387 11391 12393
rect 11609 12393 11621 12396
rect 11655 12393 11667 12427
rect 11609 12387 11667 12393
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 11977 12427 12035 12433
rect 11977 12424 11989 12427
rect 11848 12396 11989 12424
rect 11848 12384 11854 12396
rect 11977 12393 11989 12396
rect 12023 12393 12035 12427
rect 11977 12387 12035 12393
rect 12894 12384 12900 12436
rect 12952 12424 12958 12436
rect 13541 12427 13599 12433
rect 13541 12424 13553 12427
rect 12952 12396 13553 12424
rect 12952 12384 12958 12396
rect 13541 12393 13553 12396
rect 13587 12393 13599 12427
rect 13541 12387 13599 12393
rect 14826 12384 14832 12436
rect 14884 12424 14890 12436
rect 15105 12427 15163 12433
rect 15105 12424 15117 12427
rect 14884 12396 15117 12424
rect 14884 12384 14890 12396
rect 15105 12393 15117 12396
rect 15151 12393 15163 12427
rect 15105 12387 15163 12393
rect 15654 12384 15660 12436
rect 15712 12384 15718 12436
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12424 16359 12427
rect 16758 12424 16764 12436
rect 16347 12396 16764 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 18417 12427 18475 12433
rect 18417 12393 18429 12427
rect 18463 12424 18475 12427
rect 18690 12424 18696 12436
rect 18463 12396 18696 12424
rect 18463 12393 18475 12396
rect 18417 12387 18475 12393
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 19245 12427 19303 12433
rect 19245 12393 19257 12427
rect 19291 12424 19303 12427
rect 19886 12424 19892 12436
rect 19291 12396 19892 12424
rect 19291 12393 19303 12396
rect 19245 12387 19303 12393
rect 19886 12384 19892 12396
rect 19944 12384 19950 12436
rect 20438 12424 20444 12436
rect 20088 12396 20444 12424
rect 9692 12328 11468 12356
rect 9692 12300 9720 12328
rect 11440 12300 11468 12328
rect 11882 12316 11888 12368
rect 11940 12316 11946 12368
rect 14090 12356 14096 12368
rect 12176 12328 14096 12356
rect 9674 12248 9680 12300
rect 9732 12248 9738 12300
rect 10134 12248 10140 12300
rect 10192 12297 10198 12300
rect 10192 12288 10204 12297
rect 10781 12291 10839 12297
rect 10192 12260 10237 12288
rect 10192 12251 10204 12260
rect 10781 12257 10793 12291
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 10192 12248 10198 12251
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12220 10471 12223
rect 10502 12220 10508 12232
rect 10459 12192 10508 12220
rect 10459 12189 10471 12192
rect 10413 12183 10471 12189
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 10796 12152 10824 12251
rect 10962 12248 10968 12300
rect 11020 12248 11026 12300
rect 11422 12248 11428 12300
rect 11480 12248 11486 12300
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12257 11759 12291
rect 11900 12288 11928 12316
rect 12176 12297 12204 12328
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 11900 12260 12081 12288
rect 11701 12251 11759 12257
rect 12069 12257 12081 12260
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 11057 12155 11115 12161
rect 11057 12152 11069 12155
rect 10796 12124 11069 12152
rect 11057 12121 11069 12124
rect 11103 12152 11115 12155
rect 11716 12152 11744 12251
rect 12084 12220 12112 12251
rect 12250 12248 12256 12300
rect 12308 12288 12314 12300
rect 13740 12297 13768 12328
rect 14090 12316 14096 12328
rect 14148 12356 14154 12368
rect 14148 12328 14504 12356
rect 14148 12316 14154 12328
rect 14476 12300 14504 12328
rect 13998 12297 14004 12300
rect 12417 12291 12475 12297
rect 12417 12288 12429 12291
rect 12308 12260 12429 12288
rect 12308 12248 12314 12260
rect 12417 12257 12429 12260
rect 12463 12257 12475 12291
rect 12417 12251 12475 12257
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12257 13783 12291
rect 13992 12288 14004 12297
rect 13959 12260 14004 12288
rect 13725 12251 13783 12257
rect 13992 12251 14004 12260
rect 13998 12248 14004 12251
rect 14056 12248 14062 12300
rect 14458 12248 14464 12300
rect 14516 12248 14522 12300
rect 15562 12248 15568 12300
rect 15620 12248 15626 12300
rect 16206 12248 16212 12300
rect 16264 12248 16270 12300
rect 16482 12248 16488 12300
rect 16540 12288 16546 12300
rect 16945 12291 17003 12297
rect 16945 12288 16957 12291
rect 16540 12260 16957 12288
rect 16540 12248 16546 12260
rect 16945 12257 16957 12260
rect 16991 12288 17003 12291
rect 17586 12288 17592 12300
rect 16991 12260 17592 12288
rect 16991 12257 17003 12260
rect 16945 12251 17003 12257
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 19153 12291 19211 12297
rect 19153 12257 19165 12291
rect 19199 12288 19211 12291
rect 19426 12288 19432 12300
rect 19199 12260 19432 12288
rect 19199 12257 19211 12260
rect 19153 12251 19211 12257
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 19797 12291 19855 12297
rect 19797 12257 19809 12291
rect 19843 12288 19855 12291
rect 19889 12291 19947 12297
rect 19889 12288 19901 12291
rect 19843 12260 19901 12288
rect 19843 12257 19855 12260
rect 19797 12251 19855 12257
rect 19889 12257 19901 12260
rect 19935 12288 19947 12291
rect 20088 12288 20116 12396
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 22186 12384 22192 12436
rect 22244 12424 22250 12436
rect 22833 12427 22891 12433
rect 22833 12424 22845 12427
rect 22244 12396 22845 12424
rect 22244 12384 22250 12396
rect 22833 12393 22845 12396
rect 22879 12393 22891 12427
rect 22833 12387 22891 12393
rect 24765 12427 24823 12433
rect 24765 12393 24777 12427
rect 24811 12424 24823 12427
rect 28442 12424 28448 12436
rect 24811 12396 28448 12424
rect 24811 12393 24823 12396
rect 24765 12387 24823 12393
rect 19935 12260 20116 12288
rect 20165 12291 20223 12297
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 20165 12257 20177 12291
rect 20211 12257 20223 12291
rect 20165 12251 20223 12257
rect 12268 12220 12296 12248
rect 12084 12192 12296 12220
rect 11103 12124 11744 12152
rect 11103 12121 11115 12124
rect 11057 12115 11115 12121
rect 10686 12044 10692 12096
rect 10744 12044 10750 12096
rect 11716 12084 11744 12124
rect 19981 12155 20039 12161
rect 19981 12121 19993 12155
rect 20027 12152 20039 12155
rect 20180 12152 20208 12251
rect 20622 12248 20628 12300
rect 20680 12248 20686 12300
rect 20714 12248 20720 12300
rect 20772 12248 20778 12300
rect 21542 12248 21548 12300
rect 21600 12248 21606 12300
rect 22848 12288 22876 12387
rect 28442 12384 28448 12396
rect 28500 12384 28506 12436
rect 22922 12288 22928 12300
rect 22848 12260 22928 12288
rect 22922 12248 22928 12260
rect 22980 12288 22986 12300
rect 23385 12291 23443 12297
rect 23385 12288 23397 12291
rect 22980 12260 23397 12288
rect 22980 12248 22986 12260
rect 23385 12257 23397 12260
rect 23431 12257 23443 12291
rect 23641 12291 23699 12297
rect 23641 12288 23653 12291
rect 23385 12251 23443 12257
rect 23492 12260 23653 12288
rect 20809 12223 20867 12229
rect 20809 12189 20821 12223
rect 20855 12220 20867 12223
rect 23492 12220 23520 12260
rect 23641 12257 23653 12260
rect 23687 12257 23699 12291
rect 23641 12251 23699 12257
rect 20855 12192 23520 12220
rect 20855 12189 20867 12192
rect 20809 12183 20867 12189
rect 20346 12152 20352 12164
rect 20027 12124 20352 12152
rect 20027 12121 20039 12124
rect 19981 12115 20039 12121
rect 20346 12112 20352 12124
rect 20404 12152 20410 12164
rect 20533 12155 20591 12161
rect 20533 12152 20545 12155
rect 20404 12124 20545 12152
rect 20404 12112 20410 12124
rect 20533 12121 20545 12124
rect 20579 12121 20591 12155
rect 20533 12115 20591 12121
rect 12434 12084 12440 12096
rect 11716 12056 12440 12084
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 19518 12044 19524 12096
rect 19576 12084 19582 12096
rect 19705 12087 19763 12093
rect 19705 12084 19717 12087
rect 19576 12056 19717 12084
rect 19576 12044 19582 12056
rect 19705 12053 19717 12056
rect 19751 12053 19763 12087
rect 19705 12047 19763 12053
rect 20257 12087 20315 12093
rect 20257 12053 20269 12087
rect 20303 12084 20315 12087
rect 20622 12084 20628 12096
rect 20303 12056 20628 12084
rect 20303 12053 20315 12056
rect 20257 12047 20315 12053
rect 20622 12044 20628 12056
rect 20680 12084 20686 12096
rect 20824 12084 20852 12183
rect 20680 12056 20852 12084
rect 20680 12044 20686 12056
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 28258 12084 28264 12096
rect 21048 12056 28264 12084
rect 21048 12044 21054 12056
rect 28258 12044 28264 12056
rect 28316 12044 28322 12096
rect 552 11994 31372 12016
rect 552 11942 4250 11994
rect 4302 11942 4314 11994
rect 4366 11942 4378 11994
rect 4430 11942 4442 11994
rect 4494 11942 4506 11994
rect 4558 11942 11955 11994
rect 12007 11942 12019 11994
rect 12071 11942 12083 11994
rect 12135 11942 12147 11994
rect 12199 11942 12211 11994
rect 12263 11942 19660 11994
rect 19712 11942 19724 11994
rect 19776 11942 19788 11994
rect 19840 11942 19852 11994
rect 19904 11942 19916 11994
rect 19968 11942 27365 11994
rect 27417 11942 27429 11994
rect 27481 11942 27493 11994
rect 27545 11942 27557 11994
rect 27609 11942 27621 11994
rect 27673 11942 31372 11994
rect 552 11920 31372 11942
rect 9401 11883 9459 11889
rect 9401 11849 9413 11883
rect 9447 11880 9459 11883
rect 10134 11880 10140 11892
rect 9447 11852 10140 11880
rect 9447 11849 9459 11852
rect 9401 11843 9459 11849
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 11422 11840 11428 11892
rect 11480 11840 11486 11892
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 12400 11852 12725 11880
rect 12400 11840 12406 11852
rect 12713 11849 12725 11852
rect 12759 11849 12771 11883
rect 12713 11843 12771 11849
rect 15381 11883 15439 11889
rect 15381 11849 15393 11883
rect 15427 11880 15439 11883
rect 15470 11880 15476 11892
rect 15427 11852 15476 11880
rect 15427 11849 15439 11852
rect 15381 11843 15439 11849
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 18417 11883 18475 11889
rect 18417 11849 18429 11883
rect 18463 11880 18475 11883
rect 19334 11880 19340 11892
rect 18463 11852 19340 11880
rect 18463 11849 18475 11852
rect 18417 11843 18475 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 19518 11840 19524 11892
rect 19576 11840 19582 11892
rect 20346 11840 20352 11892
rect 20404 11840 20410 11892
rect 20622 11840 20628 11892
rect 20680 11840 20686 11892
rect 20898 11840 20904 11892
rect 20956 11880 20962 11892
rect 21913 11883 21971 11889
rect 21913 11880 21925 11883
rect 20956 11852 21925 11880
rect 20956 11840 20962 11852
rect 21913 11849 21925 11852
rect 21959 11880 21971 11883
rect 23569 11883 23627 11889
rect 21959 11852 22094 11880
rect 21959 11849 21971 11852
rect 21913 11843 21971 11849
rect 11440 11812 11468 11840
rect 11440 11784 12388 11812
rect 10686 11744 10692 11756
rect 9324 11716 10692 11744
rect 9030 11636 9036 11688
rect 9088 11636 9094 11688
rect 9324 11670 9352 11716
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 12360 11744 12388 11784
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 12492 11784 13032 11812
rect 12492 11772 12498 11784
rect 12268 11716 12940 11744
rect 12268 11685 12296 11716
rect 11793 11679 11851 11685
rect 9469 11673 9527 11679
rect 9469 11670 9481 11673
rect 9324 11642 9481 11670
rect 9469 11639 9481 11642
rect 9515 11639 9527 11673
rect 9469 11633 9527 11639
rect 9593 11673 9651 11679
rect 9593 11639 9605 11673
rect 9639 11639 9651 11673
rect 11793 11645 11805 11679
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11676 12587 11679
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12575 11648 12633 11676
rect 12575 11645 12587 11648
rect 12529 11639 12587 11645
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 9593 11633 9651 11639
rect 9122 11568 9128 11620
rect 9180 11568 9186 11620
rect 9140 11540 9168 11568
rect 9600 11540 9628 11633
rect 9858 11568 9864 11620
rect 9916 11568 9922 11620
rect 11808 11552 11836 11639
rect 12544 11608 12572 11639
rect 12406 11580 12572 11608
rect 9140 11512 9628 11540
rect 9674 11500 9680 11552
rect 9732 11500 9738 11552
rect 10502 11500 10508 11552
rect 10560 11540 10566 11552
rect 11149 11543 11207 11549
rect 11149 11540 11161 11543
rect 10560 11512 11161 11540
rect 10560 11500 10566 11512
rect 11149 11509 11161 11512
rect 11195 11540 11207 11543
rect 11330 11540 11336 11552
rect 11195 11512 11336 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 11790 11500 11796 11552
rect 11848 11500 11854 11552
rect 11885 11543 11943 11549
rect 11885 11509 11897 11543
rect 11931 11540 11943 11543
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11931 11512 12173 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 12161 11509 12173 11512
rect 12207 11540 12219 11543
rect 12406 11540 12434 11580
rect 12912 11552 12940 11716
rect 13004 11608 13032 11784
rect 18690 11704 18696 11756
rect 18748 11704 18754 11756
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11676 14059 11679
rect 14090 11676 14096 11688
rect 14047 11648 14096 11676
rect 14047 11645 14059 11648
rect 14001 11639 14059 11645
rect 14090 11636 14096 11648
rect 14148 11636 14154 11688
rect 17037 11679 17095 11685
rect 17037 11645 17049 11679
rect 17083 11676 17095 11679
rect 18046 11676 18052 11688
rect 17083 11648 18052 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 18046 11636 18052 11648
rect 18104 11676 18110 11688
rect 18708 11676 18736 11704
rect 18104 11648 18736 11676
rect 19536 11676 19564 11840
rect 20364 11685 20392 11840
rect 20640 11685 20668 11840
rect 20809 11815 20867 11821
rect 20809 11781 20821 11815
rect 20855 11812 20867 11815
rect 21637 11815 21695 11821
rect 21637 11812 21649 11815
rect 20855 11784 21649 11812
rect 20855 11781 20867 11784
rect 20809 11775 20867 11781
rect 21468 11685 21496 11784
rect 21637 11781 21649 11784
rect 21683 11781 21695 11815
rect 21637 11775 21695 11781
rect 19797 11679 19855 11685
rect 19797 11676 19809 11679
rect 19536 11648 19809 11676
rect 18104 11636 18110 11648
rect 19797 11645 19809 11648
rect 19843 11676 19855 11679
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 19843 11648 20085 11676
rect 19843 11645 19855 11648
rect 19797 11639 19855 11645
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 20073 11639 20131 11645
rect 20349 11679 20407 11685
rect 20349 11645 20361 11679
rect 20395 11645 20407 11679
rect 20349 11639 20407 11645
rect 20625 11679 20683 11685
rect 20625 11645 20637 11679
rect 20671 11676 20683 11679
rect 20717 11679 20775 11685
rect 20717 11676 20729 11679
rect 20671 11648 20729 11676
rect 20671 11645 20683 11648
rect 20625 11639 20683 11645
rect 20717 11645 20729 11648
rect 20763 11645 20775 11679
rect 21177 11679 21235 11685
rect 21177 11676 21189 11679
rect 20717 11639 20775 11645
rect 21008 11648 21189 11676
rect 14246 11611 14304 11617
rect 14246 11608 14258 11611
rect 13004 11580 14258 11608
rect 14246 11577 14258 11580
rect 14292 11577 14304 11611
rect 14246 11571 14304 11577
rect 17304 11611 17362 11617
rect 17304 11577 17316 11611
rect 17350 11608 17362 11611
rect 19981 11611 20039 11617
rect 19981 11608 19993 11611
rect 17350 11580 19993 11608
rect 17350 11577 17362 11580
rect 17304 11571 17362 11577
rect 19981 11577 19993 11580
rect 20027 11577 20039 11611
rect 20088 11608 20116 11639
rect 20533 11611 20591 11617
rect 20533 11608 20545 11611
rect 20088 11580 20545 11608
rect 19981 11571 20039 11577
rect 20533 11577 20545 11580
rect 20579 11577 20591 11611
rect 20533 11571 20591 11577
rect 21008 11608 21036 11648
rect 21177 11645 21189 11648
rect 21223 11645 21235 11679
rect 21177 11639 21235 11645
rect 21453 11679 21511 11685
rect 21453 11645 21465 11679
rect 21499 11645 21511 11679
rect 21453 11639 21511 11645
rect 21545 11679 21603 11685
rect 21545 11645 21557 11679
rect 21591 11645 21603 11679
rect 21652 11676 21680 11775
rect 21821 11679 21879 11685
rect 21821 11676 21833 11679
rect 21652 11648 21833 11676
rect 21545 11639 21603 11645
rect 21821 11645 21833 11648
rect 21867 11645 21879 11679
rect 21821 11639 21879 11645
rect 21560 11608 21588 11639
rect 22066 11620 22094 11852
rect 23569 11849 23581 11883
rect 23615 11880 23627 11883
rect 28534 11880 28540 11892
rect 23615 11852 28540 11880
rect 23615 11849 23627 11852
rect 23569 11843 23627 11849
rect 28534 11840 28540 11852
rect 28592 11840 28598 11892
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 21008 11580 21588 11608
rect 12207 11512 12434 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 12894 11500 12900 11552
rect 12952 11500 12958 11552
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 19705 11543 19763 11549
rect 19705 11540 19717 11543
rect 19392 11512 19717 11540
rect 19392 11500 19398 11512
rect 19705 11509 19717 11512
rect 19751 11509 19763 11543
rect 19996 11540 20024 11571
rect 20257 11543 20315 11549
rect 20257 11540 20269 11543
rect 19996 11512 20269 11540
rect 19705 11503 19763 11509
rect 20257 11509 20269 11512
rect 20303 11540 20315 11543
rect 21008 11540 21036 11580
rect 22002 11568 22008 11620
rect 22060 11608 22094 11620
rect 22434 11611 22492 11617
rect 22434 11608 22446 11611
rect 22060 11580 22446 11608
rect 22060 11568 22066 11580
rect 22434 11577 22446 11580
rect 22480 11577 22492 11611
rect 22434 11571 22492 11577
rect 20303 11512 21036 11540
rect 20303 11509 20315 11512
rect 20257 11503 20315 11509
rect 21082 11500 21088 11552
rect 21140 11500 21146 11552
rect 21358 11500 21364 11552
rect 21416 11500 21422 11552
rect 552 11450 31531 11472
rect 552 11398 8102 11450
rect 8154 11398 8166 11450
rect 8218 11398 8230 11450
rect 8282 11398 8294 11450
rect 8346 11398 8358 11450
rect 8410 11398 15807 11450
rect 15859 11398 15871 11450
rect 15923 11398 15935 11450
rect 15987 11398 15999 11450
rect 16051 11398 16063 11450
rect 16115 11398 23512 11450
rect 23564 11398 23576 11450
rect 23628 11398 23640 11450
rect 23692 11398 23704 11450
rect 23756 11398 23768 11450
rect 23820 11398 31217 11450
rect 31269 11398 31281 11450
rect 31333 11398 31345 11450
rect 31397 11398 31409 11450
rect 31461 11398 31473 11450
rect 31525 11398 31531 11450
rect 552 11376 31531 11398
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 8113 11339 8171 11345
rect 8113 11336 8125 11339
rect 6972 11308 8125 11336
rect 6972 11296 6978 11308
rect 8113 11305 8125 11308
rect 8159 11305 8171 11339
rect 8113 11299 8171 11305
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 9180 11308 9536 11336
rect 9180 11296 9186 11308
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 9226 11271 9284 11277
rect 9226 11268 9238 11271
rect 9088 11240 9238 11268
rect 9088 11228 9094 11240
rect 9226 11237 9238 11240
rect 9272 11237 9284 11271
rect 9226 11231 9284 11237
rect 9508 11200 9536 11308
rect 9674 11296 9680 11348
rect 9732 11336 9738 11348
rect 10321 11339 10379 11345
rect 10321 11336 10333 11339
rect 9732 11308 10333 11336
rect 9732 11296 9738 11308
rect 10321 11305 10333 11308
rect 10367 11305 10379 11339
rect 10321 11299 10379 11305
rect 10597 11339 10655 11345
rect 10597 11305 10609 11339
rect 10643 11336 10655 11339
rect 10962 11336 10968 11348
rect 10643 11308 10968 11336
rect 10643 11305 10655 11308
rect 10597 11299 10655 11305
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 9508 11172 9689 11200
rect 9677 11169 9689 11172
rect 9723 11200 9735 11203
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9723 11172 10057 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 10413 11203 10471 11209
rect 10192 11172 10364 11200
rect 10192 11160 10198 11172
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 10336 11132 10364 11172
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10612 11200 10640 11299
rect 10962 11296 10968 11308
rect 11020 11336 11026 11348
rect 11057 11339 11115 11345
rect 11057 11336 11069 11339
rect 11020 11308 11069 11336
rect 11020 11296 11026 11308
rect 11057 11305 11069 11308
rect 11103 11305 11115 11339
rect 11057 11299 11115 11305
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 11606 11336 11612 11348
rect 11379 11308 11612 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 14185 11339 14243 11345
rect 14185 11336 14197 11339
rect 13596 11308 14197 11336
rect 13596 11296 13602 11308
rect 14185 11305 14197 11308
rect 14231 11305 14243 11339
rect 14185 11299 14243 11305
rect 15749 11339 15807 11345
rect 15749 11305 15761 11339
rect 15795 11336 15807 11339
rect 16206 11336 16212 11348
rect 15795 11308 16212 11336
rect 15795 11305 15807 11308
rect 15749 11299 15807 11305
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 17402 11296 17408 11348
rect 17460 11336 17466 11348
rect 17497 11339 17555 11345
rect 17497 11336 17509 11339
rect 17460 11308 17509 11336
rect 17460 11296 17466 11308
rect 17497 11305 17509 11308
rect 17543 11305 17555 11339
rect 17497 11299 17555 11305
rect 20898 11296 20904 11348
rect 20956 11296 20962 11348
rect 20990 11296 20996 11348
rect 21048 11296 21054 11348
rect 21082 11296 21088 11348
rect 21140 11336 21146 11348
rect 21913 11339 21971 11345
rect 21913 11336 21925 11339
rect 21140 11308 21925 11336
rect 21140 11296 21146 11308
rect 21913 11305 21925 11308
rect 21959 11305 21971 11339
rect 22465 11339 22523 11345
rect 22465 11336 22477 11339
rect 21913 11299 21971 11305
rect 22112 11308 22477 11336
rect 11790 11228 11796 11280
rect 11848 11228 11854 11280
rect 20717 11271 20775 11277
rect 12820 11240 14136 11268
rect 10459 11172 10640 11200
rect 10689 11203 10747 11209
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10689 11169 10701 11203
rect 10735 11200 10747 11203
rect 10735 11172 10824 11200
rect 10735 11169 10747 11172
rect 10689 11163 10747 11169
rect 10796 11144 10824 11172
rect 10962 11160 10968 11212
rect 11020 11200 11026 11212
rect 11149 11203 11207 11209
rect 11149 11200 11161 11203
rect 11020 11172 11161 11200
rect 11020 11160 11026 11172
rect 11149 11169 11161 11172
rect 11195 11200 11207 11203
rect 11808 11200 11836 11228
rect 12820 11209 12848 11240
rect 14108 11212 14136 11240
rect 16132 11240 18092 11268
rect 12446 11203 12504 11209
rect 12446 11200 12458 11203
rect 11195 11172 12458 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 12446 11169 12458 11172
rect 12492 11169 12504 11203
rect 12446 11163 12504 11169
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11200 12771 11203
rect 12805 11203 12863 11209
rect 12805 11200 12817 11203
rect 12759 11172 12817 11200
rect 12759 11169 12771 11172
rect 12713 11163 12771 11169
rect 12805 11169 12817 11172
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13061 11203 13119 11209
rect 13061 11200 13073 11203
rect 12952 11172 13073 11200
rect 12952 11160 12958 11172
rect 13061 11169 13073 11172
rect 13107 11169 13119 11203
rect 13061 11163 13119 11169
rect 14090 11160 14096 11212
rect 14148 11200 14154 11212
rect 14642 11209 14648 11212
rect 14369 11203 14427 11209
rect 14369 11200 14381 11203
rect 14148 11172 14381 11200
rect 14148 11160 14154 11172
rect 14369 11169 14381 11172
rect 14415 11169 14427 11203
rect 14369 11163 14427 11169
rect 14636 11163 14648 11209
rect 14642 11160 14648 11163
rect 14700 11160 14706 11212
rect 16132 11209 16160 11240
rect 18064 11212 18092 11240
rect 20717 11237 20729 11271
rect 20763 11268 20775 11271
rect 21008 11268 21036 11296
rect 20763 11240 21036 11268
rect 20763 11237 20775 11240
rect 20717 11231 20775 11237
rect 16117 11203 16175 11209
rect 16117 11169 16129 11203
rect 16163 11169 16175 11203
rect 16373 11203 16431 11209
rect 16373 11200 16385 11203
rect 16117 11163 16175 11169
rect 16224 11172 16385 11200
rect 10778 11132 10784 11144
rect 9539 11104 9720 11132
rect 10336 11104 10784 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9692 11076 9720 11104
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 9674 11024 9680 11076
rect 9732 11024 9738 11076
rect 9769 11067 9827 11073
rect 9769 11033 9781 11067
rect 9815 11064 9827 11067
rect 10980 11064 11008 11160
rect 16224 11132 16252 11172
rect 16373 11169 16385 11172
rect 16419 11169 16431 11203
rect 16373 11163 16431 11169
rect 18046 11160 18052 11212
rect 18104 11160 18110 11212
rect 19061 11203 19119 11209
rect 19061 11169 19073 11203
rect 19107 11200 19119 11203
rect 20530 11200 20536 11212
rect 19107 11172 20536 11200
rect 19107 11169 19119 11172
rect 19061 11163 19119 11169
rect 20530 11160 20536 11172
rect 20588 11160 20594 11212
rect 20993 11203 21051 11209
rect 20993 11169 21005 11203
rect 21039 11200 21051 11203
rect 21100 11200 21128 11296
rect 21634 11228 21640 11280
rect 21692 11268 21698 11280
rect 22112 11268 22140 11308
rect 21692 11240 22140 11268
rect 21692 11228 21698 11240
rect 21269 11203 21327 11209
rect 21269 11200 21281 11203
rect 21039 11172 21281 11200
rect 21039 11169 21051 11172
rect 20993 11163 21051 11169
rect 21269 11169 21281 11172
rect 21315 11169 21327 11203
rect 21269 11163 21327 11169
rect 21358 11160 21364 11212
rect 21416 11200 21422 11212
rect 21545 11203 21603 11209
rect 21545 11200 21557 11203
rect 21416 11172 21557 11200
rect 21416 11160 21422 11172
rect 21545 11169 21557 11172
rect 21591 11200 21603 11203
rect 21821 11203 21879 11209
rect 21821 11200 21833 11203
rect 21591 11172 21833 11200
rect 21591 11169 21603 11172
rect 21545 11163 21603 11169
rect 21821 11169 21833 11172
rect 21867 11169 21879 11203
rect 21821 11163 21879 11169
rect 16132 11104 16252 11132
rect 16132 11064 16160 11104
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 21560 11132 21588 11163
rect 22002 11160 22008 11212
rect 22060 11200 22066 11212
rect 22281 11203 22339 11209
rect 22060 11160 22094 11200
rect 22281 11169 22293 11203
rect 22327 11198 22339 11203
rect 22388 11198 22416 11308
rect 22465 11305 22477 11308
rect 22511 11305 22523 11339
rect 22465 11299 22523 11305
rect 24305 11339 24363 11345
rect 24305 11305 24317 11339
rect 24351 11336 24363 11339
rect 28258 11336 28264 11348
rect 24351 11308 28264 11336
rect 24351 11305 24363 11308
rect 24305 11299 24363 11305
rect 28258 11296 28264 11308
rect 28316 11296 28322 11348
rect 22327 11170 22416 11198
rect 22557 11203 22615 11209
rect 22327 11169 22339 11170
rect 22281 11163 22339 11169
rect 22557 11169 22569 11203
rect 22603 11200 22615 11203
rect 22649 11203 22707 11209
rect 22649 11200 22661 11203
rect 22603 11172 22661 11200
rect 22603 11169 22615 11172
rect 22557 11163 22615 11169
rect 22649 11169 22661 11172
rect 22695 11169 22707 11203
rect 23181 11203 23239 11209
rect 23181 11200 23193 11203
rect 22649 11163 22707 11169
rect 22756 11172 23193 11200
rect 19392 11104 21588 11132
rect 22066 11132 22094 11160
rect 22572 11132 22600 11163
rect 22066 11104 22600 11132
rect 19392 11092 19398 11104
rect 9815 11036 11008 11064
rect 15304 11036 16160 11064
rect 21361 11067 21419 11073
rect 9815 11033 9827 11036
rect 9769 11027 9827 11033
rect 15304 11008 15332 11036
rect 21361 11033 21373 11067
rect 21407 11064 21419 11067
rect 22186 11064 22192 11076
rect 21407 11036 21956 11064
rect 21407 11033 21419 11036
rect 21361 11027 21419 11033
rect 15286 10956 15292 11008
rect 15344 10956 15350 11008
rect 21928 10996 21956 11036
rect 22066 11036 22192 11064
rect 22066 10996 22094 11036
rect 22186 11024 22192 11036
rect 22244 11064 22250 11076
rect 22756 11064 22784 11172
rect 23181 11169 23193 11172
rect 23227 11169 23239 11203
rect 23181 11163 23239 11169
rect 22922 11092 22928 11144
rect 22980 11092 22986 11144
rect 22244 11036 22784 11064
rect 22244 11024 22250 11036
rect 21928 10968 22094 10996
rect 22738 10956 22744 11008
rect 22796 10956 22802 11008
rect 552 10906 31372 10928
rect 552 10854 4250 10906
rect 4302 10854 4314 10906
rect 4366 10854 4378 10906
rect 4430 10854 4442 10906
rect 4494 10854 4506 10906
rect 4558 10854 11955 10906
rect 12007 10854 12019 10906
rect 12071 10854 12083 10906
rect 12135 10854 12147 10906
rect 12199 10854 12211 10906
rect 12263 10854 19660 10906
rect 19712 10854 19724 10906
rect 19776 10854 19788 10906
rect 19840 10854 19852 10906
rect 19904 10854 19916 10906
rect 19968 10854 27365 10906
rect 27417 10854 27429 10906
rect 27481 10854 27493 10906
rect 27545 10854 27557 10906
rect 27609 10854 27621 10906
rect 27673 10854 31372 10906
rect 552 10832 31372 10854
rect 9769 10795 9827 10801
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 9815 10764 10057 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 10045 10761 10057 10764
rect 10091 10792 10103 10795
rect 10134 10792 10140 10804
rect 10091 10764 10140 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 10321 10795 10379 10801
rect 10321 10761 10333 10795
rect 10367 10792 10379 10795
rect 10962 10792 10968 10804
rect 10367 10764 10968 10792
rect 10367 10761 10379 10764
rect 10321 10755 10379 10761
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 11204 10764 11897 10792
rect 11204 10752 11210 10764
rect 11885 10761 11897 10764
rect 11931 10761 11943 10795
rect 11885 10755 11943 10761
rect 18417 10795 18475 10801
rect 18417 10761 18429 10795
rect 18463 10792 18475 10795
rect 21266 10792 21272 10804
rect 18463 10764 21272 10792
rect 18463 10761 18475 10764
rect 18417 10755 18475 10761
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 9674 10684 9680 10736
rect 9732 10684 9738 10736
rect 14642 10684 14648 10736
rect 14700 10724 14706 10736
rect 15933 10727 15991 10733
rect 15933 10724 15945 10727
rect 14700 10696 15945 10724
rect 14700 10684 14706 10696
rect 15933 10693 15945 10696
rect 15979 10693 15991 10727
rect 15933 10687 15991 10693
rect 22005 10727 22063 10733
rect 22005 10693 22017 10727
rect 22051 10724 22063 10727
rect 22094 10724 22100 10736
rect 22051 10696 22100 10724
rect 22051 10693 22063 10696
rect 22005 10687 22063 10693
rect 22094 10684 22100 10696
rect 22152 10684 22158 10736
rect 22738 10684 22744 10736
rect 22796 10684 22802 10736
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9692 10656 9720 10684
rect 10502 10656 10508 10668
rect 9088 10628 9628 10656
rect 9692 10628 10508 10656
rect 9088 10616 9094 10628
rect 9600 10600 9628 10628
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 16574 10656 16580 10668
rect 15764 10628 16580 10656
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 9048 10560 9137 10588
rect 9048 10464 9076 10560
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9125 10551 9183 10557
rect 9582 10548 9588 10600
rect 9640 10548 9646 10600
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 9766 10588 9772 10600
rect 9723 10560 9772 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 10137 10591 10195 10597
rect 10137 10557 10149 10591
rect 10183 10588 10195 10591
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 10183 10560 10241 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 10229 10557 10241 10560
rect 10275 10557 10287 10591
rect 10229 10551 10287 10557
rect 14461 10591 14519 10597
rect 14461 10557 14473 10591
rect 14507 10557 14519 10591
rect 14461 10551 14519 10557
rect 15197 10591 15255 10597
rect 15197 10557 15209 10591
rect 15243 10588 15255 10591
rect 15286 10588 15292 10600
rect 15243 10560 15292 10588
rect 15243 10557 15255 10560
rect 15197 10551 15255 10557
rect 9217 10523 9275 10529
rect 9217 10489 9229 10523
rect 9263 10520 9275 10523
rect 9493 10523 9551 10529
rect 9493 10520 9505 10523
rect 9263 10492 9505 10520
rect 9263 10489 9275 10492
rect 9217 10483 9275 10489
rect 9493 10489 9505 10492
rect 9539 10520 9551 10523
rect 10152 10520 10180 10551
rect 9539 10492 10180 10520
rect 9539 10489 9551 10492
rect 9493 10483 9551 10489
rect 14476 10464 14504 10551
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 15764 10597 15792 10628
rect 16574 10616 16580 10628
rect 16632 10616 16638 10668
rect 18046 10616 18052 10668
rect 18104 10616 18110 10668
rect 22278 10616 22284 10668
rect 22336 10656 22342 10668
rect 22756 10656 22784 10684
rect 22336 10628 22784 10656
rect 22336 10616 22342 10628
rect 15749 10591 15807 10597
rect 15749 10557 15761 10591
rect 15795 10557 15807 10591
rect 15749 10551 15807 10557
rect 15841 10591 15899 10597
rect 15841 10557 15853 10591
rect 15887 10557 15899 10591
rect 15841 10551 15899 10557
rect 15856 10520 15884 10551
rect 15672 10492 15884 10520
rect 16592 10520 16620 10616
rect 17037 10591 17095 10597
rect 17037 10557 17049 10591
rect 17083 10588 17095 10591
rect 18064 10588 18092 10616
rect 17083 10560 18092 10588
rect 17083 10557 17095 10560
rect 17037 10551 17095 10557
rect 21634 10548 21640 10600
rect 21692 10548 21698 10600
rect 22097 10591 22155 10597
rect 22097 10557 22109 10591
rect 22143 10588 22155 10591
rect 22186 10588 22192 10600
rect 22143 10560 22192 10588
rect 22143 10557 22155 10560
rect 22097 10551 22155 10557
rect 22186 10548 22192 10560
rect 22244 10588 22250 10600
rect 22664 10597 22692 10628
rect 22373 10591 22431 10597
rect 22373 10588 22385 10591
rect 22244 10560 22385 10588
rect 22244 10548 22250 10560
rect 22373 10557 22385 10560
rect 22419 10557 22431 10591
rect 22373 10551 22431 10557
rect 22649 10591 22707 10597
rect 22649 10557 22661 10591
rect 22695 10557 22707 10591
rect 22649 10551 22707 10557
rect 22738 10548 22744 10600
rect 22796 10548 22802 10600
rect 17282 10523 17340 10529
rect 17282 10520 17294 10523
rect 16592 10492 17294 10520
rect 9030 10412 9036 10464
rect 9088 10412 9094 10464
rect 14366 10412 14372 10464
rect 14424 10412 14430 10464
rect 14458 10412 14464 10464
rect 14516 10412 14522 10464
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 15378 10452 15384 10464
rect 15335 10424 15384 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 15378 10412 15384 10424
rect 15436 10452 15442 10464
rect 15672 10461 15700 10492
rect 17282 10489 17294 10492
rect 17328 10489 17340 10523
rect 17282 10483 17340 10489
rect 21729 10523 21787 10529
rect 21729 10489 21741 10523
rect 21775 10520 21787 10523
rect 22002 10520 22008 10532
rect 21775 10492 22008 10520
rect 21775 10489 21787 10492
rect 21729 10483 21787 10489
rect 22002 10480 22008 10492
rect 22060 10520 22066 10532
rect 22557 10523 22615 10529
rect 22557 10520 22569 10523
rect 22060 10492 22569 10520
rect 22060 10480 22066 10492
rect 22557 10489 22569 10492
rect 22603 10489 22615 10523
rect 22557 10483 22615 10489
rect 15657 10455 15715 10461
rect 15657 10452 15669 10455
rect 15436 10424 15669 10452
rect 15436 10412 15442 10424
rect 15657 10421 15669 10424
rect 15703 10421 15715 10455
rect 15657 10415 15715 10421
rect 22186 10412 22192 10464
rect 22244 10452 22250 10464
rect 22830 10452 22836 10464
rect 22244 10424 22836 10452
rect 22244 10412 22250 10424
rect 22830 10412 22836 10424
rect 22888 10412 22894 10464
rect 552 10362 31531 10384
rect 552 10310 8102 10362
rect 8154 10310 8166 10362
rect 8218 10310 8230 10362
rect 8282 10310 8294 10362
rect 8346 10310 8358 10362
rect 8410 10310 15807 10362
rect 15859 10310 15871 10362
rect 15923 10310 15935 10362
rect 15987 10310 15999 10362
rect 16051 10310 16063 10362
rect 16115 10310 23512 10362
rect 23564 10310 23576 10362
rect 23628 10310 23640 10362
rect 23692 10310 23704 10362
rect 23756 10310 23768 10362
rect 23820 10310 31217 10362
rect 31269 10310 31281 10362
rect 31333 10310 31345 10362
rect 31397 10310 31409 10362
rect 31461 10310 31473 10362
rect 31525 10310 31531 10362
rect 552 10288 31531 10310
rect 7098 10208 7104 10260
rect 7156 10208 7162 10260
rect 9674 10248 9680 10260
rect 8496 10220 9680 10248
rect 8225 10115 8283 10121
rect 8225 10081 8237 10115
rect 8271 10112 8283 10115
rect 8386 10112 8392 10124
rect 8271 10084 8392 10112
rect 8271 10081 8283 10084
rect 8225 10075 8283 10081
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 8496 10121 8524 10220
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 9766 10208 9772 10260
rect 9824 10248 9830 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 9824 10220 9873 10248
rect 9824 10208 9830 10220
rect 9861 10217 9873 10220
rect 9907 10248 9919 10251
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 9907 10220 10149 10248
rect 9907 10217 9919 10220
rect 9861 10211 9919 10217
rect 10137 10217 10149 10220
rect 10183 10217 10195 10251
rect 10137 10211 10195 10217
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 15289 10251 15347 10257
rect 15289 10248 15301 10251
rect 14516 10220 15301 10248
rect 14516 10208 14522 10220
rect 15289 10217 15301 10220
rect 15335 10217 15347 10251
rect 15289 10211 15347 10217
rect 15378 10208 15384 10260
rect 15436 10208 15442 10260
rect 22186 10248 22192 10260
rect 21744 10220 22192 10248
rect 8757 10183 8815 10189
rect 8757 10149 8769 10183
rect 8803 10180 8815 10183
rect 9582 10180 9588 10192
rect 8803 10152 9588 10180
rect 8803 10149 8815 10152
rect 8757 10143 8815 10149
rect 9582 10140 9588 10152
rect 9640 10140 9646 10192
rect 9784 10180 9812 10208
rect 9692 10152 9812 10180
rect 14292 10152 14780 10180
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10081 8539 10115
rect 8481 10075 8539 10081
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 9692 10121 9720 10152
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8904 10084 9137 10112
rect 8904 10072 8910 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 9125 10075 9183 10081
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10081 9827 10115
rect 9769 10075 9827 10081
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10081 10287 10115
rect 14292 10112 14320 10152
rect 10229 10075 10287 10081
rect 12406 10084 14320 10112
rect 14553 10115 14611 10121
rect 8404 10044 8432 10072
rect 9030 10044 9036 10056
rect 8404 10016 9036 10044
rect 9030 10004 9036 10016
rect 9088 10044 9094 10056
rect 9784 10044 9812 10075
rect 9088 10016 9812 10044
rect 9088 10004 9094 10016
rect 9950 10004 9956 10056
rect 10008 10044 10014 10056
rect 10244 10044 10272 10075
rect 10008 10016 10272 10044
rect 10008 10004 10014 10016
rect 12406 9976 12434 10084
rect 14553 10081 14565 10115
rect 14599 10081 14611 10115
rect 14553 10075 14611 10081
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 13909 10047 13967 10053
rect 13909 10044 13921 10047
rect 13872 10016 13921 10044
rect 13872 10004 13878 10016
rect 13909 10013 13921 10016
rect 13955 10013 13967 10047
rect 13909 10007 13967 10013
rect 14182 10004 14188 10056
rect 14240 10004 14246 10056
rect 8496 9948 12434 9976
rect 14568 9976 14596 10075
rect 14642 10072 14648 10124
rect 14700 10072 14706 10124
rect 14752 10044 14780 10152
rect 15105 10115 15163 10121
rect 15105 10081 15117 10115
rect 15151 10112 15163 10115
rect 15286 10112 15292 10124
rect 15151 10084 15292 10112
rect 15151 10081 15163 10084
rect 15105 10075 15163 10081
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 15396 10121 15424 10208
rect 15381 10115 15439 10121
rect 15381 10081 15393 10115
rect 15427 10081 15439 10115
rect 15381 10075 15439 10081
rect 15657 10115 15715 10121
rect 15657 10081 15669 10115
rect 15703 10112 15715 10115
rect 15930 10112 15936 10124
rect 15703 10084 15936 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 16117 10115 16175 10121
rect 16117 10081 16129 10115
rect 16163 10081 16175 10115
rect 16117 10075 16175 10081
rect 16132 10044 16160 10075
rect 18046 10072 18052 10124
rect 18104 10072 18110 10124
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 21744 10121 21772 10220
rect 22186 10208 22192 10220
rect 22244 10208 22250 10260
rect 22278 10208 22284 10260
rect 22336 10208 22342 10260
rect 22741 10251 22799 10257
rect 22741 10217 22753 10251
rect 22787 10248 22799 10251
rect 22830 10248 22836 10260
rect 22787 10220 22836 10248
rect 22787 10217 22799 10220
rect 22741 10211 22799 10217
rect 22830 10208 22836 10220
rect 22888 10208 22894 10260
rect 24305 10251 24363 10257
rect 24305 10217 24317 10251
rect 24351 10248 24363 10251
rect 28258 10248 28264 10260
rect 24351 10220 28264 10248
rect 24351 10217 24363 10220
rect 24305 10211 24363 10217
rect 28258 10208 28264 10220
rect 28316 10208 28322 10260
rect 22296 10127 22324 10208
rect 23170 10183 23228 10189
rect 23170 10180 23182 10183
rect 22848 10152 23182 10180
rect 18581 10115 18639 10121
rect 18581 10112 18593 10115
rect 18196 10084 18593 10112
rect 18196 10072 18202 10084
rect 18581 10081 18593 10084
rect 18627 10081 18639 10115
rect 21453 10115 21511 10121
rect 21453 10112 21465 10115
rect 18581 10075 18639 10081
rect 21284 10084 21465 10112
rect 14752 10016 16160 10044
rect 18064 10044 18092 10072
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 18064 10016 18337 10044
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 14568 9948 14780 9976
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 8496 9908 8524 9948
rect 7248 9880 8524 9908
rect 7248 9868 7254 9880
rect 12618 9868 12624 9920
rect 12676 9868 12682 9920
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14458 9908 14464 9920
rect 13872 9880 14464 9908
rect 13872 9868 13878 9880
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 14752 9917 14780 9948
rect 14826 9936 14832 9988
rect 14884 9976 14890 9988
rect 15565 9979 15623 9985
rect 15565 9976 15577 9979
rect 14884 9948 15577 9976
rect 14884 9936 14890 9948
rect 15565 9945 15577 9948
rect 15611 9945 15623 9979
rect 15565 9939 15623 9945
rect 14737 9911 14795 9917
rect 14737 9877 14749 9911
rect 14783 9908 14795 9911
rect 14918 9908 14924 9920
rect 14783 9880 14924 9908
rect 14783 9877 14795 9880
rect 14737 9871 14795 9877
rect 14918 9868 14924 9880
rect 14976 9908 14982 9920
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14976 9880 15025 9908
rect 14976 9868 14982 9880
rect 15013 9877 15025 9880
rect 15059 9877 15071 9911
rect 15013 9871 15071 9877
rect 15286 9868 15292 9920
rect 15344 9908 15350 9920
rect 15838 9908 15844 9920
rect 15344 9880 15844 9908
rect 15344 9868 15350 9880
rect 15838 9868 15844 9880
rect 15896 9868 15902 9920
rect 17586 9868 17592 9920
rect 17644 9868 17650 9920
rect 18046 9868 18052 9920
rect 18104 9868 18110 9920
rect 19705 9911 19763 9917
rect 19705 9877 19717 9911
rect 19751 9908 19763 9911
rect 20898 9908 20904 9920
rect 19751 9880 20904 9908
rect 19751 9877 19763 9880
rect 19705 9871 19763 9877
rect 20898 9868 20904 9880
rect 20956 9868 20962 9920
rect 21284 9908 21312 10084
rect 21453 10081 21465 10084
rect 21499 10081 21511 10115
rect 21453 10075 21511 10081
rect 21729 10115 21787 10121
rect 21729 10081 21741 10115
rect 21775 10081 21787 10115
rect 21729 10075 21787 10081
rect 22002 10072 22008 10124
rect 22060 10121 22066 10124
rect 22281 10121 22339 10127
rect 22060 10112 22071 10121
rect 22060 10084 22232 10112
rect 22060 10075 22071 10084
rect 22060 10072 22066 10075
rect 21361 10047 21419 10053
rect 21361 10013 21373 10047
rect 21407 10044 21419 10047
rect 21818 10044 21824 10056
rect 21407 10016 21824 10044
rect 21407 10013 21419 10016
rect 21361 10007 21419 10013
rect 21818 10004 21824 10016
rect 21876 10004 21882 10056
rect 22204 10044 22232 10084
rect 22281 10087 22293 10121
rect 22327 10087 22339 10121
rect 22281 10081 22339 10087
rect 22370 10072 22376 10124
rect 22428 10072 22434 10124
rect 22848 10121 22876 10152
rect 23170 10149 23182 10152
rect 23216 10149 23228 10183
rect 23170 10143 23228 10149
rect 22833 10115 22891 10121
rect 22833 10081 22845 10115
rect 22879 10081 22891 10115
rect 22833 10075 22891 10081
rect 22848 10044 22876 10075
rect 22922 10072 22928 10124
rect 22980 10072 22986 10124
rect 22204 10016 22876 10044
rect 21637 9979 21695 9985
rect 21637 9945 21649 9979
rect 21683 9976 21695 9979
rect 22465 9979 22523 9985
rect 22465 9976 22477 9979
rect 21683 9948 22477 9976
rect 21683 9945 21695 9948
rect 21637 9939 21695 9945
rect 22465 9945 22477 9948
rect 22511 9945 22523 9979
rect 22465 9939 22523 9945
rect 22738 9936 22744 9988
rect 22796 9936 22802 9988
rect 21913 9911 21971 9917
rect 21913 9908 21925 9911
rect 21284 9880 21925 9908
rect 21913 9877 21925 9880
rect 21959 9908 21971 9911
rect 22094 9908 22100 9920
rect 21959 9880 22100 9908
rect 21959 9877 21971 9880
rect 21913 9871 21971 9877
rect 22094 9868 22100 9880
rect 22152 9868 22158 9920
rect 22186 9868 22192 9920
rect 22244 9908 22250 9920
rect 22756 9908 22784 9936
rect 22244 9880 22784 9908
rect 22244 9868 22250 9880
rect 552 9818 31372 9840
rect 552 9766 4250 9818
rect 4302 9766 4314 9818
rect 4366 9766 4378 9818
rect 4430 9766 4442 9818
rect 4494 9766 4506 9818
rect 4558 9766 11955 9818
rect 12007 9766 12019 9818
rect 12071 9766 12083 9818
rect 12135 9766 12147 9818
rect 12199 9766 12211 9818
rect 12263 9766 19660 9818
rect 19712 9766 19724 9818
rect 19776 9766 19788 9818
rect 19840 9766 19852 9818
rect 19904 9766 19916 9818
rect 19968 9766 27365 9818
rect 27417 9766 27429 9818
rect 27481 9766 27493 9818
rect 27545 9766 27557 9818
rect 27609 9766 27621 9818
rect 27673 9766 31372 9818
rect 552 9744 31372 9766
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 8481 9707 8539 9713
rect 8481 9704 8493 9707
rect 8444 9676 8493 9704
rect 8444 9664 8450 9676
rect 8481 9673 8493 9676
rect 8527 9673 8539 9707
rect 8481 9667 8539 9673
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 9125 9707 9183 9713
rect 9125 9704 9137 9707
rect 8904 9676 9137 9704
rect 8904 9664 8910 9676
rect 9125 9673 9137 9676
rect 9171 9673 9183 9707
rect 9125 9667 9183 9673
rect 14366 9664 14372 9716
rect 14424 9704 14430 9716
rect 14553 9707 14611 9713
rect 14553 9704 14565 9707
rect 14424 9676 14565 9704
rect 14424 9664 14430 9676
rect 14553 9673 14565 9676
rect 14599 9673 14611 9707
rect 14553 9667 14611 9673
rect 15930 9664 15936 9716
rect 15988 9704 15994 9716
rect 16117 9707 16175 9713
rect 16117 9704 16129 9707
rect 15988 9676 16129 9704
rect 15988 9664 15994 9676
rect 16117 9673 16129 9676
rect 16163 9704 16175 9707
rect 16393 9707 16451 9713
rect 16393 9704 16405 9707
rect 16163 9676 16405 9704
rect 16163 9673 16175 9676
rect 16117 9667 16175 9673
rect 16393 9673 16405 9676
rect 16439 9673 16451 9707
rect 16393 9667 16451 9673
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 16669 9707 16727 9713
rect 16669 9704 16681 9707
rect 16632 9676 16681 9704
rect 16632 9664 16638 9676
rect 16669 9673 16681 9676
rect 16715 9704 16727 9707
rect 17681 9707 17739 9713
rect 17681 9704 17693 9707
rect 16715 9676 17693 9704
rect 16715 9673 16727 9676
rect 16669 9667 16727 9673
rect 17681 9673 17693 9676
rect 17727 9673 17739 9707
rect 17681 9667 17739 9673
rect 18046 9664 18052 9716
rect 18104 9664 18110 9716
rect 20898 9664 20904 9716
rect 20956 9704 20962 9716
rect 31662 9704 31668 9716
rect 20956 9676 31668 9704
rect 20956 9664 20962 9676
rect 31662 9664 31668 9676
rect 31720 9664 31726 9716
rect 8220 9608 9260 9636
rect 8220 9509 8248 9608
rect 9232 9512 9260 9608
rect 9766 9596 9772 9648
rect 9824 9596 9830 9648
rect 13814 9636 13820 9648
rect 13280 9608 13820 9636
rect 12986 9528 12992 9580
rect 13044 9528 13050 9580
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9469 8263 9503
rect 8205 9463 8263 9469
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9469 8631 9503
rect 8573 9463 8631 9469
rect 8113 9435 8171 9441
rect 8113 9401 8125 9435
rect 8159 9432 8171 9435
rect 8478 9432 8484 9444
rect 8159 9404 8484 9432
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 8478 9392 8484 9404
rect 8536 9432 8542 9444
rect 8588 9432 8616 9463
rect 8846 9460 8852 9512
rect 8904 9500 8910 9512
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8904 9472 8953 9500
rect 8904 9460 8910 9472
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 9214 9460 9220 9512
rect 9272 9460 9278 9512
rect 13280 9509 13308 9608
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14384 9568 14412 9664
rect 16592 9568 16620 9664
rect 17221 9639 17279 9645
rect 17221 9605 17233 9639
rect 17267 9636 17279 9639
rect 18064 9636 18092 9664
rect 17267 9608 18092 9636
rect 17267 9605 17279 9608
rect 17221 9599 17279 9605
rect 14384 9540 15056 9568
rect 14384 9509 14412 9540
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9469 9367 9503
rect 10882 9503 10940 9509
rect 10882 9500 10894 9503
rect 9309 9463 9367 9469
rect 9968 9472 10894 9500
rect 9324 9432 9352 9463
rect 8536 9404 9352 9432
rect 8536 9392 8542 9404
rect 9968 9376 9996 9472
rect 10882 9469 10894 9472
rect 10928 9469 10940 9503
rect 10882 9463 10940 9469
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9469 11207 9503
rect 11149 9463 11207 9469
rect 13265 9503 13323 9509
rect 13265 9469 13277 9503
rect 13311 9469 13323 9503
rect 13265 9463 13323 9469
rect 13541 9503 13599 9509
rect 13541 9469 13553 9503
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 11164 9432 11192 9463
rect 10796 9404 11192 9432
rect 12744 9435 12802 9441
rect 10796 9376 10824 9404
rect 12744 9401 12756 9435
rect 12790 9432 12802 9435
rect 12790 9404 13124 9432
rect 12790 9401 12802 9404
rect 12744 9395 12802 9401
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 8904 9336 9413 9364
rect 8904 9324 8910 9336
rect 9401 9333 9413 9336
rect 9447 9364 9459 9367
rect 9950 9364 9956 9376
rect 9447 9336 9956 9364
rect 9447 9333 9459 9336
rect 9401 9327 9459 9333
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10778 9324 10784 9376
rect 10836 9324 10842 9376
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 11296 9336 11621 9364
rect 11296 9324 11302 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 13096 9364 13124 9404
rect 13170 9392 13176 9444
rect 13228 9432 13234 9444
rect 13556 9432 13584 9463
rect 14642 9460 14648 9512
rect 14700 9460 14706 9512
rect 14918 9460 14924 9512
rect 14976 9460 14982 9512
rect 15028 9509 15056 9540
rect 16224 9540 16620 9568
rect 16224 9509 16252 9540
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9469 15071 9503
rect 15013 9463 15071 9469
rect 16209 9503 16267 9509
rect 16209 9469 16221 9503
rect 16255 9469 16267 9503
rect 16209 9463 16267 9469
rect 16485 9503 16543 9509
rect 16485 9469 16497 9503
rect 16531 9469 16543 9503
rect 16485 9463 16543 9469
rect 16761 9503 16819 9509
rect 16761 9469 16773 9503
rect 16807 9500 16819 9503
rect 17037 9503 17095 9509
rect 17037 9500 17049 9503
rect 16807 9472 17049 9500
rect 16807 9469 16819 9472
rect 16761 9463 16819 9469
rect 17037 9469 17049 9472
rect 17083 9500 17095 9503
rect 17236 9500 17264 9599
rect 17328 9540 18368 9568
rect 17328 9512 17356 9540
rect 17083 9472 17264 9500
rect 17083 9469 17095 9472
rect 17037 9463 17095 9469
rect 15105 9435 15163 9441
rect 15105 9432 15117 9435
rect 13228 9404 13584 9432
rect 13648 9404 15117 9432
rect 13228 9392 13234 9404
rect 13648 9376 13676 9404
rect 15105 9401 15117 9404
rect 15151 9401 15163 9435
rect 16500 9432 16528 9463
rect 17310 9460 17316 9512
rect 17368 9460 17374 9512
rect 18340 9509 18368 9540
rect 17773 9503 17831 9509
rect 17773 9469 17785 9503
rect 17819 9500 17831 9503
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17819 9472 18061 9500
rect 17819 9469 17831 9472
rect 17773 9463 17831 9469
rect 18049 9469 18061 9472
rect 18095 9500 18107 9503
rect 18325 9503 18383 9509
rect 18095 9472 18276 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 17957 9435 18015 9441
rect 17957 9432 17969 9435
rect 16500 9404 17969 9432
rect 15105 9395 15163 9401
rect 17957 9401 17969 9404
rect 18003 9432 18015 9435
rect 18138 9432 18144 9444
rect 18003 9404 18144 9432
rect 18003 9401 18015 9404
rect 17957 9395 18015 9401
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18248 9441 18276 9472
rect 18325 9469 18337 9503
rect 18371 9469 18383 9503
rect 18325 9463 18383 9469
rect 18877 9503 18935 9509
rect 18877 9469 18889 9503
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9432 18291 9435
rect 18785 9435 18843 9441
rect 18785 9432 18797 9435
rect 18279 9404 18797 9432
rect 18279 9401 18291 9404
rect 18233 9395 18291 9401
rect 18785 9401 18797 9404
rect 18831 9401 18843 9435
rect 18892 9432 18920 9463
rect 18966 9460 18972 9512
rect 19024 9460 19030 9512
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 20898 9500 20904 9512
rect 19392 9472 20904 9500
rect 19392 9460 19398 9472
rect 20898 9460 20904 9472
rect 20956 9500 20962 9512
rect 22005 9503 22063 9509
rect 22005 9500 22017 9503
rect 20956 9472 22017 9500
rect 20956 9460 20962 9472
rect 22005 9469 22017 9472
rect 22051 9469 22063 9503
rect 28258 9500 28264 9512
rect 22005 9463 22063 9469
rect 22204 9472 28264 9500
rect 19426 9432 19432 9444
rect 18892 9404 19432 9432
rect 18785 9395 18843 9401
rect 19426 9392 19432 9404
rect 19484 9432 19490 9444
rect 19582 9435 19640 9441
rect 19582 9432 19594 9435
rect 19484 9404 19594 9432
rect 19484 9392 19490 9404
rect 19582 9401 19594 9404
rect 19628 9401 19640 9435
rect 19582 9395 19640 9401
rect 13262 9364 13268 9376
rect 13096 9336 13268 9364
rect 11609 9327 11667 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13630 9324 13636 9376
rect 13688 9324 13694 9376
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14277 9367 14335 9373
rect 14277 9364 14289 9367
rect 13964 9336 14289 9364
rect 13964 9324 13970 9336
rect 14277 9333 14289 9336
rect 14323 9364 14335 9367
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 14323 9336 14841 9364
rect 14323 9333 14335 9336
rect 14277 9327 14335 9333
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 15838 9324 15844 9376
rect 15896 9364 15902 9376
rect 16945 9367 17003 9373
rect 16945 9364 16957 9367
rect 15896 9336 16957 9364
rect 15896 9324 15902 9336
rect 16945 9333 16957 9336
rect 16991 9333 17003 9367
rect 18156 9364 18184 9392
rect 19061 9367 19119 9373
rect 19061 9364 19073 9367
rect 18156 9336 19073 9364
rect 16945 9327 17003 9333
rect 19061 9333 19073 9336
rect 19107 9333 19119 9367
rect 19061 9327 19119 9333
rect 20717 9367 20775 9373
rect 20717 9333 20729 9367
rect 20763 9364 20775 9367
rect 22204 9364 22232 9472
rect 28258 9460 28264 9472
rect 28316 9460 28322 9512
rect 22278 9441 22284 9444
rect 22272 9395 22284 9441
rect 22336 9432 22342 9444
rect 22336 9404 22372 9432
rect 22278 9392 22284 9395
rect 22336 9392 22342 9404
rect 20763 9336 22232 9364
rect 20763 9333 20775 9336
rect 20717 9327 20775 9333
rect 23382 9324 23388 9376
rect 23440 9324 23446 9376
rect 552 9274 31531 9296
rect 552 9222 8102 9274
rect 8154 9222 8166 9274
rect 8218 9222 8230 9274
rect 8282 9222 8294 9274
rect 8346 9222 8358 9274
rect 8410 9222 15807 9274
rect 15859 9222 15871 9274
rect 15923 9222 15935 9274
rect 15987 9222 15999 9274
rect 16051 9222 16063 9274
rect 16115 9222 23512 9274
rect 23564 9222 23576 9274
rect 23628 9222 23640 9274
rect 23692 9222 23704 9274
rect 23756 9222 23768 9274
rect 23820 9222 31217 9274
rect 31269 9222 31281 9274
rect 31333 9222 31345 9274
rect 31397 9222 31409 9274
rect 31461 9222 31473 9274
rect 31525 9222 31531 9274
rect 552 9200 31531 9222
rect 8297 9163 8355 9169
rect 8297 9129 8309 9163
rect 8343 9160 8355 9163
rect 8478 9160 8484 9172
rect 8343 9132 8484 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 8846 9120 8852 9172
rect 8904 9120 8910 9172
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9214 9160 9220 9172
rect 9171 9132 9220 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 12989 9163 13047 9169
rect 12989 9129 13001 9163
rect 13035 9160 13047 9163
rect 13170 9160 13176 9172
rect 13035 9132 13176 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 7868 9095 7926 9101
rect 7868 9061 7880 9095
rect 7914 9092 7926 9095
rect 9232 9092 9260 9120
rect 10514 9095 10572 9101
rect 10514 9092 10526 9095
rect 7914 9064 8432 9092
rect 9232 9064 10526 9092
rect 7914 9061 7926 9064
rect 7868 9055 7926 9061
rect 8404 9036 8432 9064
rect 10514 9061 10526 9064
rect 10560 9061 10572 9095
rect 10514 9055 10572 9061
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 8113 9027 8171 9033
rect 8113 9024 8125 9027
rect 8076 8996 8125 9024
rect 8076 8984 8082 8996
rect 8113 8993 8125 8996
rect 8159 8993 8171 9027
rect 8113 8987 8171 8993
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 8481 9027 8539 9033
rect 8481 9024 8493 9027
rect 8444 8996 8493 9024
rect 8444 8984 8450 8996
rect 8481 8993 8493 8996
rect 8527 8993 8539 9027
rect 8941 9027 8999 9033
rect 8941 9024 8953 9027
rect 8481 8987 8539 8993
rect 8680 8996 8953 9024
rect 6730 8848 6736 8900
rect 6788 8848 6794 8900
rect 8680 8832 8708 8996
rect 8941 8993 8953 8996
rect 8987 9024 8999 9027
rect 9033 9027 9091 9033
rect 9033 9024 9045 9027
rect 8987 8996 9045 9024
rect 8987 8993 8999 8996
rect 8941 8987 8999 8993
rect 9033 8993 9045 8996
rect 9079 8993 9091 9027
rect 9033 8987 9091 8993
rect 12805 9027 12863 9033
rect 12805 8993 12817 9027
rect 12851 9024 12863 9027
rect 13004 9024 13032 9123
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 13630 9120 13636 9172
rect 13688 9160 13694 9172
rect 17957 9163 18015 9169
rect 13688 9132 14136 9160
rect 13688 9120 13694 9132
rect 13906 9092 13912 9104
rect 13464 9064 13912 9092
rect 12851 8996 13032 9024
rect 13089 9027 13147 9033
rect 12851 8993 12863 8996
rect 12805 8987 12863 8993
rect 13089 8993 13101 9027
rect 13135 9024 13147 9027
rect 13262 9024 13268 9036
rect 13135 8996 13268 9024
rect 13135 8993 13147 8996
rect 13089 8987 13147 8993
rect 13262 8984 13268 8996
rect 13320 9024 13326 9036
rect 13464 9024 13492 9064
rect 13832 9033 13860 9064
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 14108 9033 14136 9132
rect 17957 9129 17969 9163
rect 18003 9160 18015 9163
rect 18322 9160 18328 9172
rect 18003 9132 18328 9160
rect 18003 9129 18015 9132
rect 17957 9123 18015 9129
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 18785 9163 18843 9169
rect 18785 9160 18797 9163
rect 18432 9132 18797 9160
rect 16476 9095 16534 9101
rect 16476 9061 16488 9095
rect 16522 9092 16534 9095
rect 17310 9092 17316 9104
rect 16522 9064 17316 9092
rect 16522 9061 16534 9064
rect 16476 9055 16534 9061
rect 17310 9052 17316 9064
rect 17368 9092 17374 9104
rect 18233 9095 18291 9101
rect 18233 9092 18245 9095
rect 17368 9064 18245 9092
rect 17368 9052 17374 9064
rect 18233 9061 18245 9064
rect 18279 9092 18291 9095
rect 18432 9092 18460 9132
rect 18785 9129 18797 9132
rect 18831 9129 18843 9163
rect 18785 9123 18843 9129
rect 18966 9120 18972 9172
rect 19024 9160 19030 9172
rect 19061 9163 19119 9169
rect 19061 9160 19073 9163
rect 19024 9132 19073 9160
rect 19024 9120 19030 9132
rect 19061 9129 19073 9132
rect 19107 9129 19119 9163
rect 19061 9123 19119 9129
rect 19337 9163 19395 9169
rect 19337 9129 19349 9163
rect 19383 9160 19395 9163
rect 19426 9160 19432 9172
rect 19383 9132 19432 9160
rect 19383 9129 19395 9132
rect 19337 9123 19395 9129
rect 18279 9064 18460 9092
rect 18509 9095 18567 9101
rect 18279 9061 18291 9064
rect 18233 9055 18291 9061
rect 18509 9061 18521 9095
rect 18555 9092 18567 9095
rect 18984 9092 19012 9120
rect 19352 9092 19380 9123
rect 19426 9120 19432 9132
rect 19484 9160 19490 9172
rect 19889 9163 19947 9169
rect 19889 9160 19901 9163
rect 19484 9132 19901 9160
rect 19484 9120 19490 9132
rect 19889 9129 19901 9132
rect 19935 9129 19947 9163
rect 19889 9123 19947 9129
rect 20070 9120 20076 9172
rect 20128 9120 20134 9172
rect 20088 9092 20116 9120
rect 18555 9064 19012 9092
rect 18555 9061 18567 9064
rect 18509 9055 18567 9061
rect 13320 8996 13492 9024
rect 13541 9027 13599 9033
rect 13320 8984 13326 8996
rect 13541 8993 13553 9027
rect 13587 8993 13599 9027
rect 13541 8987 13599 8993
rect 13817 9027 13875 9033
rect 13817 8993 13829 9027
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 14093 9027 14151 9033
rect 14093 8993 14105 9027
rect 14139 9024 14151 9027
rect 14369 9027 14427 9033
rect 14369 9024 14381 9027
rect 14139 8996 14381 9024
rect 14139 8993 14151 8996
rect 14093 8987 14151 8993
rect 14369 8993 14381 8996
rect 14415 9024 14427 9027
rect 14717 9027 14775 9033
rect 14717 9024 14729 9027
rect 14415 8996 14729 9024
rect 14415 8993 14427 8996
rect 14369 8987 14427 8993
rect 14717 8993 14729 8996
rect 14763 8993 14775 9027
rect 18049 9027 18107 9033
rect 18049 9024 18061 9027
rect 14717 8987 14775 8993
rect 17888 8996 18061 9024
rect 10778 8916 10784 8968
rect 10836 8916 10842 8968
rect 12713 8891 12771 8897
rect 12713 8857 12725 8891
rect 12759 8888 12771 8891
rect 13170 8888 13176 8900
rect 12759 8860 13176 8888
rect 12759 8857 12771 8860
rect 12713 8851 12771 8857
rect 13170 8848 13176 8860
rect 13228 8888 13234 8900
rect 13449 8891 13507 8897
rect 13449 8888 13461 8891
rect 13228 8860 13461 8888
rect 13228 8848 13234 8860
rect 13449 8857 13461 8860
rect 13495 8857 13507 8891
rect 13556 8888 13584 8987
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 13556 8860 13768 8888
rect 13449 8851 13507 8857
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 8662 8820 8668 8832
rect 8619 8792 8668 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 9398 8780 9404 8832
rect 9456 8780 9462 8832
rect 13740 8829 13768 8860
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 13998 8820 14004 8832
rect 13771 8792 14004 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 13998 8780 14004 8792
rect 14056 8780 14062 8832
rect 14274 8780 14280 8832
rect 14332 8780 14338 8832
rect 14476 8820 14504 8919
rect 16206 8916 16212 8968
rect 16264 8916 16270 8968
rect 17888 8888 17916 8996
rect 18049 8993 18061 8996
rect 18095 8993 18107 9027
rect 18049 8987 18107 8993
rect 18322 8984 18328 9036
rect 18380 8984 18386 9036
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 9024 18659 9027
rect 18782 9024 18788 9036
rect 18647 8996 18788 9024
rect 18647 8993 18659 8996
rect 18601 8987 18659 8993
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 18877 9027 18935 9033
rect 18877 8993 18889 9027
rect 18923 9024 18935 9027
rect 18984 9024 19012 9064
rect 19168 9064 19380 9092
rect 19720 9064 20116 9092
rect 19168 9033 19196 9064
rect 19720 9033 19748 9064
rect 18923 8996 19012 9024
rect 19153 9027 19211 9033
rect 18923 8993 18935 8996
rect 18877 8987 18935 8993
rect 19153 8993 19165 9027
rect 19199 8993 19211 9027
rect 19153 8987 19211 8993
rect 19429 9027 19487 9033
rect 19429 8993 19441 9027
rect 19475 9024 19487 9027
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19475 8996 19625 9024
rect 19475 8993 19487 8996
rect 19429 8987 19487 8993
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 8993 19763 9027
rect 19705 8987 19763 8993
rect 18414 8916 18420 8968
rect 18472 8956 18478 8968
rect 19444 8956 19472 8987
rect 19978 8984 19984 9036
rect 20036 9024 20042 9036
rect 20073 9027 20131 9033
rect 20073 9024 20085 9027
rect 20036 8996 20085 9024
rect 20036 8984 20042 8996
rect 20073 8993 20085 8996
rect 20119 8993 20131 9027
rect 20073 8987 20131 8993
rect 20533 9027 20591 9033
rect 20533 8993 20545 9027
rect 20579 9024 20591 9027
rect 20714 9024 20720 9036
rect 20579 8996 20720 9024
rect 20579 8993 20591 8996
rect 20533 8987 20591 8993
rect 20714 8984 20720 8996
rect 20772 8984 20778 9036
rect 20809 9027 20867 9033
rect 20809 8993 20821 9027
rect 20855 8993 20867 9027
rect 20809 8987 20867 8993
rect 20824 8956 20852 8987
rect 18472 8928 19472 8956
rect 20548 8928 20852 8956
rect 18472 8916 18478 8928
rect 19426 8888 19432 8900
rect 17888 8860 19432 8888
rect 19426 8848 19432 8860
rect 19484 8888 19490 8900
rect 20441 8891 20499 8897
rect 20441 8888 20453 8891
rect 19484 8860 20453 8888
rect 19484 8848 19490 8860
rect 20441 8857 20453 8860
rect 20487 8857 20499 8891
rect 20441 8851 20499 8857
rect 20548 8832 20576 8928
rect 20898 8916 20904 8968
rect 20956 8956 20962 8968
rect 21266 8956 21272 8968
rect 20956 8928 21272 8956
rect 20956 8916 20962 8928
rect 21266 8916 21272 8928
rect 21324 8956 21330 8968
rect 21453 8959 21511 8965
rect 21453 8956 21465 8959
rect 21324 8928 21465 8956
rect 21324 8916 21330 8928
rect 21453 8925 21465 8928
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 21729 8959 21787 8965
rect 21729 8956 21741 8959
rect 21692 8928 21741 8956
rect 21692 8916 21698 8928
rect 21729 8925 21741 8928
rect 21775 8925 21787 8959
rect 21729 8919 21787 8925
rect 14642 8820 14648 8832
rect 14476 8792 14648 8820
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 15841 8823 15899 8829
rect 15841 8820 15853 8823
rect 15528 8792 15853 8820
rect 15528 8780 15534 8792
rect 15841 8789 15853 8792
rect 15887 8789 15899 8823
rect 15841 8783 15899 8789
rect 17589 8823 17647 8829
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 18690 8820 18696 8832
rect 17635 8792 18696 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 20070 8820 20076 8832
rect 18840 8792 20076 8820
rect 18840 8780 18846 8792
rect 20070 8780 20076 8792
rect 20128 8820 20134 8832
rect 20165 8823 20223 8829
rect 20165 8820 20177 8823
rect 20128 8792 20177 8820
rect 20128 8780 20134 8792
rect 20165 8789 20177 8792
rect 20211 8789 20223 8823
rect 20165 8783 20223 8789
rect 20530 8780 20536 8832
rect 20588 8780 20594 8832
rect 23017 8823 23075 8829
rect 23017 8789 23029 8823
rect 23063 8820 23075 8823
rect 28442 8820 28448 8832
rect 23063 8792 28448 8820
rect 23063 8789 23075 8792
rect 23017 8783 23075 8789
rect 28442 8780 28448 8792
rect 28500 8780 28506 8832
rect 552 8730 31372 8752
rect 552 8678 4250 8730
rect 4302 8678 4314 8730
rect 4366 8678 4378 8730
rect 4430 8678 4442 8730
rect 4494 8678 4506 8730
rect 4558 8678 11955 8730
rect 12007 8678 12019 8730
rect 12071 8678 12083 8730
rect 12135 8678 12147 8730
rect 12199 8678 12211 8730
rect 12263 8678 19660 8730
rect 19712 8678 19724 8730
rect 19776 8678 19788 8730
rect 19840 8678 19852 8730
rect 19904 8678 19916 8730
rect 19968 8678 27365 8730
rect 27417 8678 27429 8730
rect 27481 8678 27493 8730
rect 27545 8678 27557 8730
rect 27609 8678 27621 8730
rect 27673 8678 31372 8730
rect 552 8656 31372 8678
rect 8662 8576 8668 8628
rect 8720 8576 8726 8628
rect 8941 8619 8999 8625
rect 8941 8585 8953 8619
rect 8987 8616 8999 8619
rect 9214 8616 9220 8628
rect 8987 8588 9220 8616
rect 8987 8585 8999 8588
rect 8941 8579 8999 8585
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 19334 8576 19340 8628
rect 19392 8576 19398 8628
rect 19794 8576 19800 8628
rect 19852 8616 19858 8628
rect 19852 8588 20852 8616
rect 19852 8576 19858 8588
rect 13633 8551 13691 8557
rect 13633 8517 13645 8551
rect 13679 8548 13691 8551
rect 14274 8548 14280 8560
rect 13679 8520 14280 8548
rect 13679 8517 13691 8520
rect 13633 8511 13691 8517
rect 14274 8508 14280 8520
rect 14332 8508 14338 8560
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 7944 8452 8125 8480
rect 7944 8421 7972 8452
rect 8113 8449 8125 8452
rect 8159 8480 8171 8483
rect 12805 8483 12863 8489
rect 8159 8452 9076 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8381 7987 8415
rect 7929 8375 7987 8381
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8478 8412 8484 8424
rect 8251 8384 8484 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8478 8372 8484 8384
rect 8536 8412 8542 8424
rect 9048 8421 9076 8452
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 12986 8480 12992 8492
rect 12851 8452 12992 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 12986 8440 12992 8452
rect 13044 8480 13050 8492
rect 19352 8480 19380 8576
rect 19786 8483 19844 8489
rect 19786 8480 19798 8483
rect 13044 8452 14688 8480
rect 19352 8452 19798 8480
rect 13044 8440 13050 8452
rect 14660 8424 14688 8452
rect 19786 8449 19798 8452
rect 19832 8449 19844 8483
rect 20824 8480 20852 8588
rect 21266 8576 21272 8628
rect 21324 8616 21330 8628
rect 21818 8616 21824 8628
rect 21324 8588 21824 8616
rect 21324 8576 21330 8588
rect 21818 8576 21824 8588
rect 21876 8616 21882 8628
rect 22649 8619 22707 8625
rect 22649 8616 22661 8619
rect 21876 8588 22661 8616
rect 21876 8576 21882 8588
rect 22649 8585 22661 8588
rect 22695 8585 22707 8619
rect 22649 8579 22707 8585
rect 21177 8551 21235 8557
rect 21177 8517 21189 8551
rect 21223 8548 21235 8551
rect 28258 8548 28264 8560
rect 21223 8520 28264 8548
rect 21223 8517 21235 8520
rect 21177 8511 21235 8517
rect 28258 8508 28264 8520
rect 28316 8508 28322 8560
rect 20824 8452 21404 8480
rect 19786 8443 19844 8449
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 8536 8384 8769 8412
rect 8536 8372 8542 8384
rect 8757 8381 8769 8384
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 9490 8412 9496 8424
rect 9079 8384 9496 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 7837 8347 7895 8353
rect 7837 8313 7849 8347
rect 7883 8344 7895 8347
rect 8386 8344 8392 8356
rect 7883 8316 8392 8344
rect 7883 8313 7895 8316
rect 7837 8307 7895 8313
rect 8386 8304 8392 8316
rect 8444 8344 8450 8356
rect 8772 8344 8800 8375
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 9732 8384 10701 8412
rect 9732 8372 9738 8384
rect 10689 8381 10701 8384
rect 10735 8412 10747 8415
rect 10778 8412 10784 8424
rect 10735 8384 10784 8412
rect 10735 8381 10747 8384
rect 10689 8375 10747 8381
rect 10778 8372 10784 8384
rect 10836 8372 10842 8424
rect 12549 8415 12607 8421
rect 12549 8381 12561 8415
rect 12595 8412 12607 8415
rect 13170 8412 13176 8424
rect 12595 8384 13176 8412
rect 12595 8381 12607 8384
rect 12549 8375 12607 8381
rect 13170 8372 13176 8384
rect 13228 8412 13234 8424
rect 13541 8415 13599 8421
rect 13541 8412 13553 8415
rect 13228 8384 13553 8412
rect 13228 8372 13234 8384
rect 13541 8381 13553 8384
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 13998 8372 14004 8424
rect 14056 8372 14062 8424
rect 14274 8372 14280 8424
rect 14332 8412 14338 8424
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 14332 8384 14381 8412
rect 14332 8372 14338 8384
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 14369 8375 14427 8381
rect 14642 8372 14648 8424
rect 14700 8372 14706 8424
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8412 19487 8415
rect 19610 8412 19616 8424
rect 19475 8384 19616 8412
rect 19475 8381 19487 8384
rect 19429 8375 19487 8381
rect 19610 8372 19616 8384
rect 19668 8372 19674 8424
rect 21376 8421 21404 8452
rect 19705 8415 19763 8421
rect 19705 8381 19717 8415
rect 19751 8412 19763 8415
rect 21361 8415 21419 8421
rect 19751 8384 20024 8412
rect 19751 8381 19763 8384
rect 19705 8375 19763 8381
rect 10422 8347 10480 8353
rect 10422 8344 10434 8347
rect 8444 8316 8708 8344
rect 8772 8316 10434 8344
rect 8444 8304 8450 8316
rect 8680 8288 8708 8316
rect 10422 8313 10434 8316
rect 10468 8313 10480 8347
rect 10422 8307 10480 8313
rect 13906 8304 13912 8356
rect 13964 8344 13970 8356
rect 14185 8347 14243 8353
rect 14185 8344 14197 8347
rect 13964 8316 14197 8344
rect 13964 8304 13970 8316
rect 14185 8313 14197 8316
rect 14231 8344 14243 8347
rect 14890 8347 14948 8353
rect 14890 8344 14902 8347
rect 14231 8316 14902 8344
rect 14231 8313 14243 8316
rect 14185 8307 14243 8313
rect 14890 8313 14902 8316
rect 14936 8313 14948 8347
rect 14890 8307 14948 8313
rect 17586 8304 17592 8356
rect 17644 8344 17650 8356
rect 19794 8344 19800 8356
rect 17644 8316 19800 8344
rect 17644 8304 17650 8316
rect 19794 8304 19800 8316
rect 19852 8304 19858 8356
rect 8662 8236 8668 8288
rect 8720 8236 8726 8288
rect 9306 8236 9312 8288
rect 9364 8236 9370 8288
rect 11422 8236 11428 8288
rect 11480 8236 11486 8288
rect 13262 8236 13268 8288
rect 13320 8236 13326 8288
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 14461 8279 14519 8285
rect 14461 8276 14473 8279
rect 13504 8248 14473 8276
rect 13504 8236 13510 8248
rect 14461 8245 14473 8248
rect 14507 8276 14519 8279
rect 14734 8276 14740 8288
rect 14507 8248 14740 8276
rect 14507 8245 14519 8248
rect 14461 8239 14519 8245
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 16025 8279 16083 8285
rect 16025 8245 16037 8279
rect 16071 8276 16083 8279
rect 16298 8276 16304 8288
rect 16071 8248 16304 8276
rect 16071 8245 16083 8248
rect 16025 8239 16083 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 19337 8279 19395 8285
rect 19337 8245 19349 8279
rect 19383 8276 19395 8279
rect 19426 8276 19432 8288
rect 19383 8248 19432 8276
rect 19383 8245 19395 8248
rect 19337 8239 19395 8245
rect 19426 8236 19432 8248
rect 19484 8236 19490 8288
rect 19613 8279 19671 8285
rect 19613 8245 19625 8279
rect 19659 8276 19671 8279
rect 19886 8276 19892 8288
rect 19659 8248 19892 8276
rect 19659 8245 19671 8248
rect 19613 8239 19671 8245
rect 19886 8236 19892 8248
rect 19944 8236 19950 8288
rect 19996 8276 20024 8384
rect 21361 8381 21373 8415
rect 21407 8412 21419 8415
rect 21542 8412 21548 8424
rect 21407 8384 21548 8412
rect 21407 8381 21419 8384
rect 21361 8375 21419 8381
rect 21542 8372 21548 8384
rect 21600 8372 21606 8424
rect 23198 8372 23204 8424
rect 23256 8372 23262 8424
rect 20070 8353 20076 8356
rect 20064 8307 20076 8353
rect 20128 8344 20134 8356
rect 20128 8316 20164 8344
rect 20070 8304 20076 8307
rect 20128 8304 20134 8316
rect 20990 8276 20996 8288
rect 19996 8248 20996 8276
rect 20990 8236 20996 8248
rect 21048 8236 21054 8288
rect 23290 8236 23296 8288
rect 23348 8236 23354 8288
rect 552 8186 31531 8208
rect 552 8134 8102 8186
rect 8154 8134 8166 8186
rect 8218 8134 8230 8186
rect 8282 8134 8294 8186
rect 8346 8134 8358 8186
rect 8410 8134 15807 8186
rect 15859 8134 15871 8186
rect 15923 8134 15935 8186
rect 15987 8134 15999 8186
rect 16051 8134 16063 8186
rect 16115 8134 23512 8186
rect 23564 8134 23576 8186
rect 23628 8134 23640 8186
rect 23692 8134 23704 8186
rect 23756 8134 23768 8186
rect 23820 8134 31217 8186
rect 31269 8134 31281 8186
rect 31333 8134 31345 8186
rect 31397 8134 31409 8186
rect 31461 8134 31473 8186
rect 31525 8134 31531 8186
rect 552 8112 31531 8134
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8478 8072 8484 8084
rect 8343 8044 8484 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 13320 8044 13461 8072
rect 13320 8032 13326 8044
rect 13449 8041 13461 8044
rect 13495 8072 13507 8075
rect 13814 8072 13820 8084
rect 13495 8044 13820 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 17586 8072 17592 8084
rect 15948 8044 17592 8072
rect 9214 8004 9220 8016
rect 7769 7976 9220 8004
rect 7769 7948 7797 7976
rect 9214 7964 9220 7976
rect 9272 7964 9278 8016
rect 9858 7964 9864 8016
rect 9916 8004 9922 8016
rect 15948 8013 15976 8044
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 19426 8032 19432 8084
rect 19484 8032 19490 8084
rect 19610 8032 19616 8084
rect 19668 8032 19674 8084
rect 19886 8032 19892 8084
rect 19944 8032 19950 8084
rect 20714 8032 20720 8084
rect 20772 8032 20778 8084
rect 20990 8032 20996 8084
rect 21048 8032 21054 8084
rect 10781 8007 10839 8013
rect 10781 8004 10793 8007
rect 9916 7976 10793 8004
rect 9916 7964 9922 7976
rect 10781 7973 10793 7976
rect 10827 8004 10839 8007
rect 15933 8007 15991 8013
rect 15933 8004 15945 8007
rect 10827 7976 15945 8004
rect 10827 7973 10839 7976
rect 10781 7967 10839 7973
rect 15933 7973 15945 7976
rect 15979 7973 15991 8007
rect 16206 8004 16212 8016
rect 15933 7967 15991 7973
rect 16132 7976 16212 8004
rect 7742 7896 7748 7948
rect 7800 7945 7806 7948
rect 7800 7899 7812 7945
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 8570 7936 8576 7948
rect 8435 7908 8576 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 7800 7896 7806 7899
rect 8018 7828 8024 7880
rect 8076 7828 8082 7880
rect 8496 7868 8524 7908
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 8665 7939 8723 7945
rect 8665 7905 8677 7939
rect 8711 7936 8723 7939
rect 8754 7936 8760 7948
rect 8711 7908 8760 7936
rect 8711 7905 8723 7908
rect 8665 7899 8723 7905
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 8941 7939 8999 7945
rect 8941 7905 8953 7939
rect 8987 7936 8999 7939
rect 10318 7936 10324 7948
rect 8987 7908 10324 7936
rect 8987 7905 8999 7908
rect 8941 7899 8999 7905
rect 10318 7896 10324 7908
rect 10376 7936 10382 7948
rect 12170 7939 12228 7945
rect 12170 7936 12182 7939
rect 10376 7908 12182 7936
rect 10376 7896 10382 7908
rect 12170 7905 12182 7908
rect 12216 7905 12228 7939
rect 12170 7899 12228 7905
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 13035 7908 13093 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13081 7905 13093 7908
rect 13127 7936 13139 7939
rect 13446 7936 13452 7948
rect 13127 7908 13452 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 13817 7939 13875 7945
rect 13817 7936 13829 7939
rect 13587 7908 13829 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 13817 7905 13829 7908
rect 13863 7936 13875 7939
rect 13906 7936 13912 7948
rect 13863 7908 13912 7936
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 13906 7896 13912 7908
rect 13964 7896 13970 7948
rect 13998 7896 14004 7948
rect 14056 7936 14062 7948
rect 16132 7945 16160 7976
rect 16206 7964 16212 7976
rect 16264 8004 16270 8016
rect 18040 8007 18098 8013
rect 16264 7976 17172 8004
rect 16264 7964 16270 7976
rect 14093 7939 14151 7945
rect 14093 7936 14105 7939
rect 14056 7908 14105 7936
rect 14056 7896 14062 7908
rect 14093 7905 14105 7908
rect 14139 7905 14151 7939
rect 14093 7899 14151 7905
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7905 16175 7939
rect 16373 7939 16431 7945
rect 16373 7936 16385 7939
rect 16117 7899 16175 7905
rect 16224 7908 16385 7936
rect 8849 7871 8907 7877
rect 8849 7868 8861 7871
rect 8496 7840 8861 7868
rect 8849 7837 8861 7840
rect 8895 7837 8907 7871
rect 8849 7831 8907 7837
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 12483 7840 14688 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 6638 7692 6644 7744
rect 6696 7692 6702 7744
rect 8036 7732 8064 7828
rect 8478 7760 8484 7812
rect 8536 7800 8542 7812
rect 8573 7803 8631 7809
rect 8573 7800 8585 7803
rect 8536 7772 8585 7800
rect 8536 7760 8542 7772
rect 8573 7769 8585 7772
rect 8619 7769 8631 7803
rect 8573 7763 8631 7769
rect 13173 7803 13231 7809
rect 13173 7769 13185 7803
rect 13219 7800 13231 7803
rect 13722 7800 13728 7812
rect 13219 7772 13728 7800
rect 13219 7769 13231 7772
rect 13173 7763 13231 7769
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 14660 7744 14688 7840
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 16224 7868 16252 7908
rect 16373 7905 16385 7908
rect 16419 7905 16431 7939
rect 16373 7899 16431 7905
rect 14792 7840 16252 7868
rect 14792 7828 14798 7840
rect 17144 7800 17172 7976
rect 18040 7973 18052 8007
rect 18086 8004 18098 8007
rect 19444 8004 19472 8032
rect 18086 7976 19472 8004
rect 19628 8004 19656 8032
rect 20162 8004 20168 8016
rect 19628 7976 20168 8004
rect 18086 7973 18098 7976
rect 18040 7967 18098 7973
rect 19444 7936 19472 7976
rect 20162 7964 20168 7976
rect 20220 8004 20226 8016
rect 20438 8004 20444 8016
rect 20220 7976 20444 8004
rect 20220 7964 20226 7976
rect 20438 7964 20444 7976
rect 20496 7964 20502 8016
rect 19981 7939 20039 7945
rect 19981 7936 19993 7939
rect 19444 7908 19993 7936
rect 19981 7905 19993 7908
rect 20027 7905 20039 7939
rect 19981 7899 20039 7905
rect 20254 7896 20260 7948
rect 20312 7896 20318 7948
rect 20349 7939 20407 7945
rect 20349 7905 20361 7939
rect 20395 7936 20407 7939
rect 20530 7936 20536 7948
rect 20395 7908 20536 7936
rect 20395 7905 20407 7908
rect 20349 7899 20407 7905
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7837 17831 7871
rect 17773 7831 17831 7837
rect 17788 7800 17816 7831
rect 17052 7772 17816 7800
rect 20165 7803 20223 7809
rect 17052 7744 17080 7772
rect 20165 7769 20177 7803
rect 20211 7800 20223 7803
rect 20364 7800 20392 7899
rect 20530 7896 20536 7908
rect 20588 7896 20594 7948
rect 20732 7936 20760 8032
rect 21008 8004 21036 8032
rect 21361 8007 21419 8013
rect 21361 8004 21373 8007
rect 21008 7976 21373 8004
rect 21100 7945 21128 7976
rect 21361 7973 21373 7976
rect 21407 8004 21419 8007
rect 21634 8004 21640 8016
rect 21407 7976 21640 8004
rect 21407 7973 21419 7976
rect 21361 7967 21419 7973
rect 21634 7964 21640 7976
rect 21692 7964 21698 8016
rect 22278 8004 22284 8016
rect 21744 7976 22284 8004
rect 21744 7945 21772 7976
rect 22278 7964 22284 7976
rect 22336 8004 22342 8016
rect 23290 8004 23296 8016
rect 22336 7976 23296 8004
rect 22336 7964 22342 7976
rect 23290 7964 23296 7976
rect 23348 7964 23354 8016
rect 20809 7939 20867 7945
rect 20809 7936 20821 7939
rect 20732 7908 20821 7936
rect 20809 7905 20821 7908
rect 20855 7936 20867 7939
rect 20993 7939 21051 7945
rect 20993 7936 21005 7939
rect 20855 7908 21005 7936
rect 20855 7905 20867 7908
rect 20809 7899 20867 7905
rect 20993 7905 21005 7908
rect 21039 7905 21051 7939
rect 20993 7899 21051 7905
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7905 21143 7939
rect 21085 7899 21143 7905
rect 21269 7939 21327 7945
rect 21269 7905 21281 7939
rect 21315 7905 21327 7939
rect 21269 7899 21327 7905
rect 21729 7939 21787 7945
rect 21729 7905 21741 7939
rect 21775 7905 21787 7939
rect 21729 7899 21787 7905
rect 20211 7772 20392 7800
rect 20211 7769 20223 7772
rect 20165 7763 20223 7769
rect 20438 7760 20444 7812
rect 20496 7800 20502 7812
rect 21284 7800 21312 7899
rect 21818 7896 21824 7948
rect 21876 7936 21882 7948
rect 21913 7939 21971 7945
rect 21913 7936 21925 7939
rect 21876 7908 21925 7936
rect 21876 7896 21882 7908
rect 21913 7905 21925 7908
rect 21959 7905 21971 7939
rect 22169 7939 22227 7945
rect 22169 7936 22181 7939
rect 21913 7899 21971 7905
rect 22020 7908 22181 7936
rect 21634 7828 21640 7880
rect 21692 7868 21698 7880
rect 22020 7868 22048 7908
rect 22169 7905 22181 7908
rect 22215 7905 22227 7939
rect 22169 7899 22227 7905
rect 21692 7840 22048 7868
rect 21692 7828 21698 7840
rect 20496 7772 21312 7800
rect 20496 7760 20502 7772
rect 9493 7735 9551 7741
rect 9493 7732 9505 7735
rect 8036 7704 9505 7732
rect 9493 7701 9505 7704
rect 9539 7732 9551 7735
rect 9674 7732 9680 7744
rect 9539 7704 9680 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 11020 7704 11069 7732
rect 11020 7692 11026 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 12894 7692 12900 7744
rect 12952 7692 12958 7744
rect 14001 7735 14059 7741
rect 14001 7701 14013 7735
rect 14047 7732 14059 7735
rect 14090 7732 14096 7744
rect 14047 7704 14096 7732
rect 14047 7701 14059 7704
rect 14001 7695 14059 7701
rect 14090 7692 14096 7704
rect 14148 7692 14154 7744
rect 14642 7692 14648 7744
rect 14700 7692 14706 7744
rect 17034 7692 17040 7744
rect 17092 7692 17098 7744
rect 17494 7692 17500 7744
rect 17552 7692 17558 7744
rect 19153 7735 19211 7741
rect 19153 7701 19165 7735
rect 19199 7732 19211 7735
rect 19978 7732 19984 7744
rect 19199 7704 19984 7732
rect 19199 7701 19211 7704
rect 19153 7695 19211 7701
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 20070 7692 20076 7744
rect 20128 7732 20134 7744
rect 20717 7735 20775 7741
rect 20717 7732 20729 7735
rect 20128 7704 20729 7732
rect 20128 7692 20134 7704
rect 20717 7701 20729 7704
rect 20763 7701 20775 7735
rect 20717 7695 20775 7701
rect 23293 7735 23351 7741
rect 23293 7701 23305 7735
rect 23339 7732 23351 7735
rect 28258 7732 28264 7744
rect 23339 7704 28264 7732
rect 23339 7701 23351 7704
rect 23293 7695 23351 7701
rect 28258 7692 28264 7704
rect 28316 7692 28322 7744
rect 552 7642 31372 7664
rect 552 7590 4250 7642
rect 4302 7590 4314 7642
rect 4366 7590 4378 7642
rect 4430 7590 4442 7642
rect 4494 7590 4506 7642
rect 4558 7590 11955 7642
rect 12007 7590 12019 7642
rect 12071 7590 12083 7642
rect 12135 7590 12147 7642
rect 12199 7590 12211 7642
rect 12263 7590 19660 7642
rect 19712 7590 19724 7642
rect 19776 7590 19788 7642
rect 19840 7590 19852 7642
rect 19904 7590 19916 7642
rect 19968 7590 27365 7642
rect 27417 7590 27429 7642
rect 27481 7590 27493 7642
rect 27545 7590 27557 7642
rect 27609 7590 27621 7642
rect 27673 7590 31372 7642
rect 552 7568 31372 7590
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7800 7500 7849 7528
rect 7800 7488 7806 7500
rect 7837 7497 7849 7500
rect 7883 7497 7895 7531
rect 7837 7491 7895 7497
rect 9125 7531 9183 7537
rect 9125 7497 9137 7531
rect 9171 7528 9183 7531
rect 10318 7528 10324 7540
rect 9171 7500 10324 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 7561 7463 7619 7469
rect 7561 7429 7573 7463
rect 7607 7460 7619 7463
rect 8754 7460 8760 7472
rect 7607 7432 8760 7460
rect 7607 7429 7619 7432
rect 7561 7423 7619 7429
rect 8754 7420 8760 7432
rect 8812 7460 8818 7472
rect 8849 7463 8907 7469
rect 8849 7460 8861 7463
rect 8812 7432 8861 7460
rect 8812 7420 8818 7432
rect 8849 7429 8861 7432
rect 8895 7429 8907 7463
rect 9140 7460 9168 7491
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 12713 7531 12771 7537
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 12894 7528 12900 7540
rect 12759 7500 12900 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 14369 7531 14427 7537
rect 14369 7497 14381 7531
rect 14415 7528 14427 7531
rect 14734 7528 14740 7540
rect 14415 7500 14740 7528
rect 14415 7497 14427 7500
rect 14369 7491 14427 7497
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 20162 7488 20168 7540
rect 20220 7528 20226 7540
rect 20257 7531 20315 7537
rect 20257 7528 20269 7531
rect 20220 7500 20269 7528
rect 20220 7488 20226 7500
rect 20257 7497 20269 7500
rect 20303 7497 20315 7531
rect 20257 7491 20315 7497
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 21634 7528 21640 7540
rect 20588 7500 21640 7528
rect 20588 7488 20594 7500
rect 21634 7488 21640 7500
rect 21692 7488 21698 7540
rect 22278 7528 22284 7540
rect 21744 7500 22284 7528
rect 8849 7423 8907 7429
rect 8956 7432 9168 7460
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 8956 7392 8984 7432
rect 9214 7420 9220 7472
rect 9272 7460 9278 7472
rect 11885 7463 11943 7469
rect 9272 7432 9674 7460
rect 9272 7420 9278 7432
rect 7800 7364 8064 7392
rect 7800 7352 7806 7364
rect 7650 7284 7656 7336
rect 7708 7284 7714 7336
rect 7926 7284 7932 7336
rect 7984 7284 7990 7336
rect 8036 7333 8064 7364
rect 8772 7364 8984 7392
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8570 7326 8576 7336
rect 8496 7324 8576 7326
rect 8159 7298 8576 7324
rect 8159 7296 8524 7298
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8570 7284 8576 7298
rect 8628 7284 8634 7336
rect 8772 7324 8800 7364
rect 9490 7352 9496 7404
rect 9548 7352 9554 7404
rect 9646 7392 9674 7432
rect 11885 7429 11897 7463
rect 11931 7460 11943 7463
rect 11974 7460 11980 7472
rect 11931 7432 11980 7460
rect 11931 7429 11943 7432
rect 11885 7423 11943 7429
rect 11974 7420 11980 7432
rect 12032 7460 12038 7472
rect 12526 7460 12532 7472
rect 12032 7432 12532 7460
rect 12032 7420 12038 7432
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 19981 7463 20039 7469
rect 12636 7432 13860 7460
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 9600 7364 10057 7392
rect 8933 7329 8991 7335
rect 8933 7326 8945 7329
rect 8864 7324 8945 7326
rect 8772 7298 8945 7324
rect 8772 7296 8892 7298
rect 8933 7295 8945 7298
rect 8979 7295 8991 7329
rect 8933 7289 8991 7295
rect 9033 7327 9091 7333
rect 9033 7293 9045 7327
rect 9079 7326 9091 7327
rect 9079 7324 9168 7326
rect 9398 7324 9404 7336
rect 9079 7298 9404 7324
rect 9079 7293 9091 7298
rect 9140 7296 9404 7298
rect 9033 7287 9091 7293
rect 9398 7284 9404 7296
rect 9456 7324 9462 7336
rect 9600 7333 9628 7364
rect 10045 7361 10057 7364
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 12636 7343 12664 7432
rect 13722 7352 13728 7404
rect 13780 7352 13786 7404
rect 13832 7401 13860 7432
rect 19981 7429 19993 7463
rect 20027 7460 20039 7463
rect 20622 7460 20628 7472
rect 20027 7432 20628 7460
rect 20027 7429 20039 7432
rect 19981 7423 20039 7429
rect 20622 7420 20628 7432
rect 20680 7460 20686 7472
rect 20680 7432 21220 7460
rect 20680 7420 20686 7432
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7392 13875 7395
rect 14090 7392 14096 7404
rect 13863 7364 14096 7392
rect 13863 7361 13875 7364
rect 13817 7355 13875 7361
rect 14090 7352 14096 7364
rect 14148 7392 14154 7404
rect 19426 7392 19432 7404
rect 14148 7364 14412 7392
rect 14148 7352 14154 7364
rect 12621 7337 12679 7343
rect 9585 7327 9643 7333
rect 9456 7296 9536 7324
rect 9456 7284 9462 7296
rect 8481 7259 8539 7265
rect 8481 7225 8493 7259
rect 8527 7256 8539 7259
rect 8662 7256 8668 7268
rect 8527 7228 8668 7256
rect 8527 7225 8539 7228
rect 8481 7219 8539 7225
rect 8662 7216 8668 7228
rect 8720 7216 8726 7268
rect 9508 7256 9536 7296
rect 9585 7293 9597 7327
rect 9631 7293 9643 7327
rect 9585 7287 9643 7293
rect 9858 7284 9864 7336
rect 9916 7284 9922 7336
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 9769 7259 9827 7265
rect 9769 7256 9781 7259
rect 9508 7228 9781 7256
rect 9769 7225 9781 7228
rect 9815 7225 9827 7259
rect 9769 7219 9827 7225
rect 8754 7148 8760 7200
rect 8812 7188 8818 7200
rect 9968 7188 9996 7287
rect 10410 7284 10416 7336
rect 10468 7284 10474 7336
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 12023 7296 12173 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12161 7293 12173 7296
rect 12207 7293 12219 7327
rect 12161 7287 12219 7293
rect 8812 7160 9996 7188
rect 12176 7188 12204 7287
rect 12250 7284 12256 7336
rect 12308 7284 12314 7336
rect 12529 7327 12587 7333
rect 12529 7293 12541 7327
rect 12575 7324 12587 7327
rect 12621 7324 12633 7337
rect 12575 7303 12633 7324
rect 12667 7303 12679 7337
rect 12575 7297 12679 7303
rect 12575 7296 12664 7297
rect 12575 7293 12587 7296
rect 12529 7287 12587 7293
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 13081 7327 13139 7333
rect 13081 7324 13093 7327
rect 12952 7296 13093 7324
rect 12952 7284 12958 7296
rect 13081 7293 13093 7296
rect 13127 7324 13139 7327
rect 13173 7327 13231 7333
rect 13173 7324 13185 7327
rect 13127 7296 13185 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 13173 7293 13185 7296
rect 13219 7293 13231 7327
rect 13740 7324 13768 7352
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 13740 7296 13921 7324
rect 13173 7287 13231 7293
rect 13909 7293 13921 7296
rect 13955 7324 13967 7327
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 13955 7296 14013 7324
rect 13955 7293 13967 7296
rect 13909 7287 13967 7293
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 14182 7284 14188 7336
rect 14240 7324 14246 7336
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 14240 7296 14289 7324
rect 14240 7284 14246 7296
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 14384 7324 14412 7364
rect 19352 7364 19432 7392
rect 15758 7327 15816 7333
rect 15758 7324 15770 7327
rect 14384 7296 15770 7324
rect 14277 7287 14335 7293
rect 15758 7293 15770 7296
rect 15804 7293 15816 7327
rect 15758 7287 15816 7293
rect 16025 7327 16083 7333
rect 16025 7293 16037 7327
rect 16071 7324 16083 7327
rect 16071 7296 17080 7324
rect 16071 7293 16083 7296
rect 16025 7287 16083 7293
rect 12989 7259 13047 7265
rect 12989 7225 13001 7259
rect 13035 7256 13047 7259
rect 13035 7228 14136 7256
rect 13035 7225 13047 7228
rect 12989 7219 13047 7225
rect 14108 7200 14136 7228
rect 17052 7200 17080 7296
rect 17586 7284 17592 7336
rect 17644 7324 17650 7336
rect 19352 7333 19380 7364
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 20364 7364 20576 7392
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 17644 7296 18521 7324
rect 17644 7284 17650 7296
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 19337 7327 19395 7333
rect 19337 7293 19349 7327
rect 19383 7293 19395 7327
rect 19337 7287 19395 7293
rect 19794 7284 19800 7336
rect 19852 7284 19858 7336
rect 20364 7333 20392 7364
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7293 19947 7327
rect 19889 7287 19947 7293
rect 20349 7327 20407 7333
rect 20349 7293 20361 7327
rect 20395 7293 20407 7327
rect 20349 7287 20407 7293
rect 20441 7327 20499 7333
rect 20441 7293 20453 7327
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 19429 7259 19487 7265
rect 19429 7225 19441 7259
rect 19475 7256 19487 7259
rect 19705 7259 19763 7265
rect 19705 7256 19717 7259
rect 19475 7228 19717 7256
rect 19475 7225 19487 7228
rect 19429 7219 19487 7225
rect 19705 7225 19717 7228
rect 19751 7256 19763 7259
rect 19904 7256 19932 7287
rect 20456 7256 20484 7287
rect 20548 7265 20576 7364
rect 20714 7284 20720 7336
rect 20772 7333 20778 7336
rect 21192 7333 21220 7432
rect 21744 7333 21772 7500
rect 22278 7488 22284 7500
rect 22336 7488 22342 7540
rect 21818 7420 21824 7472
rect 21876 7460 21882 7472
rect 21876 7432 22048 7460
rect 21876 7420 21882 7432
rect 22020 7401 22048 7432
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 20772 7324 20783 7333
rect 21177 7327 21235 7333
rect 20772 7296 20817 7324
rect 20772 7287 20783 7296
rect 21177 7293 21189 7327
rect 21223 7324 21235 7327
rect 21269 7327 21327 7333
rect 21269 7324 21281 7327
rect 21223 7296 21281 7324
rect 21223 7293 21235 7296
rect 21177 7287 21235 7293
rect 21269 7293 21281 7296
rect 21315 7293 21327 7327
rect 21269 7287 21327 7293
rect 21361 7327 21419 7333
rect 21361 7293 21373 7327
rect 21407 7324 21419 7327
rect 21729 7327 21787 7333
rect 21729 7324 21741 7327
rect 21407 7296 21741 7324
rect 21407 7293 21419 7296
rect 21361 7287 21419 7293
rect 21729 7293 21741 7296
rect 21775 7293 21787 7327
rect 21729 7287 21787 7293
rect 20772 7284 20778 7287
rect 23198 7284 23204 7336
rect 23256 7284 23262 7336
rect 19751 7228 20484 7256
rect 20533 7259 20591 7265
rect 19751 7225 19763 7228
rect 19705 7219 19763 7225
rect 20533 7225 20545 7259
rect 20579 7256 20591 7259
rect 20809 7259 20867 7265
rect 20809 7256 20821 7259
rect 20579 7228 20821 7256
rect 20579 7225 20591 7228
rect 20533 7219 20591 7225
rect 20809 7225 20821 7228
rect 20855 7256 20867 7259
rect 22272 7259 22330 7265
rect 22272 7256 22284 7259
rect 20855 7228 22284 7256
rect 20855 7225 20867 7228
rect 20809 7219 20867 7225
rect 22272 7225 22284 7228
rect 22318 7256 22330 7259
rect 23216 7256 23244 7284
rect 22318 7228 23244 7256
rect 22318 7225 22330 7228
rect 22272 7219 22330 7225
rect 12342 7188 12348 7200
rect 12176 7160 12348 7188
rect 8812 7148 8818 7160
rect 12342 7148 12348 7160
rect 12400 7188 12406 7200
rect 12437 7191 12495 7197
rect 12437 7188 12449 7191
rect 12400 7160 12449 7188
rect 12400 7148 12406 7160
rect 12437 7157 12449 7160
rect 12483 7157 12495 7191
rect 12437 7151 12495 7157
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 12584 7160 13277 7188
rect 12584 7148 12590 7160
rect 13265 7157 13277 7160
rect 13311 7157 13323 7191
rect 13265 7151 13323 7157
rect 14090 7148 14096 7200
rect 14148 7148 14154 7200
rect 14458 7148 14464 7200
rect 14516 7188 14522 7200
rect 14645 7191 14703 7197
rect 14645 7188 14657 7191
rect 14516 7160 14657 7188
rect 14516 7148 14522 7160
rect 14645 7157 14657 7160
rect 14691 7157 14703 7191
rect 14645 7151 14703 7157
rect 17034 7148 17040 7200
rect 17092 7148 17098 7200
rect 20254 7148 20260 7200
rect 20312 7188 20318 7200
rect 20714 7188 20720 7200
rect 20312 7160 20720 7188
rect 20312 7148 20318 7160
rect 20714 7148 20720 7160
rect 20772 7188 20778 7200
rect 20898 7188 20904 7200
rect 20772 7160 20904 7188
rect 20772 7148 20778 7160
rect 20898 7148 20904 7160
rect 20956 7188 20962 7200
rect 21085 7191 21143 7197
rect 21085 7188 21097 7191
rect 20956 7160 21097 7188
rect 20956 7148 20962 7160
rect 21085 7157 21097 7160
rect 21131 7157 21143 7191
rect 21085 7151 21143 7157
rect 23385 7191 23443 7197
rect 23385 7157 23397 7191
rect 23431 7188 23443 7191
rect 28258 7188 28264 7200
rect 23431 7160 28264 7188
rect 23431 7157 23443 7160
rect 23385 7151 23443 7157
rect 28258 7148 28264 7160
rect 28316 7148 28322 7200
rect 552 7098 31531 7120
rect 552 7046 8102 7098
rect 8154 7046 8166 7098
rect 8218 7046 8230 7098
rect 8282 7046 8294 7098
rect 8346 7046 8358 7098
rect 8410 7046 15807 7098
rect 15859 7046 15871 7098
rect 15923 7046 15935 7098
rect 15987 7046 15999 7098
rect 16051 7046 16063 7098
rect 16115 7046 23512 7098
rect 23564 7046 23576 7098
rect 23628 7046 23640 7098
rect 23692 7046 23704 7098
rect 23756 7046 23768 7098
rect 23820 7046 31217 7098
rect 31269 7046 31281 7098
rect 31333 7046 31345 7098
rect 31397 7046 31409 7098
rect 31461 7046 31473 7098
rect 31525 7046 31531 7098
rect 552 7024 31531 7046
rect 7650 6944 7656 6996
rect 7708 6944 7714 6996
rect 7926 6944 7932 6996
rect 7984 6984 7990 6996
rect 9398 6984 9404 6996
rect 7984 6956 9404 6984
rect 7984 6944 7990 6956
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 9858 6944 9864 6996
rect 9916 6944 9922 6996
rect 10410 6944 10416 6996
rect 10468 6944 10474 6996
rect 12342 6944 12348 6996
rect 12400 6944 12406 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 14458 6984 14464 6996
rect 12952 6956 14464 6984
rect 12952 6944 12958 6956
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 19426 6984 19432 6996
rect 19260 6956 19432 6984
rect 7668 6916 7696 6944
rect 9876 6916 9904 6944
rect 10134 6916 10140 6928
rect 7668 6888 10140 6916
rect 8956 6857 8984 6888
rect 10134 6876 10140 6888
rect 10192 6876 10198 6928
rect 8950 6851 9008 6857
rect 8950 6817 8962 6851
rect 8996 6817 9008 6851
rect 8950 6811 9008 6817
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9769 6851 9827 6857
rect 9769 6848 9781 6851
rect 9539 6820 9781 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9769 6817 9781 6820
rect 9815 6817 9827 6851
rect 9769 6811 9827 6817
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9907 6820 10057 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 10045 6817 10057 6820
rect 10091 6848 10103 6851
rect 10428 6848 10456 6944
rect 11974 6916 11980 6928
rect 11164 6888 11980 6916
rect 11164 6857 11192 6888
rect 11974 6876 11980 6888
rect 12032 6876 12038 6928
rect 10091 6820 10456 6848
rect 10505 6851 10563 6857
rect 10091 6817 10103 6820
rect 10045 6811 10103 6817
rect 10505 6817 10517 6851
rect 10551 6848 10563 6851
rect 10781 6851 10839 6857
rect 10781 6848 10793 6851
rect 10551 6820 10793 6848
rect 10551 6817 10563 6820
rect 10505 6811 10563 6817
rect 10781 6817 10793 6820
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 11149 6851 11207 6857
rect 11149 6817 11161 6851
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6848 11483 6851
rect 11701 6851 11759 6857
rect 11701 6848 11713 6851
rect 11471 6820 11713 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 11701 6817 11713 6820
rect 11747 6848 11759 6851
rect 11747 6820 11928 6848
rect 11992 6847 12020 6876
rect 11747 6817 11759 6820
rect 11701 6811 11759 6817
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6780 9275 6783
rect 9674 6780 9680 6792
rect 9263 6752 9680 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 9784 6712 9812 6811
rect 10796 6780 10824 6811
rect 10796 6752 11652 6780
rect 9784 6684 10272 6712
rect 7834 6604 7840 6656
rect 7892 6604 7898 6656
rect 10244 6644 10272 6684
rect 10612 6684 11376 6712
rect 10612 6644 10640 6684
rect 11348 6656 11376 6684
rect 11624 6656 11652 6752
rect 11900 6721 11928 6820
rect 11977 6841 12035 6847
rect 11977 6807 11989 6841
rect 12023 6807 12035 6841
rect 12250 6808 12256 6860
rect 12308 6808 12314 6860
rect 12360 6857 12388 6944
rect 13900 6919 13958 6925
rect 13900 6885 13912 6919
rect 13946 6916 13958 6919
rect 14090 6916 14096 6928
rect 13946 6888 14096 6916
rect 13946 6885 13958 6888
rect 13900 6879 13958 6885
rect 12345 6851 12403 6857
rect 12345 6817 12357 6851
rect 12391 6817 12403 6851
rect 13915 6848 13943 6879
rect 14090 6876 14096 6888
rect 14148 6876 14154 6928
rect 19260 6925 19288 6956
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 19794 6944 19800 6996
rect 19852 6984 19858 6996
rect 20349 6987 20407 6993
rect 20349 6984 20361 6987
rect 19852 6956 20361 6984
rect 19852 6944 19858 6956
rect 20349 6953 20361 6956
rect 20395 6953 20407 6987
rect 20349 6947 20407 6953
rect 19245 6919 19303 6925
rect 19245 6916 19257 6919
rect 19076 6888 19257 6916
rect 12345 6811 12403 6817
rect 12452 6820 13943 6848
rect 11977 6801 12035 6807
rect 12268 6780 12296 6808
rect 12452 6780 12480 6820
rect 17034 6808 17040 6860
rect 17092 6808 17098 6860
rect 17304 6851 17362 6857
rect 17304 6817 17316 6851
rect 17350 6848 17362 6851
rect 17350 6820 18092 6848
rect 17350 6817 17362 6820
rect 17304 6811 17362 6817
rect 12268 6752 12480 6780
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6749 13691 6783
rect 13633 6743 13691 6749
rect 11885 6715 11943 6721
rect 11885 6681 11897 6715
rect 11931 6712 11943 6715
rect 12161 6715 12219 6721
rect 12161 6712 12173 6715
rect 11931 6684 12173 6712
rect 11931 6681 11943 6684
rect 11885 6675 11943 6681
rect 12161 6681 12173 6684
rect 12207 6681 12219 6715
rect 12161 6675 12219 6681
rect 10244 6616 10640 6644
rect 10686 6604 10692 6656
rect 10744 6644 10750 6656
rect 11057 6647 11115 6653
rect 11057 6644 11069 6647
rect 10744 6616 11069 6644
rect 10744 6604 10750 6616
rect 11057 6613 11069 6616
rect 11103 6613 11115 6647
rect 11057 6607 11115 6613
rect 11330 6604 11336 6656
rect 11388 6604 11394 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 11664 6616 12449 6644
rect 11664 6604 11670 6616
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 13648 6644 13676 6743
rect 14642 6644 14648 6656
rect 13648 6616 14648 6644
rect 12437 6607 12495 6613
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 15010 6604 15016 6656
rect 15068 6604 15074 6656
rect 17052 6644 17080 6808
rect 18064 6780 18092 6820
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 18601 6851 18659 6857
rect 18601 6848 18613 6851
rect 18196 6820 18613 6848
rect 18196 6808 18202 6820
rect 18601 6817 18613 6820
rect 18647 6817 18659 6851
rect 18601 6811 18659 6817
rect 18782 6808 18788 6860
rect 18840 6848 18846 6860
rect 18877 6851 18935 6857
rect 18877 6848 18889 6851
rect 18840 6820 18889 6848
rect 18840 6808 18846 6820
rect 18877 6817 18889 6820
rect 18923 6817 18935 6851
rect 19076 6848 19104 6888
rect 19245 6885 19257 6888
rect 19291 6885 19303 6919
rect 19245 6879 19303 6885
rect 19521 6919 19579 6925
rect 19521 6885 19533 6919
rect 19567 6916 19579 6919
rect 20070 6916 20076 6928
rect 19567 6888 19932 6916
rect 19567 6885 19579 6888
rect 19521 6879 19579 6885
rect 19329 6851 19387 6857
rect 19329 6848 19341 6851
rect 18877 6811 18935 6817
rect 18984 6820 19104 6848
rect 19168 6820 19341 6848
rect 18693 6783 18751 6789
rect 18693 6780 18705 6783
rect 18064 6752 18705 6780
rect 18693 6749 18705 6752
rect 18739 6780 18751 6783
rect 18984 6780 19012 6820
rect 18739 6752 19012 6780
rect 18739 6749 18751 6752
rect 18693 6743 18751 6749
rect 19058 6712 19064 6724
rect 18432 6684 19064 6712
rect 18322 6644 18328 6656
rect 17052 6616 18328 6644
rect 18322 6604 18328 6616
rect 18380 6604 18386 6656
rect 18432 6653 18460 6684
rect 19058 6672 19064 6684
rect 19116 6672 19122 6724
rect 19168 6656 19196 6820
rect 19306 6817 19341 6820
rect 19375 6817 19387 6851
rect 19306 6811 19387 6817
rect 19426 6814 19432 6866
rect 19484 6814 19490 6866
rect 19705 6851 19763 6857
rect 19705 6817 19717 6851
rect 19751 6817 19763 6851
rect 19705 6811 19763 6817
rect 18417 6647 18475 6653
rect 18417 6613 18429 6647
rect 18463 6613 18475 6647
rect 18417 6607 18475 6613
rect 18969 6647 19027 6653
rect 18969 6613 18981 6647
rect 19015 6644 19027 6647
rect 19150 6644 19156 6656
rect 19015 6616 19156 6644
rect 19015 6613 19027 6616
rect 18969 6607 19027 6613
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 19306 6644 19334 6811
rect 19720 6644 19748 6811
rect 19904 6780 19932 6888
rect 19996 6888 20076 6916
rect 19996 6857 20024 6888
rect 20070 6876 20076 6888
rect 20128 6876 20134 6928
rect 20364 6916 20392 6947
rect 20622 6944 20628 6996
rect 20680 6984 20686 6996
rect 20680 6956 20760 6984
rect 20680 6944 20686 6956
rect 20732 6916 20760 6956
rect 20898 6944 20904 6996
rect 20956 6944 20962 6996
rect 21818 6944 21824 6996
rect 21876 6944 21882 6996
rect 21836 6916 21864 6944
rect 20364 6888 20668 6916
rect 20732 6888 20944 6916
rect 20640 6860 20668 6888
rect 19981 6851 20039 6857
rect 19981 6817 19993 6851
rect 20027 6817 20039 6851
rect 19981 6811 20039 6817
rect 20441 6851 20499 6857
rect 20441 6817 20453 6851
rect 20487 6848 20499 6851
rect 20533 6851 20591 6857
rect 20533 6848 20545 6851
rect 20487 6820 20545 6848
rect 20487 6817 20499 6820
rect 20441 6811 20499 6817
rect 20533 6817 20545 6820
rect 20579 6817 20591 6851
rect 20533 6811 20591 6817
rect 20456 6780 20484 6811
rect 20622 6808 20628 6860
rect 20680 6848 20686 6860
rect 20809 6851 20867 6857
rect 20809 6848 20821 6851
rect 20680 6820 20821 6848
rect 20680 6808 20686 6820
rect 20809 6817 20821 6820
rect 20855 6817 20867 6851
rect 20809 6811 20867 6817
rect 19904 6752 20484 6780
rect 20916 6780 20944 6888
rect 21284 6888 21864 6916
rect 21082 6808 21088 6860
rect 21140 6848 21146 6860
rect 21284 6857 21312 6888
rect 21269 6851 21327 6857
rect 21269 6848 21281 6851
rect 21140 6820 21281 6848
rect 21140 6808 21146 6820
rect 21269 6817 21281 6820
rect 21315 6817 21327 6851
rect 21525 6851 21583 6857
rect 21525 6848 21537 6851
rect 21269 6811 21327 6817
rect 21376 6820 21537 6848
rect 21376 6780 21404 6820
rect 21525 6817 21537 6820
rect 21571 6817 21583 6851
rect 21525 6811 21583 6817
rect 20916 6752 21404 6780
rect 19904 6712 19932 6752
rect 20073 6715 20131 6721
rect 20073 6712 20085 6715
rect 19904 6684 20085 6712
rect 20073 6681 20085 6684
rect 20119 6681 20131 6715
rect 20073 6675 20131 6681
rect 19306 6616 19748 6644
rect 22649 6647 22707 6653
rect 22649 6613 22661 6647
rect 22695 6644 22707 6647
rect 28258 6644 28264 6656
rect 22695 6616 28264 6644
rect 22695 6613 22707 6616
rect 22649 6607 22707 6613
rect 28258 6604 28264 6616
rect 28316 6604 28322 6656
rect 552 6554 31372 6576
rect 552 6502 4250 6554
rect 4302 6502 4314 6554
rect 4366 6502 4378 6554
rect 4430 6502 4442 6554
rect 4494 6502 4506 6554
rect 4558 6502 11955 6554
rect 12007 6502 12019 6554
rect 12071 6502 12083 6554
rect 12135 6502 12147 6554
rect 12199 6502 12211 6554
rect 12263 6502 19660 6554
rect 19712 6502 19724 6554
rect 19776 6502 19788 6554
rect 19840 6502 19852 6554
rect 19904 6502 19916 6554
rect 19968 6502 27365 6554
rect 27417 6502 27429 6554
rect 27481 6502 27493 6554
rect 27545 6502 27557 6554
rect 27609 6502 27621 6554
rect 27673 6502 31372 6554
rect 552 6480 31372 6502
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 10192 6412 10609 6440
rect 10192 6400 10198 6412
rect 10597 6409 10609 6412
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 10686 6400 10692 6452
rect 10744 6400 10750 6452
rect 10965 6443 11023 6449
rect 10965 6409 10977 6443
rect 11011 6440 11023 6443
rect 11330 6440 11336 6452
rect 11011 6412 11336 6440
rect 11011 6409 11023 6412
rect 10965 6403 11023 6409
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 9732 6208 10425 6236
rect 9732 6196 9738 6208
rect 10413 6205 10425 6208
rect 10459 6236 10471 6239
rect 10502 6236 10508 6248
rect 10459 6208 10508 6236
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 10704 6245 10732 6400
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6236 10747 6239
rect 11057 6239 11115 6245
rect 11057 6236 11069 6239
rect 10735 6208 11069 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 11057 6205 11069 6208
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 10168 6171 10226 6177
rect 10168 6137 10180 6171
rect 10214 6168 10226 6171
rect 11164 6168 11192 6412
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 17034 6440 17040 6452
rect 16132 6412 17040 6440
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 11931 6208 14565 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 14553 6205 14565 6208
rect 14599 6236 14611 6239
rect 14642 6236 14648 6248
rect 14599 6208 14648 6236
rect 14599 6205 14611 6208
rect 14553 6199 14611 6205
rect 14642 6196 14648 6208
rect 14700 6196 14706 6248
rect 16132 6245 16160 6412
rect 17034 6400 17040 6412
rect 17092 6400 17098 6452
rect 18782 6400 18788 6452
rect 18840 6400 18846 6452
rect 20070 6400 20076 6452
rect 20128 6400 20134 6452
rect 17497 6375 17555 6381
rect 17497 6341 17509 6375
rect 17543 6372 17555 6375
rect 17862 6372 17868 6384
rect 17543 6344 17868 6372
rect 17543 6341 17555 6344
rect 17497 6335 17555 6341
rect 17862 6332 17868 6344
rect 17920 6332 17926 6384
rect 18800 6372 18828 6400
rect 17972 6344 18828 6372
rect 17770 6304 17776 6316
rect 17144 6276 17776 6304
rect 16117 6239 16175 6245
rect 16117 6205 16129 6239
rect 16163 6205 16175 6239
rect 16117 6199 16175 6205
rect 16384 6239 16442 6245
rect 16384 6205 16396 6239
rect 16430 6236 16442 6239
rect 17144 6236 17172 6276
rect 17770 6264 17776 6276
rect 17828 6304 17834 6316
rect 17972 6304 18000 6344
rect 17828 6276 18000 6304
rect 17828 6264 17834 6276
rect 17972 6245 18000 6276
rect 18322 6264 18328 6316
rect 18380 6304 18386 6316
rect 18785 6307 18843 6313
rect 18785 6304 18797 6307
rect 18380 6276 18797 6304
rect 18380 6264 18386 6276
rect 18785 6273 18797 6276
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 17681 6239 17739 6245
rect 17681 6236 17693 6239
rect 16430 6208 17172 6236
rect 17236 6208 17693 6236
rect 16430 6205 16442 6208
rect 16384 6199 16442 6205
rect 10214 6140 11192 6168
rect 12152 6171 12210 6177
rect 10214 6137 10226 6140
rect 10168 6131 10226 6137
rect 12152 6137 12164 6171
rect 12198 6168 12210 6171
rect 12526 6168 12532 6180
rect 12198 6140 12532 6168
rect 12198 6137 12210 6140
rect 12152 6131 12210 6137
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 14820 6171 14878 6177
rect 14820 6137 14832 6171
rect 14866 6168 14878 6171
rect 16206 6168 16212 6180
rect 14866 6140 16212 6168
rect 14866 6137 14878 6140
rect 14820 6131 14878 6137
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 17236 6112 17264 6208
rect 17681 6205 17693 6208
rect 17727 6205 17739 6239
rect 17681 6199 17739 6205
rect 17957 6239 18015 6245
rect 17957 6205 17969 6239
rect 18003 6205 18015 6239
rect 17957 6199 18015 6205
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6236 18107 6239
rect 18138 6236 18144 6248
rect 18095 6208 18144 6236
rect 18095 6205 18107 6208
rect 18049 6199 18107 6205
rect 9033 6103 9091 6109
rect 9033 6069 9045 6103
rect 9079 6100 9091 6103
rect 9674 6100 9680 6112
rect 9079 6072 9680 6100
rect 9079 6069 9091 6072
rect 9033 6063 9091 6069
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 13265 6103 13323 6109
rect 13265 6069 13277 6103
rect 13311 6100 13323 6103
rect 13538 6100 13544 6112
rect 13311 6072 13544 6100
rect 13311 6069 13323 6072
rect 13265 6063 13323 6069
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 15933 6103 15991 6109
rect 15933 6069 15945 6103
rect 15979 6100 15991 6103
rect 16758 6100 16764 6112
rect 15979 6072 16764 6100
rect 15979 6069 15991 6072
rect 15933 6063 15991 6069
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 17218 6060 17224 6112
rect 17276 6060 17282 6112
rect 17696 6100 17724 6199
rect 17773 6171 17831 6177
rect 17773 6137 17785 6171
rect 17819 6168 17831 6171
rect 18064 6168 18092 6199
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 19052 6239 19110 6245
rect 19052 6205 19064 6239
rect 19098 6236 19110 6239
rect 20088 6236 20116 6400
rect 19098 6208 20116 6236
rect 20349 6239 20407 6245
rect 19098 6205 19110 6208
rect 19052 6199 19110 6205
rect 18248 6168 18276 6199
rect 19260 6180 19288 6208
rect 20349 6205 20361 6239
rect 20395 6236 20407 6239
rect 21082 6236 21088 6248
rect 20395 6208 21088 6236
rect 20395 6205 20407 6208
rect 20349 6199 20407 6205
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 17819 6140 18092 6168
rect 18156 6140 18276 6168
rect 17819 6137 17831 6140
rect 17773 6131 17831 6137
rect 18156 6100 18184 6140
rect 19242 6128 19248 6180
rect 19300 6128 19306 6180
rect 20622 6177 20628 6180
rect 20616 6168 20628 6177
rect 20583 6140 20628 6168
rect 20616 6131 20628 6140
rect 20622 6128 20628 6131
rect 20680 6128 20686 6180
rect 17696 6072 18184 6100
rect 18230 6060 18236 6112
rect 18288 6100 18294 6112
rect 18325 6103 18383 6109
rect 18325 6100 18337 6103
rect 18288 6072 18337 6100
rect 18288 6060 18294 6072
rect 18325 6069 18337 6072
rect 18371 6069 18383 6103
rect 18325 6063 18383 6069
rect 20165 6103 20223 6109
rect 20165 6069 20177 6103
rect 20211 6100 20223 6103
rect 20438 6100 20444 6112
rect 20211 6072 20444 6100
rect 20211 6069 20223 6072
rect 20165 6063 20223 6069
rect 20438 6060 20444 6072
rect 20496 6060 20502 6112
rect 21726 6060 21732 6112
rect 21784 6060 21790 6112
rect 552 6010 31531 6032
rect 552 5958 8102 6010
rect 8154 5958 8166 6010
rect 8218 5958 8230 6010
rect 8282 5958 8294 6010
rect 8346 5958 8358 6010
rect 8410 5958 15807 6010
rect 15859 5958 15871 6010
rect 15923 5958 15935 6010
rect 15987 5958 15999 6010
rect 16051 5958 16063 6010
rect 16115 5958 23512 6010
rect 23564 5958 23576 6010
rect 23628 5958 23640 6010
rect 23692 5958 23704 6010
rect 23756 5958 23768 6010
rect 23820 5958 31217 6010
rect 31269 5958 31281 6010
rect 31333 5958 31345 6010
rect 31397 5958 31409 6010
rect 31461 5958 31473 6010
rect 31525 5958 31531 6010
rect 552 5936 31531 5958
rect 11606 5856 11612 5908
rect 11664 5856 11670 5908
rect 16206 5856 16212 5908
rect 16264 5896 16270 5908
rect 17129 5899 17187 5905
rect 17129 5896 17141 5899
rect 16264 5868 17141 5896
rect 16264 5856 16270 5868
rect 17129 5865 17141 5868
rect 17175 5896 17187 5899
rect 17218 5896 17224 5908
rect 17175 5868 17224 5896
rect 17175 5865 17187 5868
rect 17129 5859 17187 5865
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 17770 5856 17776 5908
rect 17828 5856 17834 5908
rect 18230 5856 18236 5908
rect 18288 5896 18294 5908
rect 18288 5868 18828 5896
rect 18288 5856 18294 5868
rect 11324 5831 11382 5837
rect 11324 5797 11336 5831
rect 11370 5828 11382 5831
rect 11624 5828 11652 5856
rect 11370 5800 11652 5828
rect 11370 5797 11382 5800
rect 11324 5791 11382 5797
rect 14642 5788 14648 5840
rect 14700 5828 14706 5840
rect 14700 5800 15332 5828
rect 14700 5788 14706 5800
rect 10502 5720 10508 5772
rect 10560 5760 10566 5772
rect 15304 5769 15332 5800
rect 16500 5800 17540 5828
rect 11057 5763 11115 5769
rect 11057 5760 11069 5763
rect 10560 5732 11069 5760
rect 10560 5720 10566 5732
rect 11057 5729 11069 5732
rect 11103 5729 11115 5763
rect 11057 5723 11115 5729
rect 15033 5763 15091 5769
rect 15033 5729 15045 5763
rect 15079 5760 15091 5763
rect 15289 5763 15347 5769
rect 15079 5732 15240 5760
rect 15079 5729 15091 5732
rect 15033 5723 15091 5729
rect 15212 5692 15240 5732
rect 15289 5729 15301 5763
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5760 16359 5763
rect 16393 5763 16451 5769
rect 16393 5760 16405 5763
rect 16347 5732 16405 5760
rect 16347 5729 16359 5732
rect 16301 5723 16359 5729
rect 16393 5729 16405 5732
rect 16439 5729 16451 5763
rect 16393 5723 16451 5729
rect 15212 5664 16160 5692
rect 16132 5624 16160 5664
rect 16206 5652 16212 5704
rect 16264 5692 16270 5704
rect 16316 5692 16344 5723
rect 16264 5664 16344 5692
rect 16264 5652 16270 5664
rect 16390 5624 16396 5636
rect 16132 5596 16396 5624
rect 16390 5584 16396 5596
rect 16448 5624 16454 5636
rect 16500 5633 16528 5800
rect 16945 5763 17003 5769
rect 16945 5729 16957 5763
rect 16991 5760 17003 5763
rect 17221 5763 17279 5769
rect 17221 5760 17233 5763
rect 16991 5732 17233 5760
rect 16991 5729 17003 5732
rect 16945 5723 17003 5729
rect 17221 5729 17233 5732
rect 17267 5760 17279 5763
rect 17402 5760 17408 5772
rect 17267 5732 17408 5760
rect 17267 5729 17279 5732
rect 17221 5723 17279 5729
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 17512 5769 17540 5800
rect 18138 5788 18144 5840
rect 18196 5788 18202 5840
rect 17497 5763 17555 5769
rect 17497 5729 17509 5763
rect 17543 5760 17555 5763
rect 17586 5760 17592 5772
rect 17543 5732 17592 5760
rect 17543 5729 17555 5732
rect 17497 5723 17555 5729
rect 17586 5720 17592 5732
rect 17644 5720 17650 5772
rect 17857 5769 17915 5775
rect 17857 5766 17869 5769
rect 17788 5738 17869 5766
rect 16485 5627 16543 5633
rect 16485 5624 16497 5627
rect 16448 5596 16497 5624
rect 16448 5584 16454 5596
rect 16485 5593 16497 5596
rect 16531 5593 16543 5627
rect 16485 5587 16543 5593
rect 16853 5627 16911 5633
rect 16853 5593 16865 5627
rect 16899 5624 16911 5627
rect 17678 5624 17684 5636
rect 16899 5596 17684 5624
rect 16899 5593 16911 5596
rect 16853 5587 16911 5593
rect 17678 5584 17684 5596
rect 17736 5584 17742 5636
rect 17788 5624 17816 5738
rect 17857 5735 17869 5738
rect 17903 5735 17915 5769
rect 17857 5729 17915 5735
rect 17954 5720 17960 5772
rect 18012 5758 18018 5772
rect 18156 5760 18184 5788
rect 18233 5763 18291 5769
rect 18233 5760 18245 5763
rect 18012 5730 18055 5758
rect 18156 5732 18245 5760
rect 18012 5720 18018 5730
rect 18233 5729 18245 5732
rect 18279 5729 18291 5763
rect 18233 5723 18291 5729
rect 18506 5720 18512 5772
rect 18564 5720 18570 5772
rect 18800 5769 18828 5868
rect 19150 5856 19156 5908
rect 19208 5856 19214 5908
rect 19242 5856 19248 5908
rect 19300 5856 19306 5908
rect 18877 5831 18935 5837
rect 18877 5797 18889 5831
rect 18923 5828 18935 5831
rect 19260 5828 19288 5856
rect 18923 5800 19288 5828
rect 18923 5797 18935 5800
rect 18877 5791 18935 5797
rect 18785 5763 18843 5769
rect 18785 5729 18797 5763
rect 18831 5729 18843 5763
rect 18785 5723 18843 5729
rect 18049 5627 18107 5633
rect 18049 5624 18061 5627
rect 17788 5596 18061 5624
rect 18049 5593 18061 5596
rect 18095 5624 18107 5627
rect 18230 5624 18236 5636
rect 18095 5596 18236 5624
rect 18095 5593 18107 5596
rect 18049 5587 18107 5593
rect 18230 5584 18236 5596
rect 18288 5584 18294 5636
rect 18325 5627 18383 5633
rect 18325 5593 18337 5627
rect 18371 5624 18383 5627
rect 18892 5624 18920 5791
rect 19260 5769 19288 5800
rect 19245 5763 19303 5769
rect 19245 5729 19257 5763
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 18371 5596 18920 5624
rect 18371 5593 18383 5596
rect 18325 5587 18383 5593
rect 12342 5516 12348 5568
rect 12400 5556 12406 5568
rect 12437 5559 12495 5565
rect 12437 5556 12449 5559
rect 12400 5528 12449 5556
rect 12400 5516 12406 5528
rect 12437 5525 12449 5528
rect 12483 5525 12495 5559
rect 12437 5519 12495 5525
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5556 13967 5559
rect 14182 5556 14188 5568
rect 13955 5528 14188 5556
rect 13955 5525 13967 5528
rect 13909 5519 13967 5525
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 17402 5516 17408 5568
rect 17460 5556 17466 5568
rect 18601 5559 18659 5565
rect 18601 5556 18613 5559
rect 17460 5528 18613 5556
rect 17460 5516 17466 5528
rect 18601 5525 18613 5528
rect 18647 5525 18659 5559
rect 18601 5519 18659 5525
rect 552 5466 31372 5488
rect 552 5414 4250 5466
rect 4302 5414 4314 5466
rect 4366 5414 4378 5466
rect 4430 5414 4442 5466
rect 4494 5414 4506 5466
rect 4558 5414 11955 5466
rect 12007 5414 12019 5466
rect 12071 5414 12083 5466
rect 12135 5414 12147 5466
rect 12199 5414 12211 5466
rect 12263 5414 19660 5466
rect 19712 5414 19724 5466
rect 19776 5414 19788 5466
rect 19840 5414 19852 5466
rect 19904 5414 19916 5466
rect 19968 5414 27365 5466
rect 27417 5414 27429 5466
rect 27481 5414 27493 5466
rect 27545 5414 27557 5466
rect 27609 5414 27621 5466
rect 27673 5414 31372 5466
rect 552 5392 31372 5414
rect 15841 5355 15899 5361
rect 15841 5321 15853 5355
rect 15887 5352 15899 5355
rect 16206 5352 16212 5364
rect 15887 5324 16212 5352
rect 15887 5321 15899 5324
rect 15841 5315 15899 5321
rect 16206 5312 16212 5324
rect 16264 5352 16270 5364
rect 16485 5355 16543 5361
rect 16485 5352 16497 5355
rect 16264 5324 16497 5352
rect 16264 5312 16270 5324
rect 16485 5321 16497 5324
rect 16531 5321 16543 5355
rect 16485 5315 16543 5321
rect 16592 5188 16804 5216
rect 15657 5151 15715 5157
rect 15657 5117 15669 5151
rect 15703 5148 15715 5151
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15703 5120 15761 5148
rect 15703 5117 15715 5120
rect 15657 5111 15715 5117
rect 15749 5117 15761 5120
rect 15795 5148 15807 5151
rect 16206 5148 16212 5160
rect 15795 5120 16212 5148
rect 15795 5117 15807 5120
rect 15749 5111 15807 5117
rect 16206 5108 16212 5120
rect 16264 5148 16270 5160
rect 16592 5157 16620 5188
rect 16776 5157 16804 5188
rect 17034 5176 17040 5228
rect 17092 5176 17098 5228
rect 16301 5151 16359 5157
rect 16301 5148 16313 5151
rect 16264 5120 16313 5148
rect 16264 5108 16270 5120
rect 16301 5117 16313 5120
rect 16347 5117 16359 5151
rect 16301 5111 16359 5117
rect 16577 5151 16635 5157
rect 16577 5117 16589 5151
rect 16623 5117 16635 5151
rect 16577 5111 16635 5117
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 16761 5151 16819 5157
rect 16761 5117 16773 5151
rect 16807 5148 16819 5151
rect 17304 5151 17362 5157
rect 17304 5148 17316 5151
rect 16807 5120 17316 5148
rect 16807 5117 16819 5120
rect 16761 5111 16819 5117
rect 17304 5117 17316 5120
rect 17350 5148 17362 5151
rect 18506 5148 18512 5160
rect 17350 5120 18512 5148
rect 17350 5117 17362 5120
rect 17304 5111 17362 5117
rect 15565 5083 15623 5089
rect 15565 5049 15577 5083
rect 15611 5080 15623 5083
rect 16482 5080 16488 5092
rect 15611 5052 16488 5080
rect 15611 5049 15623 5052
rect 15565 5043 15623 5049
rect 16482 5040 16488 5052
rect 16540 5080 16546 5092
rect 16684 5080 16712 5111
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 16540 5052 16712 5080
rect 16540 5040 16546 5052
rect 18417 5015 18475 5021
rect 18417 4981 18429 5015
rect 18463 5012 18475 5015
rect 21266 5012 21272 5024
rect 18463 4984 21272 5012
rect 18463 4981 18475 4984
rect 18417 4975 18475 4981
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 552 4922 31531 4944
rect 552 4870 8102 4922
rect 8154 4870 8166 4922
rect 8218 4870 8230 4922
rect 8282 4870 8294 4922
rect 8346 4870 8358 4922
rect 8410 4870 15807 4922
rect 15859 4870 15871 4922
rect 15923 4870 15935 4922
rect 15987 4870 15999 4922
rect 16051 4870 16063 4922
rect 16115 4870 23512 4922
rect 23564 4870 23576 4922
rect 23628 4870 23640 4922
rect 23692 4870 23704 4922
rect 23756 4870 23768 4922
rect 23820 4870 31217 4922
rect 31269 4870 31281 4922
rect 31333 4870 31345 4922
rect 31397 4870 31409 4922
rect 31461 4870 31473 4922
rect 31525 4870 31531 4922
rect 552 4848 31531 4870
rect 16390 4768 16396 4820
rect 16448 4768 16454 4820
rect 16482 4768 16488 4820
rect 16540 4768 16546 4820
rect 16500 4681 16528 4768
rect 16485 4675 16543 4681
rect 16485 4641 16497 4675
rect 16531 4641 16543 4675
rect 16485 4635 16543 4641
rect 552 4378 31372 4400
rect 552 4326 4250 4378
rect 4302 4326 4314 4378
rect 4366 4326 4378 4378
rect 4430 4326 4442 4378
rect 4494 4326 4506 4378
rect 4558 4326 11955 4378
rect 12007 4326 12019 4378
rect 12071 4326 12083 4378
rect 12135 4326 12147 4378
rect 12199 4326 12211 4378
rect 12263 4326 19660 4378
rect 19712 4326 19724 4378
rect 19776 4326 19788 4378
rect 19840 4326 19852 4378
rect 19904 4326 19916 4378
rect 19968 4326 27365 4378
rect 27417 4326 27429 4378
rect 27481 4326 27493 4378
rect 27545 4326 27557 4378
rect 27609 4326 27621 4378
rect 27673 4326 31372 4378
rect 552 4304 31372 4326
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 11238 4128 11244 4140
rect 10376 4100 11244 4128
rect 10376 4088 10382 4100
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 552 3834 31531 3856
rect 552 3782 8102 3834
rect 8154 3782 8166 3834
rect 8218 3782 8230 3834
rect 8282 3782 8294 3834
rect 8346 3782 8358 3834
rect 8410 3782 15807 3834
rect 15859 3782 15871 3834
rect 15923 3782 15935 3834
rect 15987 3782 15999 3834
rect 16051 3782 16063 3834
rect 16115 3782 23512 3834
rect 23564 3782 23576 3834
rect 23628 3782 23640 3834
rect 23692 3782 23704 3834
rect 23756 3782 23768 3834
rect 23820 3782 31217 3834
rect 31269 3782 31281 3834
rect 31333 3782 31345 3834
rect 31397 3782 31409 3834
rect 31461 3782 31473 3834
rect 31525 3782 31531 3834
rect 552 3760 31531 3782
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 12618 3448 12624 3460
rect 9088 3420 12624 3448
rect 9088 3408 9094 3420
rect 12618 3408 12624 3420
rect 12676 3408 12682 3460
rect 552 3290 31372 3312
rect 552 3238 4250 3290
rect 4302 3238 4314 3290
rect 4366 3238 4378 3290
rect 4430 3238 4442 3290
rect 4494 3238 4506 3290
rect 4558 3238 11955 3290
rect 12007 3238 12019 3290
rect 12071 3238 12083 3290
rect 12135 3238 12147 3290
rect 12199 3238 12211 3290
rect 12263 3238 19660 3290
rect 19712 3238 19724 3290
rect 19776 3238 19788 3290
rect 19840 3238 19852 3290
rect 19904 3238 19916 3290
rect 19968 3238 27365 3290
rect 27417 3238 27429 3290
rect 27481 3238 27493 3290
rect 27545 3238 27557 3290
rect 27609 3238 27621 3290
rect 27673 3238 31372 3290
rect 552 3216 31372 3238
rect 552 2746 31531 2768
rect 552 2694 8102 2746
rect 8154 2694 8166 2746
rect 8218 2694 8230 2746
rect 8282 2694 8294 2746
rect 8346 2694 8358 2746
rect 8410 2694 15807 2746
rect 15859 2694 15871 2746
rect 15923 2694 15935 2746
rect 15987 2694 15999 2746
rect 16051 2694 16063 2746
rect 16115 2694 23512 2746
rect 23564 2694 23576 2746
rect 23628 2694 23640 2746
rect 23692 2694 23704 2746
rect 23756 2694 23768 2746
rect 23820 2694 31217 2746
rect 31269 2694 31281 2746
rect 31333 2694 31345 2746
rect 31397 2694 31409 2746
rect 31461 2694 31473 2746
rect 31525 2694 31531 2746
rect 552 2672 31531 2694
rect 552 2202 31372 2224
rect 552 2150 4250 2202
rect 4302 2150 4314 2202
rect 4366 2150 4378 2202
rect 4430 2150 4442 2202
rect 4494 2150 4506 2202
rect 4558 2150 11955 2202
rect 12007 2150 12019 2202
rect 12071 2150 12083 2202
rect 12135 2150 12147 2202
rect 12199 2150 12211 2202
rect 12263 2150 19660 2202
rect 19712 2150 19724 2202
rect 19776 2150 19788 2202
rect 19840 2150 19852 2202
rect 19904 2150 19916 2202
rect 19968 2150 27365 2202
rect 27417 2150 27429 2202
rect 27481 2150 27493 2202
rect 27545 2150 27557 2202
rect 27609 2150 27621 2202
rect 27673 2150 31372 2202
rect 552 2128 31372 2150
rect 552 1658 31531 1680
rect 552 1606 8102 1658
rect 8154 1606 8166 1658
rect 8218 1606 8230 1658
rect 8282 1606 8294 1658
rect 8346 1606 8358 1658
rect 8410 1606 15807 1658
rect 15859 1606 15871 1658
rect 15923 1606 15935 1658
rect 15987 1606 15999 1658
rect 16051 1606 16063 1658
rect 16115 1606 23512 1658
rect 23564 1606 23576 1658
rect 23628 1606 23640 1658
rect 23692 1606 23704 1658
rect 23756 1606 23768 1658
rect 23820 1606 31217 1658
rect 31269 1606 31281 1658
rect 31333 1606 31345 1658
rect 31397 1606 31409 1658
rect 31461 1606 31473 1658
rect 31525 1606 31531 1658
rect 552 1584 31531 1606
rect 552 1114 31372 1136
rect 552 1062 4250 1114
rect 4302 1062 4314 1114
rect 4366 1062 4378 1114
rect 4430 1062 4442 1114
rect 4494 1062 4506 1114
rect 4558 1062 11955 1114
rect 12007 1062 12019 1114
rect 12071 1062 12083 1114
rect 12135 1062 12147 1114
rect 12199 1062 12211 1114
rect 12263 1062 19660 1114
rect 19712 1062 19724 1114
rect 19776 1062 19788 1114
rect 19840 1062 19852 1114
rect 19904 1062 19916 1114
rect 19968 1062 27365 1114
rect 27417 1062 27429 1114
rect 27481 1062 27493 1114
rect 27545 1062 27557 1114
rect 27609 1062 27621 1114
rect 27673 1062 31372 1114
rect 552 1040 31372 1062
rect 16206 824 16212 876
rect 16264 864 16270 876
rect 22925 867 22983 873
rect 22925 864 22937 867
rect 16264 836 22937 864
rect 16264 824 16270 836
rect 22925 833 22937 836
rect 22971 833 22983 867
rect 22925 827 22983 833
rect 22646 756 22652 808
rect 22704 756 22710 808
rect 552 570 31531 592
rect 552 518 8102 570
rect 8154 518 8166 570
rect 8218 518 8230 570
rect 8282 518 8294 570
rect 8346 518 8358 570
rect 8410 518 15807 570
rect 15859 518 15871 570
rect 15923 518 15935 570
rect 15987 518 15999 570
rect 16051 518 16063 570
rect 16115 518 23512 570
rect 23564 518 23576 570
rect 23628 518 23640 570
rect 23692 518 23704 570
rect 23756 518 23768 570
rect 23820 518 31217 570
rect 31269 518 31281 570
rect 31333 518 31345 570
rect 31397 518 31409 570
rect 31461 518 31473 570
rect 31525 518 31531 570
rect 552 496 31531 518
rect 16022 416 16028 468
rect 16080 456 16086 468
rect 16298 456 16304 468
rect 16080 428 16304 456
rect 16080 416 16086 428
rect 16298 416 16304 428
rect 16356 416 16362 468
<< via1 >>
rect 8102 19014 8154 19066
rect 8166 19014 8218 19066
rect 8230 19014 8282 19066
rect 8294 19014 8346 19066
rect 8358 19014 8410 19066
rect 15807 19014 15859 19066
rect 15871 19014 15923 19066
rect 15935 19014 15987 19066
rect 15999 19014 16051 19066
rect 16063 19014 16115 19066
rect 23512 19014 23564 19066
rect 23576 19014 23628 19066
rect 23640 19014 23692 19066
rect 23704 19014 23756 19066
rect 23768 19014 23820 19066
rect 31217 19014 31269 19066
rect 31281 19014 31333 19066
rect 31345 19014 31397 19066
rect 31409 19014 31461 19066
rect 31473 19014 31525 19066
rect 4250 18470 4302 18522
rect 4314 18470 4366 18522
rect 4378 18470 4430 18522
rect 4442 18470 4494 18522
rect 4506 18470 4558 18522
rect 11955 18470 12007 18522
rect 12019 18470 12071 18522
rect 12083 18470 12135 18522
rect 12147 18470 12199 18522
rect 12211 18470 12263 18522
rect 19660 18470 19712 18522
rect 19724 18470 19776 18522
rect 19788 18470 19840 18522
rect 19852 18470 19904 18522
rect 19916 18470 19968 18522
rect 27365 18470 27417 18522
rect 27429 18470 27481 18522
rect 27493 18470 27545 18522
rect 27557 18470 27609 18522
rect 27621 18470 27673 18522
rect 8102 17926 8154 17978
rect 8166 17926 8218 17978
rect 8230 17926 8282 17978
rect 8294 17926 8346 17978
rect 8358 17926 8410 17978
rect 15807 17926 15859 17978
rect 15871 17926 15923 17978
rect 15935 17926 15987 17978
rect 15999 17926 16051 17978
rect 16063 17926 16115 17978
rect 23512 17926 23564 17978
rect 23576 17926 23628 17978
rect 23640 17926 23692 17978
rect 23704 17926 23756 17978
rect 23768 17926 23820 17978
rect 31217 17926 31269 17978
rect 31281 17926 31333 17978
rect 31345 17926 31397 17978
rect 31409 17926 31461 17978
rect 31473 17926 31525 17978
rect 4250 17382 4302 17434
rect 4314 17382 4366 17434
rect 4378 17382 4430 17434
rect 4442 17382 4494 17434
rect 4506 17382 4558 17434
rect 11955 17382 12007 17434
rect 12019 17382 12071 17434
rect 12083 17382 12135 17434
rect 12147 17382 12199 17434
rect 12211 17382 12263 17434
rect 19660 17382 19712 17434
rect 19724 17382 19776 17434
rect 19788 17382 19840 17434
rect 19852 17382 19904 17434
rect 19916 17382 19968 17434
rect 27365 17382 27417 17434
rect 27429 17382 27481 17434
rect 27493 17382 27545 17434
rect 27557 17382 27609 17434
rect 27621 17382 27673 17434
rect 8102 16838 8154 16890
rect 8166 16838 8218 16890
rect 8230 16838 8282 16890
rect 8294 16838 8346 16890
rect 8358 16838 8410 16890
rect 15807 16838 15859 16890
rect 15871 16838 15923 16890
rect 15935 16838 15987 16890
rect 15999 16838 16051 16890
rect 16063 16838 16115 16890
rect 23512 16838 23564 16890
rect 23576 16838 23628 16890
rect 23640 16838 23692 16890
rect 23704 16838 23756 16890
rect 23768 16838 23820 16890
rect 31217 16838 31269 16890
rect 31281 16838 31333 16890
rect 31345 16838 31397 16890
rect 31409 16838 31461 16890
rect 31473 16838 31525 16890
rect 4250 16294 4302 16346
rect 4314 16294 4366 16346
rect 4378 16294 4430 16346
rect 4442 16294 4494 16346
rect 4506 16294 4558 16346
rect 11955 16294 12007 16346
rect 12019 16294 12071 16346
rect 12083 16294 12135 16346
rect 12147 16294 12199 16346
rect 12211 16294 12263 16346
rect 19660 16294 19712 16346
rect 19724 16294 19776 16346
rect 19788 16294 19840 16346
rect 19852 16294 19904 16346
rect 19916 16294 19968 16346
rect 27365 16294 27417 16346
rect 27429 16294 27481 16346
rect 27493 16294 27545 16346
rect 27557 16294 27609 16346
rect 27621 16294 27673 16346
rect 8102 15750 8154 15802
rect 8166 15750 8218 15802
rect 8230 15750 8282 15802
rect 8294 15750 8346 15802
rect 8358 15750 8410 15802
rect 15807 15750 15859 15802
rect 15871 15750 15923 15802
rect 15935 15750 15987 15802
rect 15999 15750 16051 15802
rect 16063 15750 16115 15802
rect 23512 15750 23564 15802
rect 23576 15750 23628 15802
rect 23640 15750 23692 15802
rect 23704 15750 23756 15802
rect 23768 15750 23820 15802
rect 31217 15750 31269 15802
rect 31281 15750 31333 15802
rect 31345 15750 31397 15802
rect 31409 15750 31461 15802
rect 31473 15750 31525 15802
rect 4250 15206 4302 15258
rect 4314 15206 4366 15258
rect 4378 15206 4430 15258
rect 4442 15206 4494 15258
rect 4506 15206 4558 15258
rect 11955 15206 12007 15258
rect 12019 15206 12071 15258
rect 12083 15206 12135 15258
rect 12147 15206 12199 15258
rect 12211 15206 12263 15258
rect 19660 15206 19712 15258
rect 19724 15206 19776 15258
rect 19788 15206 19840 15258
rect 19852 15206 19904 15258
rect 19916 15206 19968 15258
rect 27365 15206 27417 15258
rect 27429 15206 27481 15258
rect 27493 15206 27545 15258
rect 27557 15206 27609 15258
rect 27621 15206 27673 15258
rect 8102 14662 8154 14714
rect 8166 14662 8218 14714
rect 8230 14662 8282 14714
rect 8294 14662 8346 14714
rect 8358 14662 8410 14714
rect 15807 14662 15859 14714
rect 15871 14662 15923 14714
rect 15935 14662 15987 14714
rect 15999 14662 16051 14714
rect 16063 14662 16115 14714
rect 23512 14662 23564 14714
rect 23576 14662 23628 14714
rect 23640 14662 23692 14714
rect 23704 14662 23756 14714
rect 23768 14662 23820 14714
rect 31217 14662 31269 14714
rect 31281 14662 31333 14714
rect 31345 14662 31397 14714
rect 31409 14662 31461 14714
rect 31473 14662 31525 14714
rect 14188 14560 14240 14612
rect 16764 14560 16816 14612
rect 13176 14467 13228 14476
rect 13176 14433 13210 14467
rect 13210 14433 13228 14467
rect 13176 14424 13228 14433
rect 14464 14467 14516 14476
rect 14464 14433 14473 14467
rect 14473 14433 14507 14467
rect 14507 14433 14516 14467
rect 14464 14424 14516 14433
rect 14740 14467 14792 14476
rect 14740 14433 14774 14467
rect 14774 14433 14792 14467
rect 14740 14424 14792 14433
rect 18604 14424 18656 14476
rect 19432 14220 19484 14272
rect 4250 14118 4302 14170
rect 4314 14118 4366 14170
rect 4378 14118 4430 14170
rect 4442 14118 4494 14170
rect 4506 14118 4558 14170
rect 11955 14118 12007 14170
rect 12019 14118 12071 14170
rect 12083 14118 12135 14170
rect 12147 14118 12199 14170
rect 12211 14118 12263 14170
rect 19660 14118 19712 14170
rect 19724 14118 19776 14170
rect 19788 14118 19840 14170
rect 19852 14118 19904 14170
rect 19916 14118 19968 14170
rect 27365 14118 27417 14170
rect 27429 14118 27481 14170
rect 27493 14118 27545 14170
rect 27557 14118 27609 14170
rect 27621 14118 27673 14170
rect 12440 14016 12492 14068
rect 14740 14016 14792 14068
rect 18052 14016 18104 14068
rect 20628 14016 20680 14068
rect 13176 13880 13228 13932
rect 11336 13812 11388 13864
rect 11428 13855 11480 13864
rect 11428 13821 11437 13855
rect 11437 13821 11471 13855
rect 11471 13821 11480 13855
rect 11428 13812 11480 13821
rect 13452 13812 13504 13864
rect 16488 13787 16540 13796
rect 10692 13676 10744 13728
rect 11152 13676 11204 13728
rect 14004 13719 14056 13728
rect 14004 13685 14013 13719
rect 14013 13685 14047 13719
rect 14047 13685 14056 13719
rect 14004 13676 14056 13685
rect 14372 13676 14424 13728
rect 16488 13753 16500 13787
rect 16500 13753 16540 13787
rect 16488 13744 16540 13753
rect 17776 13855 17828 13864
rect 17776 13821 17785 13855
rect 17785 13821 17819 13855
rect 17819 13821 17828 13855
rect 17776 13812 17828 13821
rect 17960 13812 18012 13864
rect 18604 13812 18656 13864
rect 18696 13855 18748 13864
rect 18696 13821 18705 13855
rect 18705 13821 18739 13855
rect 18739 13821 18748 13855
rect 18696 13812 18748 13821
rect 18972 13855 19024 13864
rect 18972 13821 18995 13855
rect 18995 13821 19024 13855
rect 18972 13812 19024 13821
rect 19432 13812 19484 13864
rect 15660 13676 15712 13728
rect 20444 13719 20496 13728
rect 20444 13685 20453 13719
rect 20453 13685 20487 13719
rect 20487 13685 20496 13719
rect 20444 13676 20496 13685
rect 20628 13676 20680 13728
rect 8102 13574 8154 13626
rect 8166 13574 8218 13626
rect 8230 13574 8282 13626
rect 8294 13574 8346 13626
rect 8358 13574 8410 13626
rect 15807 13574 15859 13626
rect 15871 13574 15923 13626
rect 15935 13574 15987 13626
rect 15999 13574 16051 13626
rect 16063 13574 16115 13626
rect 23512 13574 23564 13626
rect 23576 13574 23628 13626
rect 23640 13574 23692 13626
rect 23704 13574 23756 13626
rect 23768 13574 23820 13626
rect 31217 13574 31269 13626
rect 31281 13574 31333 13626
rect 31345 13574 31397 13626
rect 31409 13574 31461 13626
rect 31473 13574 31525 13626
rect 11428 13472 11480 13524
rect 13452 13472 13504 13524
rect 14004 13515 14056 13524
rect 14004 13481 14013 13515
rect 14013 13481 14047 13515
rect 14047 13481 14056 13515
rect 14004 13472 14056 13481
rect 14740 13472 14792 13524
rect 11152 13404 11204 13456
rect 13176 13404 13228 13456
rect 10140 13132 10192 13184
rect 11060 13175 11112 13184
rect 11060 13141 11069 13175
rect 11069 13141 11103 13175
rect 11103 13141 11112 13175
rect 11060 13132 11112 13141
rect 11244 13200 11296 13252
rect 11796 13175 11848 13184
rect 11796 13141 11805 13175
rect 11805 13141 11839 13175
rect 11839 13141 11848 13175
rect 11796 13132 11848 13141
rect 14004 13336 14056 13388
rect 16488 13472 16540 13524
rect 16304 13336 16356 13388
rect 15568 13268 15620 13320
rect 15660 13268 15712 13320
rect 17776 13472 17828 13524
rect 19984 13472 20036 13524
rect 21916 13472 21968 13524
rect 18696 13404 18748 13456
rect 20628 13404 20680 13456
rect 17868 13379 17920 13388
rect 17868 13345 17891 13379
rect 17891 13345 17920 13379
rect 17868 13336 17920 13345
rect 19524 13379 19576 13388
rect 19524 13345 19533 13379
rect 19533 13345 19567 13379
rect 19567 13345 19576 13379
rect 19524 13336 19576 13345
rect 19616 13379 19668 13388
rect 19616 13345 19625 13379
rect 19625 13345 19659 13379
rect 19659 13345 19668 13379
rect 19616 13336 19668 13345
rect 19432 13268 19484 13320
rect 14372 13200 14424 13252
rect 14004 13132 14056 13184
rect 16764 13132 16816 13184
rect 4250 13030 4302 13082
rect 4314 13030 4366 13082
rect 4378 13030 4430 13082
rect 4442 13030 4494 13082
rect 4506 13030 4558 13082
rect 11955 13030 12007 13082
rect 12019 13030 12071 13082
rect 12083 13030 12135 13082
rect 12147 13030 12199 13082
rect 12211 13030 12263 13082
rect 19660 13030 19712 13082
rect 19724 13030 19776 13082
rect 19788 13030 19840 13082
rect 19852 13030 19904 13082
rect 19916 13030 19968 13082
rect 27365 13030 27417 13082
rect 27429 13030 27481 13082
rect 27493 13030 27545 13082
rect 27557 13030 27609 13082
rect 27621 13030 27673 13082
rect 10784 12928 10836 12980
rect 11060 12928 11112 12980
rect 11520 12928 11572 12980
rect 11152 12767 11204 12776
rect 11152 12733 11170 12767
rect 11170 12733 11204 12767
rect 11152 12724 11204 12733
rect 11336 12724 11388 12776
rect 11796 12792 11848 12844
rect 11888 12724 11940 12776
rect 18512 12928 18564 12980
rect 18604 12928 18656 12980
rect 19432 12928 19484 12980
rect 20444 12971 20496 12980
rect 20444 12937 20453 12971
rect 20453 12937 20487 12971
rect 20487 12937 20496 12971
rect 20444 12928 20496 12937
rect 28264 12928 28316 12980
rect 28540 12928 28592 12980
rect 31668 12928 31720 12980
rect 18696 12860 18748 12912
rect 19524 12860 19576 12912
rect 20168 12860 20220 12912
rect 27988 12860 28040 12912
rect 14464 12792 14516 12844
rect 16488 12699 16540 12708
rect 16488 12665 16497 12699
rect 16497 12665 16531 12699
rect 16531 12665 16540 12699
rect 16488 12656 16540 12665
rect 10692 12588 10744 12640
rect 14004 12588 14056 12640
rect 16764 12588 16816 12640
rect 18972 12724 19024 12776
rect 19984 12792 20036 12844
rect 20536 12792 20588 12844
rect 22192 12767 22244 12776
rect 22192 12733 22201 12767
rect 22201 12733 22235 12767
rect 22235 12733 22244 12767
rect 22192 12724 22244 12733
rect 20444 12656 20496 12708
rect 19892 12631 19944 12640
rect 19892 12597 19901 12631
rect 19901 12597 19935 12631
rect 19935 12597 19944 12631
rect 19892 12588 19944 12597
rect 20168 12631 20220 12640
rect 20168 12597 20177 12631
rect 20177 12597 20211 12631
rect 20211 12597 20220 12631
rect 20168 12588 20220 12597
rect 20628 12588 20680 12640
rect 8102 12486 8154 12538
rect 8166 12486 8218 12538
rect 8230 12486 8282 12538
rect 8294 12486 8346 12538
rect 8358 12486 8410 12538
rect 15807 12486 15859 12538
rect 15871 12486 15923 12538
rect 15935 12486 15987 12538
rect 15999 12486 16051 12538
rect 16063 12486 16115 12538
rect 23512 12486 23564 12538
rect 23576 12486 23628 12538
rect 23640 12486 23692 12538
rect 23704 12486 23756 12538
rect 23768 12486 23820 12538
rect 31217 12486 31269 12538
rect 31281 12486 31333 12538
rect 31345 12486 31397 12538
rect 31409 12486 31461 12538
rect 31473 12486 31525 12538
rect 6920 12384 6972 12436
rect 11244 12384 11296 12436
rect 11796 12384 11848 12436
rect 12900 12384 12952 12436
rect 14832 12384 14884 12436
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 16764 12384 16816 12436
rect 18696 12384 18748 12436
rect 19892 12384 19944 12436
rect 11888 12316 11940 12368
rect 9680 12248 9732 12300
rect 10140 12291 10192 12300
rect 10140 12257 10158 12291
rect 10158 12257 10192 12291
rect 10140 12248 10192 12257
rect 10508 12180 10560 12232
rect 10968 12291 11020 12300
rect 10968 12257 10977 12291
rect 10977 12257 11011 12291
rect 11011 12257 11020 12291
rect 10968 12248 11020 12257
rect 11428 12291 11480 12300
rect 11428 12257 11437 12291
rect 11437 12257 11471 12291
rect 11471 12257 11480 12291
rect 11428 12248 11480 12257
rect 12256 12248 12308 12300
rect 14096 12316 14148 12368
rect 14004 12291 14056 12300
rect 14004 12257 14038 12291
rect 14038 12257 14056 12291
rect 14004 12248 14056 12257
rect 14464 12248 14516 12300
rect 15568 12291 15620 12300
rect 15568 12257 15577 12291
rect 15577 12257 15611 12291
rect 15611 12257 15620 12291
rect 15568 12248 15620 12257
rect 16212 12291 16264 12300
rect 16212 12257 16221 12291
rect 16221 12257 16255 12291
rect 16255 12257 16264 12291
rect 16212 12248 16264 12257
rect 16488 12248 16540 12300
rect 17592 12248 17644 12300
rect 19432 12248 19484 12300
rect 20444 12384 20496 12436
rect 22192 12384 22244 12436
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 20628 12291 20680 12300
rect 20628 12257 20637 12291
rect 20637 12257 20671 12291
rect 20671 12257 20680 12291
rect 20628 12248 20680 12257
rect 20720 12291 20772 12300
rect 20720 12257 20729 12291
rect 20729 12257 20763 12291
rect 20763 12257 20772 12291
rect 20720 12248 20772 12257
rect 21548 12291 21600 12300
rect 21548 12257 21557 12291
rect 21557 12257 21591 12291
rect 21591 12257 21600 12291
rect 21548 12248 21600 12257
rect 28448 12384 28500 12436
rect 22928 12248 22980 12300
rect 20352 12112 20404 12164
rect 12440 12044 12492 12096
rect 19524 12044 19576 12096
rect 20628 12044 20680 12096
rect 20996 12044 21048 12096
rect 28264 12044 28316 12096
rect 4250 11942 4302 11994
rect 4314 11942 4366 11994
rect 4378 11942 4430 11994
rect 4442 11942 4494 11994
rect 4506 11942 4558 11994
rect 11955 11942 12007 11994
rect 12019 11942 12071 11994
rect 12083 11942 12135 11994
rect 12147 11942 12199 11994
rect 12211 11942 12263 11994
rect 19660 11942 19712 11994
rect 19724 11942 19776 11994
rect 19788 11942 19840 11994
rect 19852 11942 19904 11994
rect 19916 11942 19968 11994
rect 27365 11942 27417 11994
rect 27429 11942 27481 11994
rect 27493 11942 27545 11994
rect 27557 11942 27609 11994
rect 27621 11942 27673 11994
rect 10140 11840 10192 11892
rect 11428 11840 11480 11892
rect 12348 11840 12400 11892
rect 15476 11840 15528 11892
rect 19340 11840 19392 11892
rect 19524 11840 19576 11892
rect 20352 11840 20404 11892
rect 20628 11840 20680 11892
rect 20904 11840 20956 11892
rect 9036 11679 9088 11688
rect 9036 11645 9045 11679
rect 9045 11645 9079 11679
rect 9079 11645 9088 11679
rect 9036 11636 9088 11645
rect 10692 11704 10744 11756
rect 12440 11815 12492 11824
rect 12440 11781 12449 11815
rect 12449 11781 12483 11815
rect 12483 11781 12492 11815
rect 12440 11772 12492 11781
rect 9128 11611 9180 11620
rect 9128 11577 9137 11611
rect 9137 11577 9171 11611
rect 9171 11577 9180 11611
rect 9128 11568 9180 11577
rect 9864 11611 9916 11620
rect 9864 11577 9873 11611
rect 9873 11577 9907 11611
rect 9907 11577 9916 11611
rect 9864 11568 9916 11577
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 10508 11500 10560 11552
rect 11336 11500 11388 11552
rect 11796 11500 11848 11552
rect 18696 11704 18748 11756
rect 14096 11636 14148 11688
rect 18052 11636 18104 11688
rect 28540 11840 28592 11892
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 12900 11500 12952 11552
rect 19340 11500 19392 11552
rect 22008 11568 22060 11620
rect 21088 11543 21140 11552
rect 21088 11509 21097 11543
rect 21097 11509 21131 11543
rect 21131 11509 21140 11543
rect 21088 11500 21140 11509
rect 21364 11543 21416 11552
rect 21364 11509 21373 11543
rect 21373 11509 21407 11543
rect 21407 11509 21416 11543
rect 21364 11500 21416 11509
rect 8102 11398 8154 11450
rect 8166 11398 8218 11450
rect 8230 11398 8282 11450
rect 8294 11398 8346 11450
rect 8358 11398 8410 11450
rect 15807 11398 15859 11450
rect 15871 11398 15923 11450
rect 15935 11398 15987 11450
rect 15999 11398 16051 11450
rect 16063 11398 16115 11450
rect 23512 11398 23564 11450
rect 23576 11398 23628 11450
rect 23640 11398 23692 11450
rect 23704 11398 23756 11450
rect 23768 11398 23820 11450
rect 31217 11398 31269 11450
rect 31281 11398 31333 11450
rect 31345 11398 31397 11450
rect 31409 11398 31461 11450
rect 31473 11398 31525 11450
rect 6920 11296 6972 11348
rect 9128 11296 9180 11348
rect 9036 11228 9088 11280
rect 9680 11296 9732 11348
rect 10140 11203 10192 11212
rect 10140 11169 10149 11203
rect 10149 11169 10183 11203
rect 10183 11169 10192 11203
rect 10140 11160 10192 11169
rect 10968 11296 11020 11348
rect 11612 11296 11664 11348
rect 13544 11296 13596 11348
rect 16212 11296 16264 11348
rect 17408 11296 17460 11348
rect 20904 11339 20956 11348
rect 20904 11305 20913 11339
rect 20913 11305 20947 11339
rect 20947 11305 20956 11339
rect 20904 11296 20956 11305
rect 20996 11296 21048 11348
rect 21088 11296 21140 11348
rect 11796 11228 11848 11280
rect 10968 11160 11020 11212
rect 12900 11160 12952 11212
rect 14096 11160 14148 11212
rect 14648 11203 14700 11212
rect 14648 11169 14682 11203
rect 14682 11169 14700 11203
rect 14648 11160 14700 11169
rect 10784 11092 10836 11144
rect 9680 11024 9732 11076
rect 18052 11160 18104 11212
rect 20536 11160 20588 11212
rect 21640 11271 21692 11280
rect 21640 11237 21649 11271
rect 21649 11237 21683 11271
rect 21683 11237 21692 11271
rect 21640 11228 21692 11237
rect 21364 11160 21416 11212
rect 19340 11135 19392 11144
rect 19340 11101 19349 11135
rect 19349 11101 19383 11135
rect 19383 11101 19392 11135
rect 22008 11160 22060 11212
rect 28264 11296 28316 11348
rect 19340 11092 19392 11101
rect 22192 11067 22244 11076
rect 15292 10956 15344 11008
rect 22192 11033 22201 11067
rect 22201 11033 22235 11067
rect 22235 11033 22244 11067
rect 22928 11135 22980 11144
rect 22928 11101 22937 11135
rect 22937 11101 22971 11135
rect 22971 11101 22980 11135
rect 22928 11092 22980 11101
rect 22192 11024 22244 11033
rect 22744 10999 22796 11008
rect 22744 10965 22753 10999
rect 22753 10965 22787 10999
rect 22787 10965 22796 10999
rect 22744 10956 22796 10965
rect 4250 10854 4302 10906
rect 4314 10854 4366 10906
rect 4378 10854 4430 10906
rect 4442 10854 4494 10906
rect 4506 10854 4558 10906
rect 11955 10854 12007 10906
rect 12019 10854 12071 10906
rect 12083 10854 12135 10906
rect 12147 10854 12199 10906
rect 12211 10854 12263 10906
rect 19660 10854 19712 10906
rect 19724 10854 19776 10906
rect 19788 10854 19840 10906
rect 19852 10854 19904 10906
rect 19916 10854 19968 10906
rect 27365 10854 27417 10906
rect 27429 10854 27481 10906
rect 27493 10854 27545 10906
rect 27557 10854 27609 10906
rect 27621 10854 27673 10906
rect 10140 10752 10192 10804
rect 10968 10752 11020 10804
rect 11152 10752 11204 10804
rect 21272 10752 21324 10804
rect 9680 10684 9732 10736
rect 14648 10684 14700 10736
rect 22100 10684 22152 10736
rect 22744 10684 22796 10736
rect 9036 10616 9088 10668
rect 10508 10659 10560 10668
rect 10508 10625 10517 10659
rect 10517 10625 10551 10659
rect 10551 10625 10560 10659
rect 10508 10616 10560 10625
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 9772 10548 9824 10600
rect 15292 10548 15344 10600
rect 16580 10616 16632 10668
rect 18052 10616 18104 10668
rect 22284 10659 22336 10668
rect 22284 10625 22293 10659
rect 22293 10625 22327 10659
rect 22327 10625 22336 10659
rect 22284 10616 22336 10625
rect 21640 10591 21692 10600
rect 21640 10557 21649 10591
rect 21649 10557 21683 10591
rect 21683 10557 21692 10591
rect 21640 10548 21692 10557
rect 22192 10548 22244 10600
rect 22744 10591 22796 10600
rect 22744 10557 22753 10591
rect 22753 10557 22787 10591
rect 22787 10557 22796 10591
rect 22744 10548 22796 10557
rect 9036 10412 9088 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 14464 10412 14516 10464
rect 15384 10412 15436 10464
rect 22008 10480 22060 10532
rect 22192 10412 22244 10464
rect 22836 10455 22888 10464
rect 22836 10421 22845 10455
rect 22845 10421 22879 10455
rect 22879 10421 22888 10455
rect 22836 10412 22888 10421
rect 8102 10310 8154 10362
rect 8166 10310 8218 10362
rect 8230 10310 8282 10362
rect 8294 10310 8346 10362
rect 8358 10310 8410 10362
rect 15807 10310 15859 10362
rect 15871 10310 15923 10362
rect 15935 10310 15987 10362
rect 15999 10310 16051 10362
rect 16063 10310 16115 10362
rect 23512 10310 23564 10362
rect 23576 10310 23628 10362
rect 23640 10310 23692 10362
rect 23704 10310 23756 10362
rect 23768 10310 23820 10362
rect 31217 10310 31269 10362
rect 31281 10310 31333 10362
rect 31345 10310 31397 10362
rect 31409 10310 31461 10362
rect 31473 10310 31525 10362
rect 7104 10251 7156 10260
rect 7104 10217 7113 10251
rect 7113 10217 7147 10251
rect 7147 10217 7156 10251
rect 7104 10208 7156 10217
rect 8392 10072 8444 10124
rect 9680 10208 9732 10260
rect 9772 10208 9824 10260
rect 14464 10208 14516 10260
rect 15384 10208 15436 10260
rect 9588 10183 9640 10192
rect 9588 10149 9597 10183
rect 9597 10149 9631 10183
rect 9631 10149 9640 10183
rect 9588 10140 9640 10149
rect 8852 10115 8904 10124
rect 8852 10081 8861 10115
rect 8861 10081 8895 10115
rect 8895 10081 8904 10115
rect 8852 10072 8904 10081
rect 9036 10047 9088 10056
rect 9036 10013 9045 10047
rect 9045 10013 9079 10047
rect 9079 10013 9088 10047
rect 9036 10004 9088 10013
rect 9956 10004 10008 10056
rect 13820 10004 13872 10056
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 14648 10115 14700 10124
rect 14648 10081 14657 10115
rect 14657 10081 14691 10115
rect 14691 10081 14700 10115
rect 14648 10072 14700 10081
rect 15292 10072 15344 10124
rect 15936 10115 15988 10124
rect 15936 10081 15945 10115
rect 15945 10081 15979 10115
rect 15979 10081 15988 10115
rect 15936 10072 15988 10081
rect 18052 10072 18104 10124
rect 18144 10115 18196 10124
rect 18144 10081 18153 10115
rect 18153 10081 18187 10115
rect 18187 10081 18196 10115
rect 22192 10208 22244 10260
rect 22284 10208 22336 10260
rect 22836 10208 22888 10260
rect 28264 10208 28316 10260
rect 18144 10072 18196 10081
rect 7196 9868 7248 9920
rect 12624 9911 12676 9920
rect 12624 9877 12633 9911
rect 12633 9877 12667 9911
rect 12667 9877 12676 9911
rect 12624 9868 12676 9877
rect 13820 9868 13872 9920
rect 14464 9911 14516 9920
rect 14464 9877 14473 9911
rect 14473 9877 14507 9911
rect 14507 9877 14516 9911
rect 14464 9868 14516 9877
rect 14832 9936 14884 9988
rect 14924 9868 14976 9920
rect 15292 9868 15344 9920
rect 15844 9911 15896 9920
rect 15844 9877 15853 9911
rect 15853 9877 15887 9911
rect 15887 9877 15896 9911
rect 15844 9868 15896 9877
rect 17592 9911 17644 9920
rect 17592 9877 17601 9911
rect 17601 9877 17635 9911
rect 17635 9877 17644 9911
rect 17592 9868 17644 9877
rect 18052 9911 18104 9920
rect 18052 9877 18061 9911
rect 18061 9877 18095 9911
rect 18095 9877 18104 9911
rect 18052 9868 18104 9877
rect 20904 9868 20956 9920
rect 22008 10115 22060 10124
rect 22008 10081 22025 10115
rect 22025 10081 22059 10115
rect 22059 10081 22060 10115
rect 22008 10072 22060 10081
rect 21824 10004 21876 10056
rect 22376 10115 22428 10124
rect 22376 10081 22385 10115
rect 22385 10081 22419 10115
rect 22419 10081 22428 10115
rect 22376 10072 22428 10081
rect 22928 10115 22980 10124
rect 22928 10081 22937 10115
rect 22937 10081 22971 10115
rect 22971 10081 22980 10115
rect 22928 10072 22980 10081
rect 22744 9936 22796 9988
rect 22100 9868 22152 9920
rect 22192 9911 22244 9920
rect 22192 9877 22201 9911
rect 22201 9877 22235 9911
rect 22235 9877 22244 9911
rect 22192 9868 22244 9877
rect 4250 9766 4302 9818
rect 4314 9766 4366 9818
rect 4378 9766 4430 9818
rect 4442 9766 4494 9818
rect 4506 9766 4558 9818
rect 11955 9766 12007 9818
rect 12019 9766 12071 9818
rect 12083 9766 12135 9818
rect 12147 9766 12199 9818
rect 12211 9766 12263 9818
rect 19660 9766 19712 9818
rect 19724 9766 19776 9818
rect 19788 9766 19840 9818
rect 19852 9766 19904 9818
rect 19916 9766 19968 9818
rect 27365 9766 27417 9818
rect 27429 9766 27481 9818
rect 27493 9766 27545 9818
rect 27557 9766 27609 9818
rect 27621 9766 27673 9818
rect 8392 9664 8444 9716
rect 8852 9707 8904 9716
rect 8852 9673 8861 9707
rect 8861 9673 8895 9707
rect 8895 9673 8904 9707
rect 8852 9664 8904 9673
rect 14372 9664 14424 9716
rect 15936 9664 15988 9716
rect 16580 9664 16632 9716
rect 18052 9664 18104 9716
rect 20904 9664 20956 9716
rect 31668 9664 31720 9716
rect 9772 9639 9824 9648
rect 9772 9605 9781 9639
rect 9781 9605 9815 9639
rect 9815 9605 9824 9639
rect 9772 9596 9824 9605
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 8484 9392 8536 9444
rect 8852 9460 8904 9512
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 13820 9596 13872 9648
rect 8852 9324 8904 9376
rect 9956 9324 10008 9376
rect 10784 9324 10836 9376
rect 11244 9324 11296 9376
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 14924 9503 14976 9512
rect 14924 9469 14933 9503
rect 14933 9469 14967 9503
rect 14967 9469 14976 9503
rect 14924 9460 14976 9469
rect 13176 9392 13228 9401
rect 17316 9503 17368 9512
rect 17316 9469 17325 9503
rect 17325 9469 17359 9503
rect 17359 9469 17368 9503
rect 17316 9460 17368 9469
rect 18144 9392 18196 9444
rect 18972 9503 19024 9512
rect 18972 9469 18981 9503
rect 18981 9469 19015 9503
rect 19015 9469 19024 9503
rect 18972 9460 19024 9469
rect 19340 9503 19392 9512
rect 19340 9469 19349 9503
rect 19349 9469 19383 9503
rect 19383 9469 19392 9503
rect 19340 9460 19392 9469
rect 20904 9460 20956 9512
rect 19432 9392 19484 9444
rect 13268 9324 13320 9376
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 13912 9324 13964 9376
rect 15844 9324 15896 9376
rect 28264 9460 28316 9512
rect 22284 9435 22336 9444
rect 22284 9401 22318 9435
rect 22318 9401 22336 9435
rect 22284 9392 22336 9401
rect 23388 9367 23440 9376
rect 23388 9333 23397 9367
rect 23397 9333 23431 9367
rect 23431 9333 23440 9367
rect 23388 9324 23440 9333
rect 8102 9222 8154 9274
rect 8166 9222 8218 9274
rect 8230 9222 8282 9274
rect 8294 9222 8346 9274
rect 8358 9222 8410 9274
rect 15807 9222 15859 9274
rect 15871 9222 15923 9274
rect 15935 9222 15987 9274
rect 15999 9222 16051 9274
rect 16063 9222 16115 9274
rect 23512 9222 23564 9274
rect 23576 9222 23628 9274
rect 23640 9222 23692 9274
rect 23704 9222 23756 9274
rect 23768 9222 23820 9274
rect 31217 9222 31269 9274
rect 31281 9222 31333 9274
rect 31345 9222 31397 9274
rect 31409 9222 31461 9274
rect 31473 9222 31525 9274
rect 8484 9120 8536 9172
rect 8852 9163 8904 9172
rect 8852 9129 8861 9163
rect 8861 9129 8895 9163
rect 8895 9129 8904 9163
rect 8852 9120 8904 9129
rect 9220 9120 9272 9172
rect 8024 8984 8076 9036
rect 8392 9027 8444 9036
rect 8392 8993 8401 9027
rect 8401 8993 8435 9027
rect 8435 8993 8444 9027
rect 8392 8984 8444 8993
rect 6736 8891 6788 8900
rect 6736 8857 6745 8891
rect 6745 8857 6779 8891
rect 6779 8857 6788 8891
rect 6736 8848 6788 8857
rect 13176 9120 13228 9172
rect 13636 9120 13688 9172
rect 13268 8984 13320 9036
rect 13912 9052 13964 9104
rect 18328 9120 18380 9172
rect 17316 9052 17368 9104
rect 18972 9120 19024 9172
rect 19432 9120 19484 9172
rect 20076 9120 20128 9172
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 13176 8848 13228 8900
rect 8668 8780 8720 8832
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9404 8780 9456 8789
rect 14004 8823 14056 8832
rect 14004 8789 14013 8823
rect 14013 8789 14047 8823
rect 14047 8789 14056 8823
rect 14004 8780 14056 8789
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 16212 8959 16264 8968
rect 16212 8925 16221 8959
rect 16221 8925 16255 8959
rect 16255 8925 16264 8959
rect 16212 8916 16264 8925
rect 18328 9027 18380 9036
rect 18328 8993 18337 9027
rect 18337 8993 18371 9027
rect 18371 8993 18380 9027
rect 18328 8984 18380 8993
rect 18788 8984 18840 9036
rect 18420 8916 18472 8968
rect 19984 9027 20036 9036
rect 19984 8993 19993 9027
rect 19993 8993 20027 9027
rect 20027 8993 20036 9027
rect 19984 8984 20036 8993
rect 20720 9027 20772 9036
rect 20720 8993 20729 9027
rect 20729 8993 20763 9027
rect 20763 8993 20772 9027
rect 20720 8984 20772 8993
rect 19432 8848 19484 8900
rect 20904 8916 20956 8968
rect 21272 8916 21324 8968
rect 21640 8916 21692 8968
rect 14648 8780 14700 8832
rect 15476 8780 15528 8832
rect 18696 8780 18748 8832
rect 18788 8780 18840 8832
rect 20076 8780 20128 8832
rect 20536 8780 20588 8832
rect 28448 8780 28500 8832
rect 4250 8678 4302 8730
rect 4314 8678 4366 8730
rect 4378 8678 4430 8730
rect 4442 8678 4494 8730
rect 4506 8678 4558 8730
rect 11955 8678 12007 8730
rect 12019 8678 12071 8730
rect 12083 8678 12135 8730
rect 12147 8678 12199 8730
rect 12211 8678 12263 8730
rect 19660 8678 19712 8730
rect 19724 8678 19776 8730
rect 19788 8678 19840 8730
rect 19852 8678 19904 8730
rect 19916 8678 19968 8730
rect 27365 8678 27417 8730
rect 27429 8678 27481 8730
rect 27493 8678 27545 8730
rect 27557 8678 27609 8730
rect 27621 8678 27673 8730
rect 8668 8619 8720 8628
rect 8668 8585 8677 8619
rect 8677 8585 8711 8619
rect 8711 8585 8720 8619
rect 8668 8576 8720 8585
rect 9220 8576 9272 8628
rect 19340 8576 19392 8628
rect 19800 8576 19852 8628
rect 14280 8508 14332 8560
rect 8484 8372 8536 8424
rect 12992 8440 13044 8492
rect 21272 8576 21324 8628
rect 21824 8576 21876 8628
rect 28264 8508 28316 8560
rect 8392 8304 8444 8356
rect 9496 8372 9548 8424
rect 9680 8372 9732 8424
rect 10784 8372 10836 8424
rect 13176 8415 13228 8424
rect 13176 8381 13185 8415
rect 13185 8381 13219 8415
rect 13219 8381 13228 8415
rect 13176 8372 13228 8381
rect 14004 8415 14056 8424
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 14280 8415 14332 8424
rect 14280 8381 14289 8415
rect 14289 8381 14323 8415
rect 14323 8381 14332 8415
rect 14280 8372 14332 8381
rect 14648 8415 14700 8424
rect 14648 8381 14657 8415
rect 14657 8381 14691 8415
rect 14691 8381 14700 8415
rect 14648 8372 14700 8381
rect 19616 8372 19668 8424
rect 13912 8347 13964 8356
rect 13912 8313 13921 8347
rect 13921 8313 13955 8347
rect 13955 8313 13964 8347
rect 13912 8304 13964 8313
rect 17592 8304 17644 8356
rect 19800 8304 19852 8356
rect 8668 8236 8720 8288
rect 9312 8279 9364 8288
rect 9312 8245 9321 8279
rect 9321 8245 9355 8279
rect 9355 8245 9364 8279
rect 9312 8236 9364 8245
rect 11428 8279 11480 8288
rect 11428 8245 11437 8279
rect 11437 8245 11471 8279
rect 11471 8245 11480 8279
rect 11428 8236 11480 8245
rect 13268 8279 13320 8288
rect 13268 8245 13277 8279
rect 13277 8245 13311 8279
rect 13311 8245 13320 8279
rect 13268 8236 13320 8245
rect 13452 8236 13504 8288
rect 14740 8236 14792 8288
rect 16304 8236 16356 8288
rect 19432 8236 19484 8288
rect 19892 8236 19944 8288
rect 21548 8372 21600 8424
rect 23204 8415 23256 8424
rect 23204 8381 23213 8415
rect 23213 8381 23247 8415
rect 23247 8381 23256 8415
rect 23204 8372 23256 8381
rect 20076 8347 20128 8356
rect 20076 8313 20110 8347
rect 20110 8313 20128 8347
rect 20076 8304 20128 8313
rect 20996 8236 21048 8288
rect 23296 8279 23348 8288
rect 23296 8245 23305 8279
rect 23305 8245 23339 8279
rect 23339 8245 23348 8279
rect 23296 8236 23348 8245
rect 8102 8134 8154 8186
rect 8166 8134 8218 8186
rect 8230 8134 8282 8186
rect 8294 8134 8346 8186
rect 8358 8134 8410 8186
rect 15807 8134 15859 8186
rect 15871 8134 15923 8186
rect 15935 8134 15987 8186
rect 15999 8134 16051 8186
rect 16063 8134 16115 8186
rect 23512 8134 23564 8186
rect 23576 8134 23628 8186
rect 23640 8134 23692 8186
rect 23704 8134 23756 8186
rect 23768 8134 23820 8186
rect 31217 8134 31269 8186
rect 31281 8134 31333 8186
rect 31345 8134 31397 8186
rect 31409 8134 31461 8186
rect 31473 8134 31525 8186
rect 8484 8032 8536 8084
rect 13268 8032 13320 8084
rect 13820 8032 13872 8084
rect 9220 7964 9272 8016
rect 9864 7964 9916 8016
rect 17592 8032 17644 8084
rect 19432 8032 19484 8084
rect 19616 8032 19668 8084
rect 19892 8075 19944 8084
rect 19892 8041 19901 8075
rect 19901 8041 19935 8075
rect 19935 8041 19944 8075
rect 19892 8032 19944 8041
rect 20720 8032 20772 8084
rect 20996 8032 21048 8084
rect 7748 7939 7800 7948
rect 7748 7905 7766 7939
rect 7766 7905 7800 7939
rect 7748 7896 7800 7905
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 8576 7896 8628 7948
rect 8760 7896 8812 7948
rect 10324 7896 10376 7948
rect 13452 7896 13504 7948
rect 13912 7896 13964 7948
rect 14004 7896 14056 7948
rect 16212 7964 16264 8016
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 8484 7760 8536 7812
rect 13728 7803 13780 7812
rect 13728 7769 13737 7803
rect 13737 7769 13771 7803
rect 13771 7769 13780 7803
rect 13728 7760 13780 7769
rect 14740 7828 14792 7880
rect 20168 7964 20220 8016
rect 20444 8007 20496 8016
rect 20444 7973 20453 8007
rect 20453 7973 20487 8007
rect 20487 7973 20496 8007
rect 20444 7964 20496 7973
rect 20260 7937 20312 7948
rect 20260 7903 20269 7937
rect 20269 7903 20303 7937
rect 20303 7903 20312 7937
rect 20260 7896 20312 7903
rect 20536 7896 20588 7948
rect 21640 8007 21692 8016
rect 21640 7973 21649 8007
rect 21649 7973 21683 8007
rect 21683 7973 21692 8007
rect 21640 7964 21692 7973
rect 22284 7964 22336 8016
rect 23296 7964 23348 8016
rect 20444 7760 20496 7812
rect 21824 7896 21876 7948
rect 21640 7828 21692 7880
rect 9680 7692 9732 7744
rect 10968 7692 11020 7744
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 14096 7692 14148 7744
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 17040 7692 17092 7744
rect 17500 7735 17552 7744
rect 17500 7701 17509 7735
rect 17509 7701 17543 7735
rect 17543 7701 17552 7735
rect 17500 7692 17552 7701
rect 19984 7692 20036 7744
rect 20076 7692 20128 7744
rect 28264 7692 28316 7744
rect 4250 7590 4302 7642
rect 4314 7590 4366 7642
rect 4378 7590 4430 7642
rect 4442 7590 4494 7642
rect 4506 7590 4558 7642
rect 11955 7590 12007 7642
rect 12019 7590 12071 7642
rect 12083 7590 12135 7642
rect 12147 7590 12199 7642
rect 12211 7590 12263 7642
rect 19660 7590 19712 7642
rect 19724 7590 19776 7642
rect 19788 7590 19840 7642
rect 19852 7590 19904 7642
rect 19916 7590 19968 7642
rect 27365 7590 27417 7642
rect 27429 7590 27481 7642
rect 27493 7590 27545 7642
rect 27557 7590 27609 7642
rect 27621 7590 27673 7642
rect 7748 7488 7800 7540
rect 10324 7531 10376 7540
rect 8760 7420 8812 7472
rect 10324 7497 10333 7531
rect 10333 7497 10367 7531
rect 10367 7497 10376 7531
rect 10324 7488 10376 7497
rect 12900 7488 12952 7540
rect 14740 7488 14792 7540
rect 20168 7488 20220 7540
rect 20536 7488 20588 7540
rect 21640 7531 21692 7540
rect 21640 7497 21649 7531
rect 21649 7497 21683 7531
rect 21683 7497 21692 7531
rect 21640 7488 21692 7497
rect 7748 7352 7800 7404
rect 9220 7420 9272 7472
rect 7656 7327 7708 7336
rect 7656 7293 7665 7327
rect 7665 7293 7699 7327
rect 7699 7293 7708 7327
rect 7656 7284 7708 7293
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 11980 7420 12032 7472
rect 12532 7420 12584 7472
rect 9404 7284 9456 7336
rect 13728 7352 13780 7404
rect 20628 7420 20680 7472
rect 14096 7352 14148 7404
rect 8668 7216 8720 7268
rect 9864 7327 9916 7336
rect 9864 7293 9873 7327
rect 9873 7293 9907 7327
rect 9907 7293 9916 7327
rect 9864 7284 9916 7293
rect 8760 7148 8812 7200
rect 10416 7327 10468 7336
rect 10416 7293 10425 7327
rect 10425 7293 10459 7327
rect 10459 7293 10468 7327
rect 10416 7284 10468 7293
rect 12256 7327 12308 7336
rect 12256 7293 12265 7327
rect 12265 7293 12299 7327
rect 12299 7293 12308 7327
rect 12256 7284 12308 7293
rect 12900 7284 12952 7336
rect 14188 7284 14240 7336
rect 17592 7284 17644 7336
rect 19432 7352 19484 7404
rect 19800 7327 19852 7336
rect 19800 7293 19809 7327
rect 19809 7293 19843 7327
rect 19843 7293 19852 7327
rect 19800 7284 19852 7293
rect 20720 7327 20772 7336
rect 22284 7488 22336 7540
rect 21824 7420 21876 7472
rect 20720 7293 20737 7327
rect 20737 7293 20771 7327
rect 20771 7293 20772 7327
rect 20720 7284 20772 7293
rect 23204 7284 23256 7336
rect 12348 7148 12400 7200
rect 12532 7148 12584 7200
rect 14096 7191 14148 7200
rect 14096 7157 14105 7191
rect 14105 7157 14139 7191
rect 14139 7157 14148 7191
rect 14096 7148 14148 7157
rect 14464 7148 14516 7200
rect 17040 7191 17092 7200
rect 17040 7157 17049 7191
rect 17049 7157 17083 7191
rect 17083 7157 17092 7191
rect 17040 7148 17092 7157
rect 20260 7148 20312 7200
rect 20720 7148 20772 7200
rect 20904 7148 20956 7200
rect 28264 7148 28316 7200
rect 8102 7046 8154 7098
rect 8166 7046 8218 7098
rect 8230 7046 8282 7098
rect 8294 7046 8346 7098
rect 8358 7046 8410 7098
rect 15807 7046 15859 7098
rect 15871 7046 15923 7098
rect 15935 7046 15987 7098
rect 15999 7046 16051 7098
rect 16063 7046 16115 7098
rect 23512 7046 23564 7098
rect 23576 7046 23628 7098
rect 23640 7046 23692 7098
rect 23704 7046 23756 7098
rect 23768 7046 23820 7098
rect 31217 7046 31269 7098
rect 31281 7046 31333 7098
rect 31345 7046 31397 7098
rect 31409 7046 31461 7098
rect 31473 7046 31525 7098
rect 7656 6944 7708 6996
rect 7932 6944 7984 6996
rect 9404 6987 9456 6996
rect 9404 6953 9413 6987
rect 9413 6953 9447 6987
rect 9447 6953 9456 6987
rect 9404 6944 9456 6953
rect 9864 6944 9916 6996
rect 10416 6987 10468 6996
rect 10416 6953 10425 6987
rect 10425 6953 10459 6987
rect 10459 6953 10468 6987
rect 10416 6944 10468 6953
rect 12348 6944 12400 6996
rect 12900 6944 12952 6996
rect 14464 6944 14516 6996
rect 10140 6919 10192 6928
rect 10140 6885 10149 6919
rect 10149 6885 10183 6919
rect 10183 6885 10192 6919
rect 10140 6876 10192 6885
rect 11980 6876 12032 6928
rect 9680 6740 9732 6792
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 12256 6851 12308 6860
rect 12256 6817 12265 6851
rect 12265 6817 12299 6851
rect 12299 6817 12308 6851
rect 12256 6808 12308 6817
rect 14096 6876 14148 6928
rect 19432 6944 19484 6996
rect 19800 6987 19852 6996
rect 19800 6953 19809 6987
rect 19809 6953 19843 6987
rect 19843 6953 19852 6987
rect 19800 6944 19852 6953
rect 17040 6851 17092 6860
rect 17040 6817 17049 6851
rect 17049 6817 17083 6851
rect 17083 6817 17092 6851
rect 17040 6808 17092 6817
rect 10692 6647 10744 6656
rect 10692 6613 10701 6647
rect 10701 6613 10735 6647
rect 10735 6613 10744 6647
rect 10692 6604 10744 6613
rect 11336 6647 11388 6656
rect 11336 6613 11345 6647
rect 11345 6613 11379 6647
rect 11379 6613 11388 6647
rect 11336 6604 11388 6613
rect 11612 6647 11664 6656
rect 11612 6613 11621 6647
rect 11621 6613 11655 6647
rect 11655 6613 11664 6647
rect 11612 6604 11664 6613
rect 14648 6604 14700 6656
rect 15016 6647 15068 6656
rect 15016 6613 15025 6647
rect 15025 6613 15059 6647
rect 15059 6613 15068 6647
rect 15016 6604 15068 6613
rect 18144 6808 18196 6860
rect 18788 6808 18840 6860
rect 18328 6604 18380 6656
rect 19064 6672 19116 6724
rect 19432 6857 19484 6866
rect 19432 6823 19441 6857
rect 19441 6823 19475 6857
rect 19475 6823 19484 6857
rect 19432 6814 19484 6823
rect 19156 6604 19208 6656
rect 20076 6876 20128 6928
rect 20628 6987 20680 6996
rect 20628 6953 20637 6987
rect 20637 6953 20671 6987
rect 20671 6953 20680 6987
rect 20628 6944 20680 6953
rect 20904 6987 20956 6996
rect 20904 6953 20913 6987
rect 20913 6953 20947 6987
rect 20947 6953 20956 6987
rect 20904 6944 20956 6953
rect 21824 6944 21876 6996
rect 20628 6808 20680 6860
rect 21088 6808 21140 6860
rect 28264 6604 28316 6656
rect 4250 6502 4302 6554
rect 4314 6502 4366 6554
rect 4378 6502 4430 6554
rect 4442 6502 4494 6554
rect 4506 6502 4558 6554
rect 11955 6502 12007 6554
rect 12019 6502 12071 6554
rect 12083 6502 12135 6554
rect 12147 6502 12199 6554
rect 12211 6502 12263 6554
rect 19660 6502 19712 6554
rect 19724 6502 19776 6554
rect 19788 6502 19840 6554
rect 19852 6502 19904 6554
rect 19916 6502 19968 6554
rect 27365 6502 27417 6554
rect 27429 6502 27481 6554
rect 27493 6502 27545 6554
rect 27557 6502 27609 6554
rect 27621 6502 27673 6554
rect 10140 6400 10192 6452
rect 10692 6400 10744 6452
rect 9680 6196 9732 6248
rect 10508 6196 10560 6248
rect 11336 6400 11388 6452
rect 14648 6196 14700 6248
rect 17040 6400 17092 6452
rect 18788 6400 18840 6452
rect 20076 6400 20128 6452
rect 17868 6332 17920 6384
rect 17776 6264 17828 6316
rect 18328 6264 18380 6316
rect 12532 6128 12584 6180
rect 16212 6128 16264 6180
rect 9680 6060 9732 6112
rect 13544 6060 13596 6112
rect 16764 6060 16816 6112
rect 17224 6060 17276 6112
rect 18144 6196 18196 6248
rect 21088 6196 21140 6248
rect 19248 6128 19300 6180
rect 20628 6171 20680 6180
rect 20628 6137 20662 6171
rect 20662 6137 20680 6171
rect 20628 6128 20680 6137
rect 18236 6060 18288 6112
rect 20444 6060 20496 6112
rect 21732 6103 21784 6112
rect 21732 6069 21741 6103
rect 21741 6069 21775 6103
rect 21775 6069 21784 6103
rect 21732 6060 21784 6069
rect 8102 5958 8154 6010
rect 8166 5958 8218 6010
rect 8230 5958 8282 6010
rect 8294 5958 8346 6010
rect 8358 5958 8410 6010
rect 15807 5958 15859 6010
rect 15871 5958 15923 6010
rect 15935 5958 15987 6010
rect 15999 5958 16051 6010
rect 16063 5958 16115 6010
rect 23512 5958 23564 6010
rect 23576 5958 23628 6010
rect 23640 5958 23692 6010
rect 23704 5958 23756 6010
rect 23768 5958 23820 6010
rect 31217 5958 31269 6010
rect 31281 5958 31333 6010
rect 31345 5958 31397 6010
rect 31409 5958 31461 6010
rect 31473 5958 31525 6010
rect 11612 5856 11664 5908
rect 16212 5899 16264 5908
rect 16212 5865 16221 5899
rect 16221 5865 16255 5899
rect 16255 5865 16264 5899
rect 16212 5856 16264 5865
rect 17224 5856 17276 5908
rect 17776 5899 17828 5908
rect 17776 5865 17785 5899
rect 17785 5865 17819 5899
rect 17819 5865 17828 5899
rect 17776 5856 17828 5865
rect 18236 5856 18288 5908
rect 14648 5788 14700 5840
rect 10508 5720 10560 5772
rect 16212 5652 16264 5704
rect 16396 5584 16448 5636
rect 17408 5720 17460 5772
rect 18144 5788 18196 5840
rect 17592 5720 17644 5772
rect 17684 5584 17736 5636
rect 17960 5761 18012 5772
rect 17960 5727 17969 5761
rect 17969 5727 18003 5761
rect 18003 5727 18012 5761
rect 17960 5720 18012 5727
rect 18512 5763 18564 5772
rect 18512 5729 18521 5763
rect 18521 5729 18555 5763
rect 18555 5729 18564 5763
rect 18512 5720 18564 5729
rect 19156 5899 19208 5908
rect 19156 5865 19165 5899
rect 19165 5865 19199 5899
rect 19199 5865 19208 5899
rect 19156 5856 19208 5865
rect 19248 5856 19300 5908
rect 18236 5584 18288 5636
rect 12348 5516 12400 5568
rect 14188 5516 14240 5568
rect 17408 5559 17460 5568
rect 17408 5525 17417 5559
rect 17417 5525 17451 5559
rect 17451 5525 17460 5559
rect 17408 5516 17460 5525
rect 4250 5414 4302 5466
rect 4314 5414 4366 5466
rect 4378 5414 4430 5466
rect 4442 5414 4494 5466
rect 4506 5414 4558 5466
rect 11955 5414 12007 5466
rect 12019 5414 12071 5466
rect 12083 5414 12135 5466
rect 12147 5414 12199 5466
rect 12211 5414 12263 5466
rect 19660 5414 19712 5466
rect 19724 5414 19776 5466
rect 19788 5414 19840 5466
rect 19852 5414 19904 5466
rect 19916 5414 19968 5466
rect 27365 5414 27417 5466
rect 27429 5414 27481 5466
rect 27493 5414 27545 5466
rect 27557 5414 27609 5466
rect 27621 5414 27673 5466
rect 16212 5312 16264 5364
rect 16212 5108 16264 5160
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 16488 5040 16540 5092
rect 18512 5108 18564 5160
rect 21272 4972 21324 5024
rect 8102 4870 8154 4922
rect 8166 4870 8218 4922
rect 8230 4870 8282 4922
rect 8294 4870 8346 4922
rect 8358 4870 8410 4922
rect 15807 4870 15859 4922
rect 15871 4870 15923 4922
rect 15935 4870 15987 4922
rect 15999 4870 16051 4922
rect 16063 4870 16115 4922
rect 23512 4870 23564 4922
rect 23576 4870 23628 4922
rect 23640 4870 23692 4922
rect 23704 4870 23756 4922
rect 23768 4870 23820 4922
rect 31217 4870 31269 4922
rect 31281 4870 31333 4922
rect 31345 4870 31397 4922
rect 31409 4870 31461 4922
rect 31473 4870 31525 4922
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 16488 4768 16540 4820
rect 4250 4326 4302 4378
rect 4314 4326 4366 4378
rect 4378 4326 4430 4378
rect 4442 4326 4494 4378
rect 4506 4326 4558 4378
rect 11955 4326 12007 4378
rect 12019 4326 12071 4378
rect 12083 4326 12135 4378
rect 12147 4326 12199 4378
rect 12211 4326 12263 4378
rect 19660 4326 19712 4378
rect 19724 4326 19776 4378
rect 19788 4326 19840 4378
rect 19852 4326 19904 4378
rect 19916 4326 19968 4378
rect 27365 4326 27417 4378
rect 27429 4326 27481 4378
rect 27493 4326 27545 4378
rect 27557 4326 27609 4378
rect 27621 4326 27673 4378
rect 10324 4088 10376 4140
rect 11244 4088 11296 4140
rect 8102 3782 8154 3834
rect 8166 3782 8218 3834
rect 8230 3782 8282 3834
rect 8294 3782 8346 3834
rect 8358 3782 8410 3834
rect 15807 3782 15859 3834
rect 15871 3782 15923 3834
rect 15935 3782 15987 3834
rect 15999 3782 16051 3834
rect 16063 3782 16115 3834
rect 23512 3782 23564 3834
rect 23576 3782 23628 3834
rect 23640 3782 23692 3834
rect 23704 3782 23756 3834
rect 23768 3782 23820 3834
rect 31217 3782 31269 3834
rect 31281 3782 31333 3834
rect 31345 3782 31397 3834
rect 31409 3782 31461 3834
rect 31473 3782 31525 3834
rect 9036 3408 9088 3460
rect 12624 3408 12676 3460
rect 4250 3238 4302 3290
rect 4314 3238 4366 3290
rect 4378 3238 4430 3290
rect 4442 3238 4494 3290
rect 4506 3238 4558 3290
rect 11955 3238 12007 3290
rect 12019 3238 12071 3290
rect 12083 3238 12135 3290
rect 12147 3238 12199 3290
rect 12211 3238 12263 3290
rect 19660 3238 19712 3290
rect 19724 3238 19776 3290
rect 19788 3238 19840 3290
rect 19852 3238 19904 3290
rect 19916 3238 19968 3290
rect 27365 3238 27417 3290
rect 27429 3238 27481 3290
rect 27493 3238 27545 3290
rect 27557 3238 27609 3290
rect 27621 3238 27673 3290
rect 8102 2694 8154 2746
rect 8166 2694 8218 2746
rect 8230 2694 8282 2746
rect 8294 2694 8346 2746
rect 8358 2694 8410 2746
rect 15807 2694 15859 2746
rect 15871 2694 15923 2746
rect 15935 2694 15987 2746
rect 15999 2694 16051 2746
rect 16063 2694 16115 2746
rect 23512 2694 23564 2746
rect 23576 2694 23628 2746
rect 23640 2694 23692 2746
rect 23704 2694 23756 2746
rect 23768 2694 23820 2746
rect 31217 2694 31269 2746
rect 31281 2694 31333 2746
rect 31345 2694 31397 2746
rect 31409 2694 31461 2746
rect 31473 2694 31525 2746
rect 4250 2150 4302 2202
rect 4314 2150 4366 2202
rect 4378 2150 4430 2202
rect 4442 2150 4494 2202
rect 4506 2150 4558 2202
rect 11955 2150 12007 2202
rect 12019 2150 12071 2202
rect 12083 2150 12135 2202
rect 12147 2150 12199 2202
rect 12211 2150 12263 2202
rect 19660 2150 19712 2202
rect 19724 2150 19776 2202
rect 19788 2150 19840 2202
rect 19852 2150 19904 2202
rect 19916 2150 19968 2202
rect 27365 2150 27417 2202
rect 27429 2150 27481 2202
rect 27493 2150 27545 2202
rect 27557 2150 27609 2202
rect 27621 2150 27673 2202
rect 8102 1606 8154 1658
rect 8166 1606 8218 1658
rect 8230 1606 8282 1658
rect 8294 1606 8346 1658
rect 8358 1606 8410 1658
rect 15807 1606 15859 1658
rect 15871 1606 15923 1658
rect 15935 1606 15987 1658
rect 15999 1606 16051 1658
rect 16063 1606 16115 1658
rect 23512 1606 23564 1658
rect 23576 1606 23628 1658
rect 23640 1606 23692 1658
rect 23704 1606 23756 1658
rect 23768 1606 23820 1658
rect 31217 1606 31269 1658
rect 31281 1606 31333 1658
rect 31345 1606 31397 1658
rect 31409 1606 31461 1658
rect 31473 1606 31525 1658
rect 4250 1062 4302 1114
rect 4314 1062 4366 1114
rect 4378 1062 4430 1114
rect 4442 1062 4494 1114
rect 4506 1062 4558 1114
rect 11955 1062 12007 1114
rect 12019 1062 12071 1114
rect 12083 1062 12135 1114
rect 12147 1062 12199 1114
rect 12211 1062 12263 1114
rect 19660 1062 19712 1114
rect 19724 1062 19776 1114
rect 19788 1062 19840 1114
rect 19852 1062 19904 1114
rect 19916 1062 19968 1114
rect 27365 1062 27417 1114
rect 27429 1062 27481 1114
rect 27493 1062 27545 1114
rect 27557 1062 27609 1114
rect 27621 1062 27673 1114
rect 16212 824 16264 876
rect 22652 799 22704 808
rect 22652 765 22661 799
rect 22661 765 22695 799
rect 22695 765 22704 799
rect 22652 756 22704 765
rect 8102 518 8154 570
rect 8166 518 8218 570
rect 8230 518 8282 570
rect 8294 518 8346 570
rect 8358 518 8410 570
rect 15807 518 15859 570
rect 15871 518 15923 570
rect 15935 518 15987 570
rect 15999 518 16051 570
rect 16063 518 16115 570
rect 23512 518 23564 570
rect 23576 518 23628 570
rect 23640 518 23692 570
rect 23704 518 23756 570
rect 23768 518 23820 570
rect 31217 518 31269 570
rect 31281 518 31333 570
rect 31345 518 31397 570
rect 31409 518 31461 570
rect 31473 518 31525 570
rect 16028 416 16080 468
rect 16304 416 16356 468
<< metal2 >>
rect 10966 19600 11022 20000
rect 11610 19600 11666 20000
rect 12254 19600 12310 20000
rect 12898 19600 12954 20000
rect 13542 19600 13598 20000
rect 14186 19600 14242 20000
rect 14830 19600 14886 20000
rect 15474 19600 15530 20000
rect 16118 19600 16174 20000
rect 16762 19600 16818 20000
rect 17406 19600 17462 20000
rect 18050 19600 18106 20000
rect 18694 19600 18750 20000
rect 19338 19600 19394 20000
rect 19982 19600 20038 20000
rect 20626 19600 20682 20000
rect 21270 19600 21326 20000
rect 21914 19600 21970 20000
rect 8102 19068 8410 19077
rect 8102 19066 8108 19068
rect 8164 19066 8188 19068
rect 8244 19066 8268 19068
rect 8324 19066 8348 19068
rect 8404 19066 8410 19068
rect 8164 19014 8166 19066
rect 8346 19014 8348 19066
rect 8102 19012 8108 19014
rect 8164 19012 8188 19014
rect 8244 19012 8268 19014
rect 8324 19012 8348 19014
rect 8404 19012 8410 19014
rect 8102 19003 8410 19012
rect 4250 18524 4558 18533
rect 4250 18522 4256 18524
rect 4312 18522 4336 18524
rect 4392 18522 4416 18524
rect 4472 18522 4496 18524
rect 4552 18522 4558 18524
rect 4312 18470 4314 18522
rect 4494 18470 4496 18522
rect 4250 18468 4256 18470
rect 4312 18468 4336 18470
rect 4392 18468 4416 18470
rect 4472 18468 4496 18470
rect 4552 18468 4558 18470
rect 4250 18459 4558 18468
rect 8102 17980 8410 17989
rect 8102 17978 8108 17980
rect 8164 17978 8188 17980
rect 8244 17978 8268 17980
rect 8324 17978 8348 17980
rect 8404 17978 8410 17980
rect 8164 17926 8166 17978
rect 8346 17926 8348 17978
rect 8102 17924 8108 17926
rect 8164 17924 8188 17926
rect 8244 17924 8268 17926
rect 8324 17924 8348 17926
rect 8404 17924 8410 17926
rect 8102 17915 8410 17924
rect 4250 17436 4558 17445
rect 4250 17434 4256 17436
rect 4312 17434 4336 17436
rect 4392 17434 4416 17436
rect 4472 17434 4496 17436
rect 4552 17434 4558 17436
rect 4312 17382 4314 17434
rect 4494 17382 4496 17434
rect 4250 17380 4256 17382
rect 4312 17380 4336 17382
rect 4392 17380 4416 17382
rect 4472 17380 4496 17382
rect 4552 17380 4558 17382
rect 4250 17371 4558 17380
rect 8102 16892 8410 16901
rect 8102 16890 8108 16892
rect 8164 16890 8188 16892
rect 8244 16890 8268 16892
rect 8324 16890 8348 16892
rect 8404 16890 8410 16892
rect 8164 16838 8166 16890
rect 8346 16838 8348 16890
rect 8102 16836 8108 16838
rect 8164 16836 8188 16838
rect 8244 16836 8268 16838
rect 8324 16836 8348 16838
rect 8404 16836 8410 16838
rect 8102 16827 8410 16836
rect 10980 16574 11008 19600
rect 10796 16546 11008 16574
rect 4250 16348 4558 16357
rect 4250 16346 4256 16348
rect 4312 16346 4336 16348
rect 4392 16346 4416 16348
rect 4472 16346 4496 16348
rect 4552 16346 4558 16348
rect 4312 16294 4314 16346
rect 4494 16294 4496 16346
rect 4250 16292 4256 16294
rect 4312 16292 4336 16294
rect 4392 16292 4416 16294
rect 4472 16292 4496 16294
rect 4552 16292 4558 16294
rect 4250 16283 4558 16292
rect 8102 15804 8410 15813
rect 8102 15802 8108 15804
rect 8164 15802 8188 15804
rect 8244 15802 8268 15804
rect 8324 15802 8348 15804
rect 8404 15802 8410 15804
rect 8164 15750 8166 15802
rect 8346 15750 8348 15802
rect 8102 15748 8108 15750
rect 8164 15748 8188 15750
rect 8244 15748 8268 15750
rect 8324 15748 8348 15750
rect 8404 15748 8410 15750
rect 8102 15739 8410 15748
rect 4250 15260 4558 15269
rect 4250 15258 4256 15260
rect 4312 15258 4336 15260
rect 4392 15258 4416 15260
rect 4472 15258 4496 15260
rect 4552 15258 4558 15260
rect 4312 15206 4314 15258
rect 4494 15206 4496 15258
rect 4250 15204 4256 15206
rect 4312 15204 4336 15206
rect 4392 15204 4416 15206
rect 4472 15204 4496 15206
rect 4552 15204 4558 15206
rect 4250 15195 4558 15204
rect 8102 14716 8410 14725
rect 8102 14714 8108 14716
rect 8164 14714 8188 14716
rect 8244 14714 8268 14716
rect 8324 14714 8348 14716
rect 8404 14714 8410 14716
rect 8164 14662 8166 14714
rect 8346 14662 8348 14714
rect 8102 14660 8108 14662
rect 8164 14660 8188 14662
rect 8244 14660 8268 14662
rect 8324 14660 8348 14662
rect 8404 14660 8410 14662
rect 8102 14651 8410 14660
rect 4250 14172 4558 14181
rect 4250 14170 4256 14172
rect 4312 14170 4336 14172
rect 4392 14170 4416 14172
rect 4472 14170 4496 14172
rect 4552 14170 4558 14172
rect 4312 14118 4314 14170
rect 4494 14118 4496 14170
rect 4250 14116 4256 14118
rect 4312 14116 4336 14118
rect 4392 14116 4416 14118
rect 4472 14116 4496 14118
rect 4552 14116 4558 14118
rect 4250 14107 4558 14116
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 8102 13628 8410 13637
rect 8102 13626 8108 13628
rect 8164 13626 8188 13628
rect 8244 13626 8268 13628
rect 8324 13626 8348 13628
rect 8404 13626 8410 13628
rect 8164 13574 8166 13626
rect 8346 13574 8348 13626
rect 8102 13572 8108 13574
rect 8164 13572 8188 13574
rect 8244 13572 8268 13574
rect 8324 13572 8348 13574
rect 8404 13572 8410 13574
rect 8102 13563 8410 13572
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 4250 13084 4558 13093
rect 4250 13082 4256 13084
rect 4312 13082 4336 13084
rect 4392 13082 4416 13084
rect 4472 13082 4496 13084
rect 4552 13082 4558 13084
rect 4312 13030 4314 13082
rect 4494 13030 4496 13082
rect 4250 13028 4256 13030
rect 4312 13028 4336 13030
rect 4392 13028 4416 13030
rect 4472 13028 4496 13030
rect 4552 13028 4558 13030
rect 4250 13019 4558 13028
rect 8102 12540 8410 12549
rect 8102 12538 8108 12540
rect 8164 12538 8188 12540
rect 8244 12538 8268 12540
rect 8324 12538 8348 12540
rect 8404 12538 8410 12540
rect 8164 12486 8166 12538
rect 8346 12486 8348 12538
rect 8102 12484 8108 12486
rect 8164 12484 8188 12486
rect 8244 12484 8268 12486
rect 8324 12484 8348 12486
rect 8404 12484 8410 12486
rect 8102 12475 8410 12484
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6932 12345 6960 12378
rect 6918 12336 6974 12345
rect 10152 12306 10180 13126
rect 10704 12646 10732 13670
rect 10796 12986 10824 16546
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 13462 11192 13670
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12986 11100 13126
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11164 12782 11192 13398
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 6918 12271 6974 12280
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 4250 11996 4558 12005
rect 4250 11994 4256 11996
rect 4312 11994 4336 11996
rect 4392 11994 4416 11996
rect 4472 11994 4496 11996
rect 4552 11994 4558 11996
rect 4312 11942 4314 11994
rect 4494 11942 4496 11994
rect 4250 11940 4256 11942
rect 4312 11940 4336 11942
rect 4392 11940 4416 11942
rect 4472 11940 4496 11942
rect 4552 11940 4558 11942
rect 4250 11931 4558 11940
rect 9036 11688 9088 11694
rect 6918 11656 6974 11665
rect 9036 11630 9088 11636
rect 6918 11591 6974 11600
rect 6932 11354 6960 11591
rect 8102 11452 8410 11461
rect 8102 11450 8108 11452
rect 8164 11450 8188 11452
rect 8244 11450 8268 11452
rect 8324 11450 8348 11452
rect 8404 11450 8410 11452
rect 8164 11398 8166 11450
rect 8346 11398 8348 11450
rect 8102 11396 8108 11398
rect 8164 11396 8188 11398
rect 8244 11396 8268 11398
rect 8324 11396 8348 11398
rect 8404 11396 8410 11398
rect 8102 11387 8410 11396
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 9048 11286 9076 11630
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9140 11354 9168 11562
rect 9692 11558 9720 12242
rect 10152 11898 10180 12242
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 11354 9720 11494
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 4250 10908 4558 10917
rect 4250 10906 4256 10908
rect 4312 10906 4336 10908
rect 4392 10906 4416 10908
rect 4472 10906 4496 10908
rect 4552 10906 4558 10908
rect 4312 10854 4314 10906
rect 4494 10854 4496 10906
rect 4250 10852 4256 10854
rect 4312 10852 4336 10854
rect 4392 10852 4416 10854
rect 4472 10852 4496 10854
rect 4552 10852 4558 10854
rect 4250 10843 4558 10852
rect 9048 10674 9076 11222
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10742 9720 11018
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8102 10364 8410 10373
rect 8102 10362 8108 10364
rect 8164 10362 8188 10364
rect 8244 10362 8268 10364
rect 8324 10362 8348 10364
rect 8404 10362 8410 10364
rect 8164 10310 8166 10362
rect 8346 10310 8348 10362
rect 8102 10308 8108 10310
rect 8164 10308 8188 10310
rect 8244 10308 8268 10310
rect 8324 10308 8348 10310
rect 8404 10308 8410 10310
rect 7102 10296 7158 10305
rect 8102 10299 8410 10308
rect 7102 10231 7104 10240
rect 7156 10231 7158 10240
rect 7104 10202 7156 10208
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 4250 9820 4558 9829
rect 4250 9818 4256 9820
rect 4312 9818 4336 9820
rect 4392 9818 4416 9820
rect 4472 9818 4496 9820
rect 4552 9818 4558 9820
rect 4312 9766 4314 9818
rect 4494 9766 4496 9818
rect 4250 9764 4256 9766
rect 4312 9764 4336 9766
rect 4392 9764 4416 9766
rect 4472 9764 4496 9766
rect 4552 9764 4558 9766
rect 4250 9755 4558 9764
rect 6734 8936 6790 8945
rect 6734 8871 6736 8880
rect 6788 8871 6790 8880
rect 6736 8842 6788 8848
rect 4250 8732 4558 8741
rect 4250 8730 4256 8732
rect 4312 8730 4336 8732
rect 4392 8730 4416 8732
rect 4472 8730 4496 8732
rect 4552 8730 4558 8732
rect 4312 8678 4314 8730
rect 4494 8678 4496 8730
rect 4250 8676 4256 8678
rect 4312 8676 4336 8678
rect 4392 8676 4416 8678
rect 4472 8676 4496 8678
rect 4552 8676 4558 8678
rect 4250 8667 4558 8676
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 4250 7644 4558 7653
rect 4250 7642 4256 7644
rect 4312 7642 4336 7644
rect 4392 7642 4416 7644
rect 4472 7642 4496 7644
rect 4552 7642 4558 7644
rect 4312 7590 4314 7642
rect 4494 7590 4496 7642
rect 4250 7588 4256 7590
rect 4312 7588 4336 7590
rect 4392 7588 4416 7590
rect 4472 7588 4496 7590
rect 4552 7588 4558 7590
rect 4250 7579 4558 7588
rect 6656 6905 6684 7686
rect 6642 6896 6698 6905
rect 6642 6831 6698 6840
rect 4250 6556 4558 6565
rect 4250 6554 4256 6556
rect 4312 6554 4336 6556
rect 4392 6554 4416 6556
rect 4472 6554 4496 6556
rect 4552 6554 4558 6556
rect 4312 6502 4314 6554
rect 4494 6502 4496 6554
rect 4250 6500 4256 6502
rect 4312 6500 4336 6502
rect 4392 6500 4416 6502
rect 4472 6500 4496 6502
rect 4552 6500 4558 6502
rect 4250 6491 4558 6500
rect 4250 5468 4558 5477
rect 4250 5466 4256 5468
rect 4312 5466 4336 5468
rect 4392 5466 4416 5468
rect 4472 5466 4496 5468
rect 4552 5466 4558 5468
rect 4312 5414 4314 5466
rect 4494 5414 4496 5466
rect 4250 5412 4256 5414
rect 4312 5412 4336 5414
rect 4392 5412 4416 5414
rect 4472 5412 4496 5414
rect 4552 5412 4558 5414
rect 4250 5403 4558 5412
rect 4250 4380 4558 4389
rect 4250 4378 4256 4380
rect 4312 4378 4336 4380
rect 4392 4378 4416 4380
rect 4472 4378 4496 4380
rect 4552 4378 4558 4380
rect 4312 4326 4314 4378
rect 4494 4326 4496 4378
rect 4250 4324 4256 4326
rect 4312 4324 4336 4326
rect 4392 4324 4416 4326
rect 4472 4324 4496 4326
rect 4552 4324 4558 4326
rect 4250 4315 4558 4324
rect 4250 3292 4558 3301
rect 4250 3290 4256 3292
rect 4312 3290 4336 3292
rect 4392 3290 4416 3292
rect 4472 3290 4496 3292
rect 4552 3290 4558 3292
rect 4312 3238 4314 3290
rect 4494 3238 4496 3290
rect 4250 3236 4256 3238
rect 4312 3236 4336 3238
rect 4392 3236 4416 3238
rect 4472 3236 4496 3238
rect 4552 3236 4558 3238
rect 4250 3227 4558 3236
rect 7208 2774 7236 9862
rect 8404 9722 8432 10066
rect 8864 9722 8892 10066
rect 9048 10062 9076 10406
rect 9600 10198 9628 10542
rect 9692 10266 9720 10678
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9784 10266 9812 10542
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 9772 9648 9824 9654
rect 9770 9616 9772 9625
rect 9824 9616 9826 9625
rect 9770 9551 9826 9560
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8102 9276 8410 9285
rect 8102 9274 8108 9276
rect 8164 9274 8188 9276
rect 8244 9274 8268 9276
rect 8324 9274 8348 9276
rect 8404 9274 8410 9276
rect 8164 9222 8166 9274
rect 8346 9222 8348 9274
rect 8102 9220 8108 9222
rect 8164 9220 8188 9222
rect 8244 9220 8268 9222
rect 8324 9220 8348 9222
rect 8404 9220 8410 9222
rect 8102 9211 8410 9220
rect 8496 9178 8524 9386
rect 8864 9382 8892 9454
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8864 9178 8892 9318
rect 9232 9178 9260 9454
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7760 7546 7788 7890
rect 8036 7886 8064 8978
rect 8404 8362 8432 8978
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8634 8708 8774
rect 9232 8634 9260 9114
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8102 8188 8410 8197
rect 8102 8186 8108 8188
rect 8164 8186 8188 8188
rect 8244 8186 8268 8188
rect 8324 8186 8348 8188
rect 8404 8186 8410 8188
rect 8164 8134 8166 8186
rect 8346 8134 8348 8186
rect 8102 8132 8108 8134
rect 8164 8132 8188 8134
rect 8244 8132 8268 8134
rect 8324 8132 8348 8134
rect 8404 8132 8410 8134
rect 8102 8123 8410 8132
rect 8496 8090 8524 8366
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8496 7818 8524 8026
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7760 7410 7788 7482
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 8588 7342 8616 7890
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 7668 7002 7696 7278
rect 7944 7002 7972 7278
rect 8680 7274 8708 8230
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8772 7478 8800 7890
rect 9232 7478 9260 7958
rect 9324 7857 9352 8230
rect 9416 7993 9444 8774
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9402 7984 9458 7993
rect 9402 7919 9458 7928
rect 9310 7848 9366 7857
rect 9310 7783 9366 7792
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8772 7206 8800 7414
rect 9508 7410 9536 8366
rect 9692 7750 9720 8366
rect 9876 8022 9904 11562
rect 10520 11558 10548 12174
rect 10704 12102 10732 12582
rect 11256 12442 11284 13194
rect 11348 12782 11376 13806
rect 11440 13530 11468 13806
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11440 13002 11468 13466
rect 11440 12986 11560 13002
rect 11440 12980 11572 12986
rect 11440 12974 11520 12980
rect 11520 12922 11572 12928
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11762 10732 12038
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10152 10810 10180 11154
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10520 10674 10548 11494
rect 10980 11354 11008 12242
rect 11348 11558 11376 12718
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11440 11898 11468 12242
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11624 11354 11652 19600
rect 12268 18714 12296 19600
rect 12268 18686 12388 18714
rect 11955 18524 12263 18533
rect 11955 18522 11961 18524
rect 12017 18522 12041 18524
rect 12097 18522 12121 18524
rect 12177 18522 12201 18524
rect 12257 18522 12263 18524
rect 12017 18470 12019 18522
rect 12199 18470 12201 18522
rect 11955 18468 11961 18470
rect 12017 18468 12041 18470
rect 12097 18468 12121 18470
rect 12177 18468 12201 18470
rect 12257 18468 12263 18470
rect 11955 18459 12263 18468
rect 11955 17436 12263 17445
rect 11955 17434 11961 17436
rect 12017 17434 12041 17436
rect 12097 17434 12121 17436
rect 12177 17434 12201 17436
rect 12257 17434 12263 17436
rect 12017 17382 12019 17434
rect 12199 17382 12201 17434
rect 11955 17380 11961 17382
rect 12017 17380 12041 17382
rect 12097 17380 12121 17382
rect 12177 17380 12201 17382
rect 12257 17380 12263 17382
rect 11955 17371 12263 17380
rect 11955 16348 12263 16357
rect 11955 16346 11961 16348
rect 12017 16346 12041 16348
rect 12097 16346 12121 16348
rect 12177 16346 12201 16348
rect 12257 16346 12263 16348
rect 12017 16294 12019 16346
rect 12199 16294 12201 16346
rect 11955 16292 11961 16294
rect 12017 16292 12041 16294
rect 12097 16292 12121 16294
rect 12177 16292 12201 16294
rect 12257 16292 12263 16294
rect 11955 16283 12263 16292
rect 11955 15260 12263 15269
rect 11955 15258 11961 15260
rect 12017 15258 12041 15260
rect 12097 15258 12121 15260
rect 12177 15258 12201 15260
rect 12257 15258 12263 15260
rect 12017 15206 12019 15258
rect 12199 15206 12201 15258
rect 11955 15204 11961 15206
rect 12017 15204 12041 15206
rect 12097 15204 12121 15206
rect 12177 15204 12201 15206
rect 12257 15204 12263 15206
rect 11955 15195 12263 15204
rect 11955 14172 12263 14181
rect 11955 14170 11961 14172
rect 12017 14170 12041 14172
rect 12097 14170 12121 14172
rect 12177 14170 12201 14172
rect 12257 14170 12263 14172
rect 12017 14118 12019 14170
rect 12199 14118 12201 14170
rect 11955 14116 11961 14118
rect 12017 14116 12041 14118
rect 12097 14116 12121 14118
rect 12177 14116 12201 14118
rect 12257 14116 12263 14118
rect 11955 14107 12263 14116
rect 12360 14090 12388 18686
rect 12360 14074 12480 14090
rect 12360 14068 12492 14074
rect 12360 14062 12440 14068
rect 12440 14010 12492 14016
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11808 12850 11836 13126
rect 11955 13084 12263 13093
rect 11955 13082 11961 13084
rect 12017 13082 12041 13084
rect 12097 13082 12121 13084
rect 12177 13082 12201 13084
rect 12257 13082 12263 13084
rect 12017 13030 12019 13082
rect 12199 13030 12201 13082
rect 11955 13028 11961 13030
rect 12017 13028 12041 13030
rect 12097 13028 12121 13030
rect 12177 13028 12201 13030
rect 12257 13028 12263 13030
rect 11955 13019 12263 13028
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11808 12442 11836 12786
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11900 12374 11928 12718
rect 12912 12442 12940 19600
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13188 13938 13216 14418
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13188 13462 13216 13874
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13464 13530 13492 13806
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12268 12084 12296 12242
rect 12440 12096 12492 12102
rect 12268 12056 12388 12084
rect 11955 11996 12263 12005
rect 11955 11994 11961 11996
rect 12017 11994 12041 11996
rect 12097 11994 12121 11996
rect 12177 11994 12201 11996
rect 12257 11994 12263 11996
rect 12017 11942 12019 11994
rect 12199 11942 12201 11994
rect 11955 11940 11961 11942
rect 12017 11940 12041 11942
rect 12097 11940 12121 11942
rect 12177 11940 12201 11942
rect 12257 11940 12263 11942
rect 11955 11931 12263 11940
rect 12360 11898 12388 12056
rect 12440 12038 12492 12044
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12452 11830 12480 12038
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11808 11286 11836 11494
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 12912 11218 12940 11494
rect 13556 11354 13584 19600
rect 14200 14618 14228 19600
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14016 13530 14044 13670
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14016 13190 14044 13330
rect 14384 13258 14412 13670
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 12646 14044 13126
rect 14476 12850 14504 14418
rect 14752 14074 14780 14418
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14752 13530 14780 14010
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14016 12306 14044 12582
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 14108 11694 14136 12310
rect 14476 12306 14504 12786
rect 14844 12442 14872 19600
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 15488 11898 15516 19600
rect 16132 19258 16160 19600
rect 16132 19230 16252 19258
rect 15807 19068 16115 19077
rect 15807 19066 15813 19068
rect 15869 19066 15893 19068
rect 15949 19066 15973 19068
rect 16029 19066 16053 19068
rect 16109 19066 16115 19068
rect 15869 19014 15871 19066
rect 16051 19014 16053 19066
rect 15807 19012 15813 19014
rect 15869 19012 15893 19014
rect 15949 19012 15973 19014
rect 16029 19012 16053 19014
rect 16109 19012 16115 19014
rect 15807 19003 16115 19012
rect 15807 17980 16115 17989
rect 15807 17978 15813 17980
rect 15869 17978 15893 17980
rect 15949 17978 15973 17980
rect 16029 17978 16053 17980
rect 16109 17978 16115 17980
rect 15869 17926 15871 17978
rect 16051 17926 16053 17978
rect 15807 17924 15813 17926
rect 15869 17924 15893 17926
rect 15949 17924 15973 17926
rect 16029 17924 16053 17926
rect 16109 17924 16115 17926
rect 15807 17915 16115 17924
rect 15807 16892 16115 16901
rect 15807 16890 15813 16892
rect 15869 16890 15893 16892
rect 15949 16890 15973 16892
rect 16029 16890 16053 16892
rect 16109 16890 16115 16892
rect 15869 16838 15871 16890
rect 16051 16838 16053 16890
rect 15807 16836 15813 16838
rect 15869 16836 15893 16838
rect 15949 16836 15973 16838
rect 16029 16836 16053 16838
rect 16109 16836 16115 16838
rect 15807 16827 16115 16836
rect 15807 15804 16115 15813
rect 15807 15802 15813 15804
rect 15869 15802 15893 15804
rect 15949 15802 15973 15804
rect 16029 15802 16053 15804
rect 16109 15802 16115 15804
rect 15869 15750 15871 15802
rect 16051 15750 16053 15802
rect 15807 15748 15813 15750
rect 15869 15748 15893 15750
rect 15949 15748 15973 15750
rect 16029 15748 16053 15750
rect 16109 15748 16115 15750
rect 15807 15739 16115 15748
rect 15807 14716 16115 14725
rect 15807 14714 15813 14716
rect 15869 14714 15893 14716
rect 15949 14714 15973 14716
rect 16029 14714 16053 14716
rect 16109 14714 16115 14716
rect 15869 14662 15871 14714
rect 16051 14662 16053 14714
rect 15807 14660 15813 14662
rect 15869 14660 15893 14662
rect 15949 14660 15973 14662
rect 16029 14660 16053 14662
rect 16109 14660 16115 14662
rect 15807 14651 16115 14660
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 13326 15700 13670
rect 15807 13628 16115 13637
rect 15807 13626 15813 13628
rect 15869 13626 15893 13628
rect 15949 13626 15973 13628
rect 16029 13626 16053 13628
rect 16109 13626 16115 13628
rect 15869 13574 15871 13626
rect 16051 13574 16053 13626
rect 15807 13572 15813 13574
rect 15869 13572 15893 13574
rect 15949 13572 15973 13574
rect 16029 13572 16053 13574
rect 16109 13572 16115 13574
rect 15807 13563 16115 13572
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15580 12306 15608 13262
rect 15672 12442 15700 13262
rect 15807 12540 16115 12549
rect 15807 12538 15813 12540
rect 15869 12538 15893 12540
rect 15949 12538 15973 12540
rect 16029 12538 16053 12540
rect 16109 12538 16115 12540
rect 15869 12486 15871 12538
rect 16051 12486 16053 12538
rect 15807 12484 15813 12486
rect 15869 12484 15893 12486
rect 15949 12484 15973 12486
rect 16029 12484 16053 12486
rect 16109 12484 16115 12486
rect 15807 12475 16115 12484
rect 15660 12436 15712 12442
rect 16224 12434 16252 19230
rect 16776 14618 16804 19600
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16500 13530 16528 13738
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 15660 12378 15712 12384
rect 16132 12406 16252 12434
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 16132 11642 16160 12406
rect 16212 12300 16264 12306
rect 16316 12288 16344 13330
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 16500 12306 16528 12650
rect 16776 12646 16804 13126
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16776 12442 16804 12582
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16264 12260 16344 12288
rect 16488 12300 16540 12306
rect 16212 12242 16264 12248
rect 16488 12242 16540 12248
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 14108 11218 14136 11630
rect 16132 11614 16252 11642
rect 15807 11452 16115 11461
rect 15807 11450 15813 11452
rect 15869 11450 15893 11452
rect 15949 11450 15973 11452
rect 16029 11450 16053 11452
rect 16109 11450 16115 11452
rect 15869 11398 15871 11450
rect 16051 11398 16053 11450
rect 15807 11396 15813 11398
rect 15869 11396 15893 11398
rect 15949 11396 15973 11398
rect 16029 11396 16053 11398
rect 16109 11396 16115 11398
rect 15807 11387 16115 11396
rect 16224 11354 16252 11614
rect 17420 11354 17448 19600
rect 18064 14074 18092 19600
rect 18708 14634 18736 19600
rect 18524 14606 18736 14634
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17776 13864 17828 13870
rect 17960 13864 18012 13870
rect 17776 13806 17828 13812
rect 17880 13812 17960 13818
rect 17880 13806 18012 13812
rect 17788 13530 17816 13806
rect 17880 13790 18000 13806
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17880 13394 17908 13790
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 18524 12986 18552 14606
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18616 13870 18644 14418
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18616 12986 18644 13806
rect 18708 13462 18736 13806
rect 18696 13456 18748 13462
rect 18696 13398 18748 13404
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18708 12918 18736 13398
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18708 12442 18736 12854
rect 18984 12782 19012 13806
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10796 10674 10824 11086
rect 10980 10810 11008 11154
rect 14108 11098 14136 11154
rect 14108 11070 14228 11098
rect 11955 10908 12263 10917
rect 11955 10906 11961 10908
rect 12017 10906 12041 10908
rect 12097 10906 12121 10908
rect 12177 10906 12201 10908
rect 12257 10906 12263 10908
rect 12017 10854 12019 10906
rect 12199 10854 12201 10906
rect 11955 10852 11961 10854
rect 12017 10852 12041 10854
rect 12097 10852 12121 10854
rect 12177 10852 12201 10854
rect 12257 10852 12263 10854
rect 11150 10840 11206 10849
rect 11955 10843 12263 10852
rect 10968 10804 11020 10810
rect 11150 10775 11152 10784
rect 10968 10746 11020 10752
rect 11204 10775 11206 10784
rect 11152 10746 11204 10752
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 14200 10062 14228 11070
rect 14660 10742 14688 11154
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 9968 9382 9996 9998
rect 13832 9926 13860 9998
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 11955 9820 12263 9829
rect 11955 9818 11961 9820
rect 12017 9818 12041 9820
rect 12097 9818 12121 9820
rect 12177 9818 12201 9820
rect 12257 9818 12263 9820
rect 12017 9766 12019 9818
rect 12199 9766 12201 9818
rect 11955 9764 11961 9766
rect 12017 9764 12041 9766
rect 12097 9764 12121 9766
rect 12177 9764 12201 9766
rect 12257 9764 12263 9766
rect 11955 9755 12263 9764
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 10796 8974 10824 9318
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10796 8430 10824 8910
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8102 7100 8410 7109
rect 8102 7098 8108 7100
rect 8164 7098 8188 7100
rect 8244 7098 8268 7100
rect 8324 7098 8348 7100
rect 8404 7098 8410 7100
rect 8164 7046 8166 7098
rect 8346 7046 8348 7098
rect 8102 7044 8108 7046
rect 8164 7044 8188 7046
rect 8244 7044 8268 7046
rect 8324 7044 8348 7046
rect 8404 7044 8410 7046
rect 8102 7035 8410 7044
rect 9416 7002 9444 7278
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9692 6798 9720 7686
rect 10336 7546 10364 7890
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 9876 7002 9904 7278
rect 10428 7002 10456 7278
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7852 6225 7880 6598
rect 9692 6254 9720 6734
rect 10152 6458 10180 6870
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10704 6458 10732 6598
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 9680 6248 9732 6254
rect 7838 6216 7894 6225
rect 9680 6190 9732 6196
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 7838 6151 7894 6160
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 8102 6012 8410 6021
rect 8102 6010 8108 6012
rect 8164 6010 8188 6012
rect 8244 6010 8268 6012
rect 8324 6010 8348 6012
rect 8404 6010 8410 6012
rect 8164 5958 8166 6010
rect 8346 5958 8348 6010
rect 8102 5956 8108 5958
rect 8164 5956 8188 5958
rect 8244 5956 8268 5958
rect 8324 5956 8348 5958
rect 8404 5956 8410 5958
rect 8102 5947 8410 5956
rect 8102 4924 8410 4933
rect 8102 4922 8108 4924
rect 8164 4922 8188 4924
rect 8244 4922 8268 4924
rect 8324 4922 8348 4924
rect 8404 4922 8410 4924
rect 8164 4870 8166 4922
rect 8346 4870 8348 4922
rect 8102 4868 8108 4870
rect 8164 4868 8188 4870
rect 8244 4868 8268 4870
rect 8324 4868 8348 4870
rect 8404 4868 8410 4870
rect 8102 4859 8410 4868
rect 8102 3836 8410 3845
rect 8102 3834 8108 3836
rect 8164 3834 8188 3836
rect 8244 3834 8268 3836
rect 8324 3834 8348 3836
rect 8404 3834 8410 3836
rect 8164 3782 8166 3834
rect 8346 3782 8348 3834
rect 8102 3780 8108 3782
rect 8164 3780 8188 3782
rect 8244 3780 8268 3782
rect 8324 3780 8348 3782
rect 8404 3780 8410 3782
rect 8102 3771 8410 3780
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 7116 2746 7236 2774
rect 8102 2748 8410 2757
rect 8102 2746 8108 2748
rect 8164 2746 8188 2748
rect 8244 2746 8268 2748
rect 8324 2746 8348 2748
rect 8404 2746 8410 2748
rect 4250 2204 4558 2213
rect 4250 2202 4256 2204
rect 4312 2202 4336 2204
rect 4392 2202 4416 2204
rect 4472 2202 4496 2204
rect 4552 2202 4558 2204
rect 4312 2150 4314 2202
rect 4494 2150 4496 2202
rect 4250 2148 4256 2150
rect 4312 2148 4336 2150
rect 4392 2148 4416 2150
rect 4472 2148 4496 2150
rect 4552 2148 4558 2150
rect 4250 2139 4558 2148
rect 4250 1116 4558 1125
rect 4250 1114 4256 1116
rect 4312 1114 4336 1116
rect 4392 1114 4416 1116
rect 4472 1114 4496 1116
rect 4552 1114 4558 1116
rect 4312 1062 4314 1114
rect 4494 1062 4496 1114
rect 4250 1060 4256 1062
rect 4312 1060 4336 1062
rect 4392 1060 4416 1062
rect 4472 1060 4496 1062
rect 4552 1060 4558 1062
rect 4250 1051 4558 1060
rect 7116 400 7144 2746
rect 8164 2694 8166 2746
rect 8346 2694 8348 2746
rect 8102 2692 8108 2694
rect 8164 2692 8188 2694
rect 8244 2692 8268 2694
rect 8324 2692 8348 2694
rect 8404 2692 8410 2694
rect 8102 2683 8410 2692
rect 8102 1660 8410 1669
rect 8102 1658 8108 1660
rect 8164 1658 8188 1660
rect 8244 1658 8268 1660
rect 8324 1658 8348 1660
rect 8404 1658 8410 1660
rect 8164 1606 8166 1658
rect 8346 1606 8348 1658
rect 8102 1604 8108 1606
rect 8164 1604 8188 1606
rect 8244 1604 8268 1606
rect 8324 1604 8348 1606
rect 8404 1604 8410 1606
rect 8102 1595 8410 1604
rect 8102 572 8410 581
rect 8102 570 8108 572
rect 8164 570 8188 572
rect 8244 570 8268 572
rect 8324 570 8348 572
rect 8404 570 8410 572
rect 8164 518 8166 570
rect 8346 518 8348 570
rect 8102 516 8108 518
rect 8164 516 8188 518
rect 8244 516 8268 518
rect 8324 516 8348 518
rect 8404 516 8410 518
rect 8102 507 8410 516
rect 9048 400 9076 3402
rect 9692 400 9720 6054
rect 10520 5778 10548 6190
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10336 400 10364 4082
rect 10980 400 11008 7686
rect 11256 4146 11284 9318
rect 11955 8732 12263 8741
rect 11955 8730 11961 8732
rect 12017 8730 12041 8732
rect 12097 8730 12121 8732
rect 12177 8730 12201 8732
rect 12257 8730 12263 8732
rect 12017 8678 12019 8730
rect 12199 8678 12201 8730
rect 11955 8676 11961 8678
rect 12017 8676 12041 8678
rect 12097 8676 12121 8678
rect 12177 8676 12201 8678
rect 12257 8676 12263 8678
rect 11955 8667 12263 8676
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11348 6458 11376 6598
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11440 2774 11468 8230
rect 11955 7644 12263 7653
rect 11955 7642 11961 7644
rect 12017 7642 12041 7644
rect 12097 7642 12121 7644
rect 12177 7642 12201 7644
rect 12257 7642 12263 7644
rect 12017 7590 12019 7642
rect 12199 7590 12201 7642
rect 11955 7588 11961 7590
rect 12017 7588 12041 7590
rect 12097 7588 12121 7590
rect 12177 7588 12201 7590
rect 12257 7588 12263 7590
rect 11955 7579 12263 7588
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 11992 6934 12020 7414
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 12268 6866 12296 7278
rect 12544 7206 12572 7414
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12360 7002 12388 7142
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11624 5914 11652 6598
rect 11955 6556 12263 6565
rect 11955 6554 11961 6556
rect 12017 6554 12041 6556
rect 12097 6554 12121 6556
rect 12177 6554 12201 6556
rect 12257 6554 12263 6556
rect 12017 6502 12019 6554
rect 12199 6502 12201 6554
rect 11955 6500 11961 6502
rect 12017 6500 12041 6502
rect 12097 6500 12121 6502
rect 12177 6500 12201 6502
rect 12257 6500 12263 6502
rect 11955 6491 12263 6500
rect 12544 6186 12572 7142
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 11955 5468 12263 5477
rect 11955 5466 11961 5468
rect 12017 5466 12041 5468
rect 12097 5466 12121 5468
rect 12177 5466 12201 5468
rect 12257 5466 12263 5468
rect 12017 5414 12019 5466
rect 12199 5414 12201 5466
rect 11955 5412 11961 5414
rect 12017 5412 12041 5414
rect 12097 5412 12121 5414
rect 12177 5412 12201 5414
rect 12257 5412 12263 5414
rect 11955 5403 12263 5412
rect 11955 4380 12263 4389
rect 11955 4378 11961 4380
rect 12017 4378 12041 4380
rect 12097 4378 12121 4380
rect 12177 4378 12201 4380
rect 12257 4378 12263 4380
rect 12017 4326 12019 4378
rect 12199 4326 12201 4378
rect 11955 4324 11961 4326
rect 12017 4324 12041 4326
rect 12097 4324 12121 4326
rect 12177 4324 12201 4326
rect 12257 4324 12263 4326
rect 11955 4315 12263 4324
rect 11955 3292 12263 3301
rect 11955 3290 11961 3292
rect 12017 3290 12041 3292
rect 12097 3290 12121 3292
rect 12177 3290 12201 3292
rect 12257 3290 12263 3292
rect 12017 3238 12019 3290
rect 12199 3238 12201 3290
rect 11955 3236 11961 3238
rect 12017 3236 12041 3238
rect 12097 3236 12121 3238
rect 12177 3236 12201 3238
rect 12257 3236 12263 3238
rect 11955 3227 12263 3236
rect 11440 2746 11652 2774
rect 11624 400 11652 2746
rect 11955 2204 12263 2213
rect 11955 2202 11961 2204
rect 12017 2202 12041 2204
rect 12097 2202 12121 2204
rect 12177 2202 12201 2204
rect 12257 2202 12263 2204
rect 12017 2150 12019 2202
rect 12199 2150 12201 2202
rect 11955 2148 11961 2150
rect 12017 2148 12041 2150
rect 12097 2148 12121 2150
rect 12177 2148 12201 2150
rect 12257 2148 12263 2150
rect 11955 2139 12263 2148
rect 11955 1116 12263 1125
rect 11955 1114 11961 1116
rect 12017 1114 12041 1116
rect 12097 1114 12121 1116
rect 12177 1114 12201 1116
rect 12257 1114 12263 1116
rect 12017 1062 12019 1114
rect 12199 1062 12201 1114
rect 11955 1060 11961 1062
rect 12017 1060 12041 1062
rect 12097 1060 12121 1062
rect 12177 1060 12201 1062
rect 12257 1060 12263 1062
rect 11955 1051 12263 1060
rect 12360 898 12388 5510
rect 12636 3466 12664 9862
rect 13832 9654 13860 9862
rect 14384 9722 14412 10406
rect 14476 10266 14504 10406
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14476 9926 14504 10202
rect 14660 10130 14688 10678
rect 15304 10606 15332 10950
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15304 10130 15332 10542
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15396 10266 15424 10406
rect 15807 10364 16115 10373
rect 15807 10362 15813 10364
rect 15869 10362 15893 10364
rect 15949 10362 15973 10364
rect 16029 10362 16053 10364
rect 16109 10362 16115 10364
rect 15869 10310 15871 10362
rect 16051 10310 16053 10362
rect 15807 10308 15813 10310
rect 15869 10308 15893 10310
rect 15949 10308 15973 10310
rect 16029 10308 16053 10310
rect 16109 10308 16115 10310
rect 15807 10299 16115 10308
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 14660 10010 14688 10066
rect 14660 9994 14872 10010
rect 14660 9988 14884 9994
rect 14660 9982 14832 9988
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13004 8498 13032 9522
rect 14660 9518 14688 9982
rect 14832 9930 14884 9936
rect 15304 9926 15332 10066
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 14936 9518 14964 9862
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 9178 13216 9386
rect 15856 9382 15884 9862
rect 15948 9722 15976 10066
rect 16592 9722 16620 10610
rect 17604 9926 17632 12242
rect 18708 11762 18736 12378
rect 19352 11898 19380 19600
rect 19660 18524 19968 18533
rect 19660 18522 19666 18524
rect 19722 18522 19746 18524
rect 19802 18522 19826 18524
rect 19882 18522 19906 18524
rect 19962 18522 19968 18524
rect 19722 18470 19724 18522
rect 19904 18470 19906 18522
rect 19660 18468 19666 18470
rect 19722 18468 19746 18470
rect 19802 18468 19826 18470
rect 19882 18468 19906 18470
rect 19962 18468 19968 18470
rect 19660 18459 19968 18468
rect 19660 17436 19968 17445
rect 19660 17434 19666 17436
rect 19722 17434 19746 17436
rect 19802 17434 19826 17436
rect 19882 17434 19906 17436
rect 19962 17434 19968 17436
rect 19722 17382 19724 17434
rect 19904 17382 19906 17434
rect 19660 17380 19666 17382
rect 19722 17380 19746 17382
rect 19802 17380 19826 17382
rect 19882 17380 19906 17382
rect 19962 17380 19968 17382
rect 19660 17371 19968 17380
rect 19660 16348 19968 16357
rect 19660 16346 19666 16348
rect 19722 16346 19746 16348
rect 19802 16346 19826 16348
rect 19882 16346 19906 16348
rect 19962 16346 19968 16348
rect 19722 16294 19724 16346
rect 19904 16294 19906 16346
rect 19660 16292 19666 16294
rect 19722 16292 19746 16294
rect 19802 16292 19826 16294
rect 19882 16292 19906 16294
rect 19962 16292 19968 16294
rect 19660 16283 19968 16292
rect 19660 15260 19968 15269
rect 19660 15258 19666 15260
rect 19722 15258 19746 15260
rect 19802 15258 19826 15260
rect 19882 15258 19906 15260
rect 19962 15258 19968 15260
rect 19722 15206 19724 15258
rect 19904 15206 19906 15258
rect 19660 15204 19666 15206
rect 19722 15204 19746 15206
rect 19802 15204 19826 15206
rect 19882 15204 19906 15206
rect 19962 15204 19968 15206
rect 19660 15195 19968 15204
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19444 13870 19472 14214
rect 19660 14172 19968 14181
rect 19660 14170 19666 14172
rect 19722 14170 19746 14172
rect 19802 14170 19826 14172
rect 19882 14170 19906 14172
rect 19962 14170 19968 14172
rect 19722 14118 19724 14170
rect 19904 14118 19906 14170
rect 19660 14116 19666 14118
rect 19722 14116 19746 14118
rect 19802 14116 19826 14118
rect 19882 14116 19906 14118
rect 19962 14116 19968 14118
rect 19660 14107 19968 14116
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 13326 19472 13806
rect 19996 13530 20024 19600
rect 20640 14074 20668 19600
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19444 12986 19472 13262
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19444 12306 19472 12922
rect 19536 12918 19564 13330
rect 19628 13274 19656 13330
rect 19628 13246 20024 13274
rect 19660 13084 19968 13093
rect 19660 13082 19666 13084
rect 19722 13082 19746 13084
rect 19802 13082 19826 13084
rect 19882 13082 19906 13084
rect 19962 13082 19968 13084
rect 19722 13030 19724 13082
rect 19904 13030 19906 13082
rect 19660 13028 19666 13030
rect 19722 13028 19746 13030
rect 19802 13028 19826 13030
rect 19882 13028 19906 13030
rect 19962 13028 19968 13030
rect 19660 13019 19968 13028
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19996 12850 20024 13246
rect 20456 12986 20484 13670
rect 20640 13462 20668 13670
rect 20628 13456 20680 13462
rect 20628 13398 20680 13404
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 20180 12646 20208 12854
rect 20456 12714 20484 12922
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 19904 12442 19932 12582
rect 20456 12442 20484 12650
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19536 11898 19564 12038
rect 19660 11996 19968 12005
rect 19660 11994 19666 11996
rect 19722 11994 19746 11996
rect 19802 11994 19826 11996
rect 19882 11994 19906 11996
rect 19962 11994 19968 11996
rect 19722 11942 19724 11994
rect 19904 11942 19906 11994
rect 19660 11940 19666 11942
rect 19722 11940 19746 11942
rect 19802 11940 19826 11942
rect 19882 11940 19906 11942
rect 19962 11940 19968 11942
rect 19660 11931 19968 11940
rect 20364 11898 20392 12106
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18064 11218 18092 11630
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 18064 10674 18092 11154
rect 19352 11150 19380 11494
rect 20548 11218 20576 12786
rect 20640 12730 20668 13398
rect 20640 12702 20760 12730
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20640 12306 20668 12582
rect 20732 12306 20760 12702
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 20640 11898 20668 12038
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20916 11354 20944 11834
rect 21008 11354 21036 12038
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 21100 11354 21128 11494
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19660 10908 19968 10917
rect 19660 10906 19666 10908
rect 19722 10906 19746 10908
rect 19802 10906 19826 10908
rect 19882 10906 19906 10908
rect 19962 10906 19968 10908
rect 19722 10854 19724 10906
rect 19904 10854 19906 10906
rect 19660 10852 19666 10854
rect 19722 10852 19746 10854
rect 19802 10852 19826 10854
rect 19882 10852 19906 10854
rect 19962 10852 19968 10854
rect 19660 10843 19968 10852
rect 21284 10810 21312 19600
rect 21928 13530 21956 19600
rect 23512 19068 23820 19077
rect 23512 19066 23518 19068
rect 23574 19066 23598 19068
rect 23654 19066 23678 19068
rect 23734 19066 23758 19068
rect 23814 19066 23820 19068
rect 23574 19014 23576 19066
rect 23756 19014 23758 19066
rect 23512 19012 23518 19014
rect 23574 19012 23598 19014
rect 23654 19012 23678 19014
rect 23734 19012 23758 19014
rect 23814 19012 23820 19014
rect 23512 19003 23820 19012
rect 31217 19068 31525 19077
rect 31217 19066 31223 19068
rect 31279 19066 31303 19068
rect 31359 19066 31383 19068
rect 31439 19066 31463 19068
rect 31519 19066 31525 19068
rect 31279 19014 31281 19066
rect 31461 19014 31463 19066
rect 31217 19012 31223 19014
rect 31279 19012 31303 19014
rect 31359 19012 31383 19014
rect 31439 19012 31463 19014
rect 31519 19012 31525 19014
rect 31217 19003 31525 19012
rect 27365 18524 27673 18533
rect 27365 18522 27371 18524
rect 27427 18522 27451 18524
rect 27507 18522 27531 18524
rect 27587 18522 27611 18524
rect 27667 18522 27673 18524
rect 27427 18470 27429 18522
rect 27609 18470 27611 18522
rect 27365 18468 27371 18470
rect 27427 18468 27451 18470
rect 27507 18468 27531 18470
rect 27587 18468 27611 18470
rect 27667 18468 27673 18470
rect 27365 18459 27673 18468
rect 23512 17980 23820 17989
rect 23512 17978 23518 17980
rect 23574 17978 23598 17980
rect 23654 17978 23678 17980
rect 23734 17978 23758 17980
rect 23814 17978 23820 17980
rect 23574 17926 23576 17978
rect 23756 17926 23758 17978
rect 23512 17924 23518 17926
rect 23574 17924 23598 17926
rect 23654 17924 23678 17926
rect 23734 17924 23758 17926
rect 23814 17924 23820 17926
rect 23512 17915 23820 17924
rect 31217 17980 31525 17989
rect 31217 17978 31223 17980
rect 31279 17978 31303 17980
rect 31359 17978 31383 17980
rect 31439 17978 31463 17980
rect 31519 17978 31525 17980
rect 31279 17926 31281 17978
rect 31461 17926 31463 17978
rect 31217 17924 31223 17926
rect 31279 17924 31303 17926
rect 31359 17924 31383 17926
rect 31439 17924 31463 17926
rect 31519 17924 31525 17926
rect 31217 17915 31525 17924
rect 27365 17436 27673 17445
rect 27365 17434 27371 17436
rect 27427 17434 27451 17436
rect 27507 17434 27531 17436
rect 27587 17434 27611 17436
rect 27667 17434 27673 17436
rect 27427 17382 27429 17434
rect 27609 17382 27611 17434
rect 27365 17380 27371 17382
rect 27427 17380 27451 17382
rect 27507 17380 27531 17382
rect 27587 17380 27611 17382
rect 27667 17380 27673 17382
rect 27365 17371 27673 17380
rect 23512 16892 23820 16901
rect 23512 16890 23518 16892
rect 23574 16890 23598 16892
rect 23654 16890 23678 16892
rect 23734 16890 23758 16892
rect 23814 16890 23820 16892
rect 23574 16838 23576 16890
rect 23756 16838 23758 16890
rect 23512 16836 23518 16838
rect 23574 16836 23598 16838
rect 23654 16836 23678 16838
rect 23734 16836 23758 16838
rect 23814 16836 23820 16838
rect 23512 16827 23820 16836
rect 31217 16892 31525 16901
rect 31217 16890 31223 16892
rect 31279 16890 31303 16892
rect 31359 16890 31383 16892
rect 31439 16890 31463 16892
rect 31519 16890 31525 16892
rect 31279 16838 31281 16890
rect 31461 16838 31463 16890
rect 31217 16836 31223 16838
rect 31279 16836 31303 16838
rect 31359 16836 31383 16838
rect 31439 16836 31463 16838
rect 31519 16836 31525 16838
rect 31217 16827 31525 16836
rect 27365 16348 27673 16357
rect 27365 16346 27371 16348
rect 27427 16346 27451 16348
rect 27507 16346 27531 16348
rect 27587 16346 27611 16348
rect 27667 16346 27673 16348
rect 27427 16294 27429 16346
rect 27609 16294 27611 16346
rect 27365 16292 27371 16294
rect 27427 16292 27451 16294
rect 27507 16292 27531 16294
rect 27587 16292 27611 16294
rect 27667 16292 27673 16294
rect 27365 16283 27673 16292
rect 23512 15804 23820 15813
rect 23512 15802 23518 15804
rect 23574 15802 23598 15804
rect 23654 15802 23678 15804
rect 23734 15802 23758 15804
rect 23814 15802 23820 15804
rect 23574 15750 23576 15802
rect 23756 15750 23758 15802
rect 23512 15748 23518 15750
rect 23574 15748 23598 15750
rect 23654 15748 23678 15750
rect 23734 15748 23758 15750
rect 23814 15748 23820 15750
rect 23512 15739 23820 15748
rect 31217 15804 31525 15813
rect 31217 15802 31223 15804
rect 31279 15802 31303 15804
rect 31359 15802 31383 15804
rect 31439 15802 31463 15804
rect 31519 15802 31525 15804
rect 31279 15750 31281 15802
rect 31461 15750 31463 15802
rect 31217 15748 31223 15750
rect 31279 15748 31303 15750
rect 31359 15748 31383 15750
rect 31439 15748 31463 15750
rect 31519 15748 31525 15750
rect 31217 15739 31525 15748
rect 27365 15260 27673 15269
rect 27365 15258 27371 15260
rect 27427 15258 27451 15260
rect 27507 15258 27531 15260
rect 27587 15258 27611 15260
rect 27667 15258 27673 15260
rect 27427 15206 27429 15258
rect 27609 15206 27611 15258
rect 27365 15204 27371 15206
rect 27427 15204 27451 15206
rect 27507 15204 27531 15206
rect 27587 15204 27611 15206
rect 27667 15204 27673 15206
rect 27365 15195 27673 15204
rect 27986 15056 28042 15065
rect 27986 14991 28042 15000
rect 23512 14716 23820 14725
rect 23512 14714 23518 14716
rect 23574 14714 23598 14716
rect 23654 14714 23678 14716
rect 23734 14714 23758 14716
rect 23814 14714 23820 14716
rect 23574 14662 23576 14714
rect 23756 14662 23758 14714
rect 23512 14660 23518 14662
rect 23574 14660 23598 14662
rect 23654 14660 23678 14662
rect 23734 14660 23758 14662
rect 23814 14660 23820 14662
rect 23512 14651 23820 14660
rect 27365 14172 27673 14181
rect 27365 14170 27371 14172
rect 27427 14170 27451 14172
rect 27507 14170 27531 14172
rect 27587 14170 27611 14172
rect 27667 14170 27673 14172
rect 27427 14118 27429 14170
rect 27609 14118 27611 14170
rect 27365 14116 27371 14118
rect 27427 14116 27451 14118
rect 27507 14116 27531 14118
rect 27587 14116 27611 14118
rect 27667 14116 27673 14118
rect 27365 14107 27673 14116
rect 23512 13628 23820 13637
rect 23512 13626 23518 13628
rect 23574 13626 23598 13628
rect 23654 13626 23678 13628
rect 23734 13626 23758 13628
rect 23814 13626 23820 13628
rect 23574 13574 23576 13626
rect 23756 13574 23758 13626
rect 23512 13572 23518 13574
rect 23574 13572 23598 13574
rect 23654 13572 23678 13574
rect 23734 13572 23758 13574
rect 23814 13572 23820 13574
rect 23512 13563 23820 13572
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 27365 13084 27673 13093
rect 27365 13082 27371 13084
rect 27427 13082 27451 13084
rect 27507 13082 27531 13084
rect 27587 13082 27611 13084
rect 27667 13082 27673 13084
rect 27427 13030 27429 13082
rect 27609 13030 27611 13082
rect 27365 13028 27371 13030
rect 27427 13028 27451 13030
rect 27507 13028 27531 13030
rect 27587 13028 27611 13030
rect 27667 13028 27673 13030
rect 27365 13019 27673 13028
rect 28000 12918 28028 14991
rect 31217 14716 31525 14725
rect 31217 14714 31223 14716
rect 31279 14714 31303 14716
rect 31359 14714 31383 14716
rect 31439 14714 31463 14716
rect 31519 14714 31525 14716
rect 31279 14662 31281 14714
rect 31461 14662 31463 14714
rect 31217 14660 31223 14662
rect 31279 14660 31303 14662
rect 31359 14660 31383 14662
rect 31439 14660 31463 14662
rect 31519 14660 31525 14662
rect 31217 14651 31525 14660
rect 28446 14376 28502 14385
rect 28446 14311 28502 14320
rect 28262 13016 28318 13025
rect 28262 12951 28264 12960
rect 28316 12951 28318 12960
rect 28264 12922 28316 12928
rect 27988 12912 28040 12918
rect 27988 12854 28040 12860
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22204 12442 22232 12718
rect 23512 12540 23820 12549
rect 23512 12538 23518 12540
rect 23574 12538 23598 12540
rect 23654 12538 23678 12540
rect 23734 12538 23758 12540
rect 23814 12538 23820 12540
rect 23574 12486 23576 12538
rect 23756 12486 23758 12538
rect 23512 12484 23518 12486
rect 23574 12484 23598 12486
rect 23654 12484 23678 12486
rect 23734 12484 23758 12486
rect 23814 12484 23820 12486
rect 23512 12475 23820 12484
rect 28460 12442 28488 14311
rect 31666 13696 31722 13705
rect 31217 13628 31525 13637
rect 31666 13631 31722 13640
rect 31217 13626 31223 13628
rect 31279 13626 31303 13628
rect 31359 13626 31383 13628
rect 31439 13626 31463 13628
rect 31519 13626 31525 13628
rect 31279 13574 31281 13626
rect 31461 13574 31463 13626
rect 31217 13572 31223 13574
rect 31279 13572 31303 13574
rect 31359 13572 31383 13574
rect 31439 13572 31463 13574
rect 31519 13572 31525 13574
rect 31217 13563 31525 13572
rect 31680 12986 31708 13631
rect 28540 12980 28592 12986
rect 28540 12922 28592 12928
rect 31668 12980 31720 12986
rect 31668 12922 31720 12928
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 28448 12436 28500 12442
rect 28448 12378 28500 12384
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 11218 21404 11494
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18064 10130 18092 10610
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13280 9042 13308 9318
rect 13648 9178 13676 9318
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13924 9110 13952 9318
rect 15807 9276 16115 9285
rect 15807 9274 15813 9276
rect 15869 9274 15893 9276
rect 15949 9274 15973 9276
rect 16029 9274 16053 9276
rect 16109 9274 16115 9276
rect 15869 9222 15871 9274
rect 16051 9222 16053 9274
rect 15807 9220 15813 9222
rect 15869 9220 15893 9222
rect 15949 9220 15973 9222
rect 16029 9220 16053 9222
rect 16109 9220 16115 9222
rect 15807 9211 16115 9220
rect 17328 9110 17356 9454
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13188 8430 13216 8842
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 14016 8430 14044 8774
rect 14292 8566 14320 8774
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14292 8430 14320 8502
rect 14660 8430 14688 8774
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13280 8090 13308 8230
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13464 7954 13492 8230
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13832 7834 13860 8026
rect 13924 7954 13952 8298
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14016 7834 14044 7890
rect 13728 7812 13780 7818
rect 13832 7806 14228 7834
rect 13728 7754 13780 7760
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 7546 12940 7686
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12912 7342 12940 7482
rect 13740 7410 13768 7754
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7410 14136 7686
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14200 7342 14228 7806
rect 14660 7750 14688 8366
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14752 7886 14780 8230
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12268 870 12388 898
rect 12268 400 12296 870
rect 12912 400 12940 6938
rect 14108 6934 14136 7142
rect 14476 7002 14504 7142
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14096 6928 14148 6934
rect 14096 6870 14148 6876
rect 14660 6662 14688 7686
rect 14752 7546 14780 7822
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14660 6254 14688 6598
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13556 400 13584 6054
rect 14660 5846 14688 6190
rect 14648 5840 14700 5846
rect 14648 5782 14700 5788
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14200 400 14228 5510
rect 15028 2774 15056 6598
rect 14844 2746 15056 2774
rect 14844 400 14872 2746
rect 15488 400 15516 8774
rect 15807 8188 16115 8197
rect 15807 8186 15813 8188
rect 15869 8186 15893 8188
rect 15949 8186 15973 8188
rect 16029 8186 16053 8188
rect 16109 8186 16115 8188
rect 15869 8134 15871 8186
rect 16051 8134 16053 8186
rect 15807 8132 15813 8134
rect 15869 8132 15893 8134
rect 15949 8132 15973 8134
rect 16029 8132 16053 8134
rect 16109 8132 16115 8134
rect 15807 8123 16115 8132
rect 16224 8022 16252 8910
rect 17604 8362 17632 9862
rect 18064 9722 18092 9862
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 18156 9450 18184 10066
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 19660 9820 19968 9829
rect 19660 9818 19666 9820
rect 19722 9818 19746 9820
rect 19802 9818 19826 9820
rect 19882 9818 19906 9820
rect 19962 9818 19968 9820
rect 19722 9766 19724 9818
rect 19904 9766 19906 9818
rect 19660 9764 19666 9766
rect 19722 9764 19746 9766
rect 19802 9764 19826 9766
rect 19882 9764 19906 9766
rect 19962 9764 19968 9766
rect 19660 9755 19968 9764
rect 20916 9722 20944 9862
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18984 9178 19012 9454
rect 18328 9172 18380 9178
rect 18972 9172 19024 9178
rect 18380 9132 18460 9160
rect 18328 9114 18380 9120
rect 18340 9042 18368 9114
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18432 8974 18460 9132
rect 18972 9114 19024 9120
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18800 8838 18828 8978
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 15807 7100 16115 7109
rect 15807 7098 15813 7100
rect 15869 7098 15893 7100
rect 15949 7098 15973 7100
rect 16029 7098 16053 7100
rect 16109 7098 16115 7100
rect 15869 7046 15871 7098
rect 16051 7046 16053 7098
rect 15807 7044 15813 7046
rect 15869 7044 15893 7046
rect 15949 7044 15973 7046
rect 16029 7044 16053 7046
rect 16109 7044 16115 7046
rect 15807 7035 16115 7044
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 15807 6012 16115 6021
rect 15807 6010 15813 6012
rect 15869 6010 15893 6012
rect 15949 6010 15973 6012
rect 16029 6010 16053 6012
rect 16109 6010 16115 6012
rect 15869 5958 15871 6010
rect 16051 5958 16053 6010
rect 15807 5956 15813 5958
rect 15869 5956 15893 5958
rect 15949 5956 15973 5958
rect 16029 5956 16053 5958
rect 16109 5956 16115 5958
rect 15807 5947 16115 5956
rect 16224 5914 16252 6122
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16224 5370 16252 5646
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 15807 4924 16115 4933
rect 15807 4922 15813 4924
rect 15869 4922 15893 4924
rect 15949 4922 15973 4924
rect 16029 4922 16053 4924
rect 16109 4922 16115 4924
rect 15869 4870 15871 4922
rect 16051 4870 16053 4922
rect 15807 4868 15813 4870
rect 15869 4868 15893 4870
rect 15949 4868 15973 4870
rect 16029 4868 16053 4870
rect 16109 4868 16115 4870
rect 15807 4859 16115 4868
rect 15807 3836 16115 3845
rect 15807 3834 15813 3836
rect 15869 3834 15893 3836
rect 15949 3834 15973 3836
rect 16029 3834 16053 3836
rect 16109 3834 16115 3836
rect 15869 3782 15871 3834
rect 16051 3782 16053 3834
rect 15807 3780 15813 3782
rect 15869 3780 15893 3782
rect 15949 3780 15973 3782
rect 16029 3780 16053 3782
rect 16109 3780 16115 3782
rect 15807 3771 16115 3780
rect 15807 2748 16115 2757
rect 15807 2746 15813 2748
rect 15869 2746 15893 2748
rect 15949 2746 15973 2748
rect 16029 2746 16053 2748
rect 16109 2746 16115 2748
rect 15869 2694 15871 2746
rect 16051 2694 16053 2746
rect 15807 2692 15813 2694
rect 15869 2692 15893 2694
rect 15949 2692 15973 2694
rect 16029 2692 16053 2694
rect 16109 2692 16115 2694
rect 15807 2683 16115 2692
rect 15807 1660 16115 1669
rect 15807 1658 15813 1660
rect 15869 1658 15893 1660
rect 15949 1658 15973 1660
rect 16029 1658 16053 1660
rect 16109 1658 16115 1660
rect 15869 1606 15871 1658
rect 16051 1606 16053 1658
rect 15807 1604 15813 1606
rect 15869 1604 15893 1606
rect 15949 1604 15973 1606
rect 16029 1604 16053 1606
rect 16109 1604 16115 1606
rect 15807 1595 16115 1604
rect 16224 882 16252 5102
rect 16212 876 16264 882
rect 16212 818 16264 824
rect 15807 572 16115 581
rect 15807 570 15813 572
rect 15869 570 15893 572
rect 15949 570 15973 572
rect 16029 570 16053 572
rect 16109 570 16115 572
rect 15869 518 15871 570
rect 16051 518 16053 570
rect 15807 516 15813 518
rect 15869 516 15893 518
rect 15949 516 15973 518
rect 16029 516 16053 518
rect 16109 516 16115 518
rect 15807 507 16115 516
rect 16316 474 16344 8230
rect 17604 8090 17632 8298
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17052 7206 17080 7686
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17052 6866 17080 7142
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17052 6458 17080 6802
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16396 5636 16448 5642
rect 16396 5578 16448 5584
rect 16408 4826 16436 5578
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16500 4826 16528 5034
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16028 468 16080 474
rect 16304 468 16356 474
rect 16080 428 16160 456
rect 16028 410 16080 416
rect 16132 400 16160 428
rect 16304 410 16356 416
rect 16776 400 16804 6054
rect 17052 5234 17080 6394
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17236 5914 17264 6054
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17420 5574 17448 5714
rect 17408 5568 17460 5574
rect 17408 5510 17460 5516
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17512 2802 17540 7686
rect 17604 7342 17632 8026
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 17880 6446 18092 6474
rect 17880 6390 17908 6446
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17788 5914 17816 6258
rect 17776 5908 17828 5914
rect 17696 5868 17776 5896
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17604 5534 17632 5714
rect 17696 5642 17724 5868
rect 17776 5850 17828 5856
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17972 5534 18000 5714
rect 17604 5506 18000 5534
rect 17420 2774 17540 2802
rect 17420 400 17448 2774
rect 18064 400 18092 6446
rect 18156 6254 18184 6802
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18340 6322 18368 6598
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18156 5846 18184 6190
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18248 5914 18276 6054
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18144 5840 18196 5846
rect 18144 5782 18196 5788
rect 18248 5642 18276 5850
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18236 5636 18288 5642
rect 18236 5578 18288 5584
rect 18524 5166 18552 5714
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18708 400 18736 8774
rect 19352 8634 19380 9454
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19444 9178 19472 9386
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19444 8294 19472 8842
rect 19660 8732 19968 8741
rect 19660 8730 19666 8732
rect 19722 8730 19746 8732
rect 19802 8730 19826 8732
rect 19882 8730 19906 8732
rect 19962 8730 19968 8732
rect 19722 8678 19724 8730
rect 19904 8678 19906 8730
rect 19660 8676 19666 8678
rect 19722 8676 19746 8678
rect 19802 8676 19826 8678
rect 19882 8676 19906 8678
rect 19962 8676 19968 8678
rect 19660 8667 19968 8676
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19444 8090 19472 8230
rect 19628 8090 19656 8366
rect 19812 8362 19840 8570
rect 19996 8514 20024 8978
rect 20088 8838 20116 9114
rect 20720 9036 20772 9042
rect 20720 8978 20772 8984
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 19904 8486 20024 8514
rect 19800 8356 19852 8362
rect 19800 8298 19852 8304
rect 19904 8294 19932 8486
rect 20088 8362 20116 8774
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19904 8090 19932 8230
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 20088 7750 20116 8298
rect 20168 8016 20220 8022
rect 20168 7958 20220 7964
rect 20444 8016 20496 8022
rect 20444 7958 20496 7964
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 19660 7644 19968 7653
rect 19660 7642 19666 7644
rect 19722 7642 19746 7644
rect 19802 7642 19826 7644
rect 19882 7642 19906 7644
rect 19962 7642 19968 7644
rect 19722 7590 19724 7642
rect 19904 7590 19906 7642
rect 19660 7588 19666 7590
rect 19722 7588 19746 7590
rect 19802 7588 19826 7590
rect 19882 7588 19906 7590
rect 19962 7588 19968 7590
rect 19660 7579 19968 7588
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19444 7002 19472 7346
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19812 7002 19840 7278
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19444 6872 19472 6938
rect 19432 6866 19484 6872
rect 18788 6860 18840 6866
rect 19432 6808 19484 6814
rect 18788 6802 18840 6808
rect 18800 6458 18828 6802
rect 19076 6730 19380 6746
rect 19064 6724 19380 6730
rect 19116 6718 19380 6724
rect 19064 6666 19116 6672
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 19168 5914 19196 6598
rect 19248 6180 19300 6186
rect 19248 6122 19300 6128
rect 19260 5914 19288 6122
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19352 400 19380 6718
rect 19660 6556 19968 6565
rect 19660 6554 19666 6556
rect 19722 6554 19746 6556
rect 19802 6554 19826 6556
rect 19882 6554 19906 6556
rect 19962 6554 19968 6556
rect 19722 6502 19724 6554
rect 19904 6502 19906 6554
rect 19660 6500 19666 6502
rect 19722 6500 19746 6502
rect 19802 6500 19826 6502
rect 19882 6500 19906 6502
rect 19962 6500 19968 6502
rect 19660 6491 19968 6500
rect 19660 5468 19968 5477
rect 19660 5466 19666 5468
rect 19722 5466 19746 5468
rect 19802 5466 19826 5468
rect 19882 5466 19906 5468
rect 19962 5466 19968 5468
rect 19722 5414 19724 5466
rect 19904 5414 19906 5466
rect 19660 5412 19666 5414
rect 19722 5412 19746 5414
rect 19802 5412 19826 5414
rect 19882 5412 19906 5414
rect 19962 5412 19968 5414
rect 19660 5403 19968 5412
rect 19660 4380 19968 4389
rect 19660 4378 19666 4380
rect 19722 4378 19746 4380
rect 19802 4378 19826 4380
rect 19882 4378 19906 4380
rect 19962 4378 19968 4380
rect 19722 4326 19724 4378
rect 19904 4326 19906 4378
rect 19660 4324 19666 4326
rect 19722 4324 19746 4326
rect 19802 4324 19826 4326
rect 19882 4324 19906 4326
rect 19962 4324 19968 4326
rect 19660 4315 19968 4324
rect 19660 3292 19968 3301
rect 19660 3290 19666 3292
rect 19722 3290 19746 3292
rect 19802 3290 19826 3292
rect 19882 3290 19906 3292
rect 19962 3290 19968 3292
rect 19722 3238 19724 3290
rect 19904 3238 19906 3290
rect 19660 3236 19666 3238
rect 19722 3236 19746 3238
rect 19802 3236 19826 3238
rect 19882 3236 19906 3238
rect 19962 3236 19968 3238
rect 19660 3227 19968 3236
rect 19660 2204 19968 2213
rect 19660 2202 19666 2204
rect 19722 2202 19746 2204
rect 19802 2202 19826 2204
rect 19882 2202 19906 2204
rect 19962 2202 19968 2204
rect 19722 2150 19724 2202
rect 19904 2150 19906 2202
rect 19660 2148 19666 2150
rect 19722 2148 19746 2150
rect 19802 2148 19826 2150
rect 19882 2148 19906 2150
rect 19962 2148 19968 2150
rect 19660 2139 19968 2148
rect 19660 1116 19968 1125
rect 19660 1114 19666 1116
rect 19722 1114 19746 1116
rect 19802 1114 19826 1116
rect 19882 1114 19906 1116
rect 19962 1114 19968 1116
rect 19722 1062 19724 1114
rect 19904 1062 19906 1114
rect 19660 1060 19666 1062
rect 19722 1060 19746 1062
rect 19802 1060 19826 1062
rect 19882 1060 19906 1062
rect 19962 1060 19968 1062
rect 19660 1051 19968 1060
rect 19996 400 20024 7686
rect 20180 7546 20208 7958
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20272 7206 20300 7890
rect 20456 7818 20484 7958
rect 20548 7954 20576 8774
rect 20732 8090 20760 8978
rect 20916 8974 20944 9454
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21284 8634 21312 8910
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21560 8430 21588 12242
rect 22204 11762 22232 12378
rect 28262 12336 28318 12345
rect 22928 12300 22980 12306
rect 28262 12271 28318 12280
rect 22928 12242 22980 12248
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21652 10606 21680 11222
rect 22020 11218 22048 11562
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 22940 11150 22968 12242
rect 28276 12102 28304 12271
rect 28264 12096 28316 12102
rect 28264 12038 28316 12044
rect 27365 11996 27673 12005
rect 27365 11994 27371 11996
rect 27427 11994 27451 11996
rect 27507 11994 27531 11996
rect 27587 11994 27611 11996
rect 27667 11994 27673 11996
rect 27427 11942 27429 11994
rect 27609 11942 27611 11994
rect 27365 11940 27371 11942
rect 27427 11940 27451 11942
rect 27507 11940 27531 11942
rect 27587 11940 27611 11942
rect 27667 11940 27673 11942
rect 27365 11931 27673 11940
rect 28552 11898 28580 12922
rect 31217 12540 31525 12549
rect 31217 12538 31223 12540
rect 31279 12538 31303 12540
rect 31359 12538 31383 12540
rect 31439 12538 31463 12540
rect 31519 12538 31525 12540
rect 31279 12486 31281 12538
rect 31461 12486 31463 12538
rect 31217 12484 31223 12486
rect 31279 12484 31303 12486
rect 31359 12484 31383 12486
rect 31439 12484 31463 12486
rect 31519 12484 31525 12486
rect 31217 12475 31525 12484
rect 28540 11892 28592 11898
rect 28540 11834 28592 11840
rect 28262 11656 28318 11665
rect 28262 11591 28318 11600
rect 23512 11452 23820 11461
rect 23512 11450 23518 11452
rect 23574 11450 23598 11452
rect 23654 11450 23678 11452
rect 23734 11450 23758 11452
rect 23814 11450 23820 11452
rect 23574 11398 23576 11450
rect 23756 11398 23758 11450
rect 23512 11396 23518 11398
rect 23574 11396 23598 11398
rect 23654 11396 23678 11398
rect 23734 11396 23758 11398
rect 23814 11396 23820 11398
rect 23512 11387 23820 11396
rect 28276 11354 28304 11591
rect 31217 11452 31525 11461
rect 31217 11450 31223 11452
rect 31279 11450 31303 11452
rect 31359 11450 31383 11452
rect 31439 11450 31463 11452
rect 31519 11450 31525 11452
rect 31279 11398 31281 11450
rect 31461 11398 31463 11450
rect 31217 11396 31223 11398
rect 31279 11396 31303 11398
rect 31359 11396 31383 11398
rect 31439 11396 31463 11398
rect 31519 11396 31525 11398
rect 31217 11387 31525 11396
rect 28264 11348 28316 11354
rect 28264 11290 28316 11296
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22192 11076 22244 11082
rect 22192 11018 22244 11024
rect 22100 10736 22152 10742
rect 22100 10678 22152 10684
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 22020 10130 22048 10474
rect 22112 10146 22140 10678
rect 22204 10606 22232 11018
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22756 10742 22784 10950
rect 22744 10736 22796 10742
rect 22744 10678 22796 10684
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 22204 10266 22232 10406
rect 22296 10266 22324 10610
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22112 10130 22416 10146
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22112 10124 22428 10130
rect 22112 10118 22376 10124
rect 21824 10056 21876 10062
rect 21876 10004 21956 10010
rect 21824 9998 21956 10004
rect 21836 9982 21956 9998
rect 21928 9738 21956 9982
rect 22112 9926 22140 10118
rect 22376 10066 22428 10072
rect 22756 9994 22784 10542
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22848 10266 22876 10406
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22940 10130 22968 11086
rect 28262 10976 28318 10985
rect 27365 10908 27673 10917
rect 28262 10911 28318 10920
rect 27365 10906 27371 10908
rect 27427 10906 27451 10908
rect 27507 10906 27531 10908
rect 27587 10906 27611 10908
rect 27667 10906 27673 10908
rect 27427 10854 27429 10906
rect 27609 10854 27611 10906
rect 27365 10852 27371 10854
rect 27427 10852 27451 10854
rect 27507 10852 27531 10854
rect 27587 10852 27611 10854
rect 27667 10852 27673 10854
rect 27365 10843 27673 10852
rect 23512 10364 23820 10373
rect 23512 10362 23518 10364
rect 23574 10362 23598 10364
rect 23654 10362 23678 10364
rect 23734 10362 23758 10364
rect 23814 10362 23820 10364
rect 23574 10310 23576 10362
rect 23756 10310 23758 10362
rect 23512 10308 23518 10310
rect 23574 10308 23598 10310
rect 23654 10308 23678 10310
rect 23734 10308 23758 10310
rect 23814 10308 23820 10310
rect 23512 10299 23820 10308
rect 28276 10266 28304 10911
rect 31217 10364 31525 10373
rect 31217 10362 31223 10364
rect 31279 10362 31303 10364
rect 31359 10362 31383 10364
rect 31439 10362 31463 10364
rect 31519 10362 31525 10364
rect 31279 10310 31281 10362
rect 31461 10310 31463 10362
rect 31217 10308 31223 10310
rect 31279 10308 31303 10310
rect 31359 10308 31383 10310
rect 31439 10308 31463 10310
rect 31519 10308 31525 10310
rect 31217 10299 31525 10308
rect 31666 10296 31722 10305
rect 28264 10260 28316 10266
rect 31666 10231 31722 10240
rect 28264 10202 28316 10208
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 22744 9988 22796 9994
rect 22744 9930 22796 9936
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 22204 9738 22232 9862
rect 27365 9820 27673 9829
rect 27365 9818 27371 9820
rect 27427 9818 27451 9820
rect 27507 9818 27531 9820
rect 27587 9818 27611 9820
rect 27667 9818 27673 9820
rect 27427 9766 27429 9818
rect 27609 9766 27611 9818
rect 27365 9764 27371 9766
rect 27427 9764 27451 9766
rect 27507 9764 27531 9766
rect 27587 9764 27611 9766
rect 27667 9764 27673 9766
rect 27365 9755 27673 9764
rect 21928 9710 22232 9738
rect 31680 9722 31708 10231
rect 22204 9466 22232 9710
rect 31668 9716 31720 9722
rect 31668 9658 31720 9664
rect 28262 9616 28318 9625
rect 28262 9551 28318 9560
rect 28276 9518 28304 9551
rect 28264 9512 28316 9518
rect 22204 9450 22324 9466
rect 28264 9454 28316 9460
rect 22204 9444 22336 9450
rect 22204 9438 22284 9444
rect 22284 9386 22336 9392
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 21008 8090 21036 8230
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21652 8022 21680 8910
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21836 7954 21864 8570
rect 23400 8537 23428 9318
rect 23512 9276 23820 9285
rect 23512 9274 23518 9276
rect 23574 9274 23598 9276
rect 23654 9274 23678 9276
rect 23734 9274 23758 9276
rect 23814 9274 23820 9276
rect 23574 9222 23576 9274
rect 23756 9222 23758 9274
rect 23512 9220 23518 9222
rect 23574 9220 23598 9222
rect 23654 9220 23678 9222
rect 23734 9220 23758 9222
rect 23814 9220 23820 9222
rect 23512 9211 23820 9220
rect 31217 9276 31525 9285
rect 31217 9274 31223 9276
rect 31279 9274 31303 9276
rect 31359 9274 31383 9276
rect 31439 9274 31463 9276
rect 31519 9274 31525 9276
rect 31279 9222 31281 9274
rect 31461 9222 31463 9274
rect 31217 9220 31223 9222
rect 31279 9220 31303 9222
rect 31359 9220 31383 9222
rect 31439 9220 31463 9222
rect 31519 9220 31525 9222
rect 31217 9211 31525 9220
rect 28262 8936 28318 8945
rect 28262 8871 28318 8880
rect 27365 8732 27673 8741
rect 27365 8730 27371 8732
rect 27427 8730 27451 8732
rect 27507 8730 27531 8732
rect 27587 8730 27611 8732
rect 27667 8730 27673 8732
rect 27427 8678 27429 8730
rect 27609 8678 27611 8730
rect 27365 8676 27371 8678
rect 27427 8676 27451 8678
rect 27507 8676 27531 8678
rect 27587 8676 27611 8678
rect 27667 8676 27673 8678
rect 27365 8667 27673 8676
rect 28276 8566 28304 8871
rect 28448 8832 28500 8838
rect 28448 8774 28500 8780
rect 28264 8560 28316 8566
rect 23386 8528 23442 8537
rect 28264 8502 28316 8508
rect 23386 8463 23442 8472
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20548 7546 20576 7890
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21652 7546 21680 7822
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21836 7478 21864 7890
rect 22296 7546 22324 7958
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 21824 7472 21876 7478
rect 21824 7414 21876 7420
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20640 7002 20668 7414
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20732 7206 20760 7278
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 7002 20944 7142
rect 21836 7002 21864 7414
rect 23216 7342 23244 8366
rect 23296 8288 23348 8294
rect 23296 8230 23348 8236
rect 23308 8022 23336 8230
rect 23512 8188 23820 8197
rect 23512 8186 23518 8188
rect 23574 8186 23598 8188
rect 23654 8186 23678 8188
rect 23734 8186 23758 8188
rect 23814 8186 23820 8188
rect 23574 8134 23576 8186
rect 23756 8134 23758 8186
rect 23512 8132 23518 8134
rect 23574 8132 23598 8134
rect 23654 8132 23678 8134
rect 23734 8132 23758 8134
rect 23814 8132 23820 8134
rect 23512 8123 23820 8132
rect 23296 8016 23348 8022
rect 23296 7958 23348 7964
rect 28264 7744 28316 7750
rect 28264 7686 28316 7692
rect 27365 7644 27673 7653
rect 27365 7642 27371 7644
rect 27427 7642 27451 7644
rect 27507 7642 27531 7644
rect 27587 7642 27611 7644
rect 27667 7642 27673 7644
rect 27427 7590 27429 7642
rect 27609 7590 27611 7642
rect 27365 7588 27371 7590
rect 27427 7588 27451 7590
rect 27507 7588 27531 7590
rect 27587 7588 27611 7590
rect 27667 7588 27673 7590
rect 27365 7579 27673 7588
rect 28276 7585 28304 7686
rect 28262 7576 28318 7585
rect 28262 7511 28318 7520
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 28264 7200 28316 7206
rect 28264 7142 28316 7148
rect 23512 7100 23820 7109
rect 23512 7098 23518 7100
rect 23574 7098 23598 7100
rect 23654 7098 23678 7100
rect 23734 7098 23758 7100
rect 23814 7098 23820 7100
rect 23574 7046 23576 7098
rect 23756 7046 23758 7098
rect 23512 7044 23518 7046
rect 23574 7044 23598 7046
rect 23654 7044 23678 7046
rect 23734 7044 23758 7046
rect 23814 7044 23820 7046
rect 23512 7035 23820 7044
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 21824 6996 21876 7002
rect 21824 6938 21876 6944
rect 20076 6928 20128 6934
rect 28276 6905 28304 7142
rect 20076 6870 20128 6876
rect 28262 6896 28318 6905
rect 20088 6458 20116 6870
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 21088 6860 21140 6866
rect 28262 6831 28318 6840
rect 21088 6802 21140 6808
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20640 6186 20668 6802
rect 21100 6254 21128 6802
rect 28264 6656 28316 6662
rect 28264 6598 28316 6604
rect 27365 6556 27673 6565
rect 27365 6554 27371 6556
rect 27427 6554 27451 6556
rect 27507 6554 27531 6556
rect 27587 6554 27611 6556
rect 27667 6554 27673 6556
rect 27427 6502 27429 6554
rect 27609 6502 27611 6554
rect 27365 6500 27371 6502
rect 27427 6500 27451 6502
rect 27507 6500 27531 6502
rect 27587 6500 27611 6502
rect 27667 6500 27673 6502
rect 27365 6491 27673 6500
rect 21088 6248 21140 6254
rect 28276 6225 28304 6598
rect 21088 6190 21140 6196
rect 28262 6216 28318 6225
rect 20628 6180 20680 6186
rect 28262 6151 28318 6160
rect 20628 6122 20680 6128
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 20456 5534 20484 6054
rect 21744 5534 21772 6054
rect 23512 6012 23820 6021
rect 23512 6010 23518 6012
rect 23574 6010 23598 6012
rect 23654 6010 23678 6012
rect 23734 6010 23758 6012
rect 23814 6010 23820 6012
rect 23574 5958 23576 6010
rect 23756 5958 23758 6010
rect 23512 5956 23518 5958
rect 23574 5956 23598 5958
rect 23654 5956 23678 5958
rect 23734 5956 23758 5958
rect 23814 5956 23820 5958
rect 23512 5947 23820 5956
rect 28460 5545 28488 8774
rect 31666 8528 31722 8537
rect 31666 8463 31722 8472
rect 31680 8265 31708 8463
rect 31666 8256 31722 8265
rect 31217 8188 31525 8197
rect 31666 8191 31722 8200
rect 31217 8186 31223 8188
rect 31279 8186 31303 8188
rect 31359 8186 31383 8188
rect 31439 8186 31463 8188
rect 31519 8186 31525 8188
rect 31279 8134 31281 8186
rect 31461 8134 31463 8186
rect 31217 8132 31223 8134
rect 31279 8132 31303 8134
rect 31359 8132 31383 8134
rect 31439 8132 31463 8134
rect 31519 8132 31525 8134
rect 31217 8123 31525 8132
rect 31217 7100 31525 7109
rect 31217 7098 31223 7100
rect 31279 7098 31303 7100
rect 31359 7098 31383 7100
rect 31439 7098 31463 7100
rect 31519 7098 31525 7100
rect 31279 7046 31281 7098
rect 31461 7046 31463 7098
rect 31217 7044 31223 7046
rect 31279 7044 31303 7046
rect 31359 7044 31383 7046
rect 31439 7044 31463 7046
rect 31519 7044 31525 7046
rect 31217 7035 31525 7044
rect 31217 6012 31525 6021
rect 31217 6010 31223 6012
rect 31279 6010 31303 6012
rect 31359 6010 31383 6012
rect 31439 6010 31463 6012
rect 31519 6010 31525 6012
rect 31279 5958 31281 6010
rect 31461 5958 31463 6010
rect 31217 5956 31223 5958
rect 31279 5956 31303 5958
rect 31359 5956 31383 5958
rect 31439 5956 31463 5958
rect 31519 5956 31525 5958
rect 31217 5947 31525 5956
rect 28446 5536 28502 5545
rect 20456 5506 20668 5534
rect 21744 5506 21956 5534
rect 20640 400 20668 5506
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21284 400 21312 4966
rect 21928 400 21956 5506
rect 27365 5468 27673 5477
rect 28446 5471 28502 5480
rect 27365 5466 27371 5468
rect 27427 5466 27451 5468
rect 27507 5466 27531 5468
rect 27587 5466 27611 5468
rect 27667 5466 27673 5468
rect 27427 5414 27429 5466
rect 27609 5414 27611 5466
rect 27365 5412 27371 5414
rect 27427 5412 27451 5414
rect 27507 5412 27531 5414
rect 27587 5412 27611 5414
rect 27667 5412 27673 5414
rect 27365 5403 27673 5412
rect 23512 4924 23820 4933
rect 23512 4922 23518 4924
rect 23574 4922 23598 4924
rect 23654 4922 23678 4924
rect 23734 4922 23758 4924
rect 23814 4922 23820 4924
rect 23574 4870 23576 4922
rect 23756 4870 23758 4922
rect 23512 4868 23518 4870
rect 23574 4868 23598 4870
rect 23654 4868 23678 4870
rect 23734 4868 23758 4870
rect 23814 4868 23820 4870
rect 23512 4859 23820 4868
rect 31217 4924 31525 4933
rect 31217 4922 31223 4924
rect 31279 4922 31303 4924
rect 31359 4922 31383 4924
rect 31439 4922 31463 4924
rect 31519 4922 31525 4924
rect 31279 4870 31281 4922
rect 31461 4870 31463 4922
rect 31217 4868 31223 4870
rect 31279 4868 31303 4870
rect 31359 4868 31383 4870
rect 31439 4868 31463 4870
rect 31519 4868 31525 4870
rect 31217 4859 31525 4868
rect 27365 4380 27673 4389
rect 27365 4378 27371 4380
rect 27427 4378 27451 4380
rect 27507 4378 27531 4380
rect 27587 4378 27611 4380
rect 27667 4378 27673 4380
rect 27427 4326 27429 4378
rect 27609 4326 27611 4378
rect 27365 4324 27371 4326
rect 27427 4324 27451 4326
rect 27507 4324 27531 4326
rect 27587 4324 27611 4326
rect 27667 4324 27673 4326
rect 27365 4315 27673 4324
rect 23512 3836 23820 3845
rect 23512 3834 23518 3836
rect 23574 3834 23598 3836
rect 23654 3834 23678 3836
rect 23734 3834 23758 3836
rect 23814 3834 23820 3836
rect 23574 3782 23576 3834
rect 23756 3782 23758 3834
rect 23512 3780 23518 3782
rect 23574 3780 23598 3782
rect 23654 3780 23678 3782
rect 23734 3780 23758 3782
rect 23814 3780 23820 3782
rect 23512 3771 23820 3780
rect 31217 3836 31525 3845
rect 31217 3834 31223 3836
rect 31279 3834 31303 3836
rect 31359 3834 31383 3836
rect 31439 3834 31463 3836
rect 31519 3834 31525 3836
rect 31279 3782 31281 3834
rect 31461 3782 31463 3834
rect 31217 3780 31223 3782
rect 31279 3780 31303 3782
rect 31359 3780 31383 3782
rect 31439 3780 31463 3782
rect 31519 3780 31525 3782
rect 31217 3771 31525 3780
rect 27365 3292 27673 3301
rect 27365 3290 27371 3292
rect 27427 3290 27451 3292
rect 27507 3290 27531 3292
rect 27587 3290 27611 3292
rect 27667 3290 27673 3292
rect 27427 3238 27429 3290
rect 27609 3238 27611 3290
rect 27365 3236 27371 3238
rect 27427 3236 27451 3238
rect 27507 3236 27531 3238
rect 27587 3236 27611 3238
rect 27667 3236 27673 3238
rect 27365 3227 27673 3236
rect 23512 2748 23820 2757
rect 23512 2746 23518 2748
rect 23574 2746 23598 2748
rect 23654 2746 23678 2748
rect 23734 2746 23758 2748
rect 23814 2746 23820 2748
rect 23574 2694 23576 2746
rect 23756 2694 23758 2746
rect 23512 2692 23518 2694
rect 23574 2692 23598 2694
rect 23654 2692 23678 2694
rect 23734 2692 23758 2694
rect 23814 2692 23820 2694
rect 23512 2683 23820 2692
rect 31217 2748 31525 2757
rect 31217 2746 31223 2748
rect 31279 2746 31303 2748
rect 31359 2746 31383 2748
rect 31439 2746 31463 2748
rect 31519 2746 31525 2748
rect 31279 2694 31281 2746
rect 31461 2694 31463 2746
rect 31217 2692 31223 2694
rect 31279 2692 31303 2694
rect 31359 2692 31383 2694
rect 31439 2692 31463 2694
rect 31519 2692 31525 2694
rect 31217 2683 31525 2692
rect 27365 2204 27673 2213
rect 27365 2202 27371 2204
rect 27427 2202 27451 2204
rect 27507 2202 27531 2204
rect 27587 2202 27611 2204
rect 27667 2202 27673 2204
rect 27427 2150 27429 2202
rect 27609 2150 27611 2202
rect 27365 2148 27371 2150
rect 27427 2148 27451 2150
rect 27507 2148 27531 2150
rect 27587 2148 27611 2150
rect 27667 2148 27673 2150
rect 27365 2139 27673 2148
rect 23512 1660 23820 1669
rect 23512 1658 23518 1660
rect 23574 1658 23598 1660
rect 23654 1658 23678 1660
rect 23734 1658 23758 1660
rect 23814 1658 23820 1660
rect 23574 1606 23576 1658
rect 23756 1606 23758 1658
rect 23512 1604 23518 1606
rect 23574 1604 23598 1606
rect 23654 1604 23678 1606
rect 23734 1604 23758 1606
rect 23814 1604 23820 1606
rect 23512 1595 23820 1604
rect 31217 1660 31525 1669
rect 31217 1658 31223 1660
rect 31279 1658 31303 1660
rect 31359 1658 31383 1660
rect 31439 1658 31463 1660
rect 31519 1658 31525 1660
rect 31279 1606 31281 1658
rect 31461 1606 31463 1658
rect 31217 1604 31223 1606
rect 31279 1604 31303 1606
rect 31359 1604 31383 1606
rect 31439 1604 31463 1606
rect 31519 1604 31525 1606
rect 31217 1595 31525 1604
rect 27365 1116 27673 1125
rect 27365 1114 27371 1116
rect 27427 1114 27451 1116
rect 27507 1114 27531 1116
rect 27587 1114 27611 1116
rect 27667 1114 27673 1116
rect 27427 1062 27429 1114
rect 27609 1062 27611 1114
rect 27365 1060 27371 1062
rect 27427 1060 27451 1062
rect 27507 1060 27531 1062
rect 27587 1060 27611 1062
rect 27667 1060 27673 1062
rect 27365 1051 27673 1060
rect 22652 808 22704 814
rect 22652 750 22704 756
rect 22664 490 22692 750
rect 23512 572 23820 581
rect 23512 570 23518 572
rect 23574 570 23598 572
rect 23654 570 23678 572
rect 23734 570 23758 572
rect 23814 570 23820 572
rect 23574 518 23576 570
rect 23756 518 23758 570
rect 23512 516 23518 518
rect 23574 516 23598 518
rect 23654 516 23678 518
rect 23734 516 23758 518
rect 23814 516 23820 518
rect 23512 507 23820 516
rect 31217 572 31525 581
rect 31217 570 31223 572
rect 31279 570 31303 572
rect 31359 570 31383 572
rect 31439 570 31463 572
rect 31519 570 31525 572
rect 31279 518 31281 570
rect 31461 518 31463 570
rect 31217 516 31223 518
rect 31279 516 31303 518
rect 31359 516 31383 518
rect 31439 516 31463 518
rect 31519 516 31525 518
rect 31217 507 31525 516
rect 22572 462 22692 490
rect 22572 400 22600 462
rect 7102 0 7158 400
rect 9034 0 9090 400
rect 9678 0 9734 400
rect 10322 0 10378 400
rect 10966 0 11022 400
rect 11610 0 11666 400
rect 12254 0 12310 400
rect 12898 0 12954 400
rect 13542 0 13598 400
rect 14186 0 14242 400
rect 14830 0 14886 400
rect 15474 0 15530 400
rect 16118 0 16174 400
rect 16762 0 16818 400
rect 17406 0 17462 400
rect 18050 0 18106 400
rect 18694 0 18750 400
rect 19338 0 19394 400
rect 19982 0 20038 400
rect 20626 0 20682 400
rect 21270 0 21326 400
rect 21914 0 21970 400
rect 22558 0 22614 400
<< via2 >>
rect 8108 19066 8164 19068
rect 8188 19066 8244 19068
rect 8268 19066 8324 19068
rect 8348 19066 8404 19068
rect 8108 19014 8154 19066
rect 8154 19014 8164 19066
rect 8188 19014 8218 19066
rect 8218 19014 8230 19066
rect 8230 19014 8244 19066
rect 8268 19014 8282 19066
rect 8282 19014 8294 19066
rect 8294 19014 8324 19066
rect 8348 19014 8358 19066
rect 8358 19014 8404 19066
rect 8108 19012 8164 19014
rect 8188 19012 8244 19014
rect 8268 19012 8324 19014
rect 8348 19012 8404 19014
rect 4256 18522 4312 18524
rect 4336 18522 4392 18524
rect 4416 18522 4472 18524
rect 4496 18522 4552 18524
rect 4256 18470 4302 18522
rect 4302 18470 4312 18522
rect 4336 18470 4366 18522
rect 4366 18470 4378 18522
rect 4378 18470 4392 18522
rect 4416 18470 4430 18522
rect 4430 18470 4442 18522
rect 4442 18470 4472 18522
rect 4496 18470 4506 18522
rect 4506 18470 4552 18522
rect 4256 18468 4312 18470
rect 4336 18468 4392 18470
rect 4416 18468 4472 18470
rect 4496 18468 4552 18470
rect 8108 17978 8164 17980
rect 8188 17978 8244 17980
rect 8268 17978 8324 17980
rect 8348 17978 8404 17980
rect 8108 17926 8154 17978
rect 8154 17926 8164 17978
rect 8188 17926 8218 17978
rect 8218 17926 8230 17978
rect 8230 17926 8244 17978
rect 8268 17926 8282 17978
rect 8282 17926 8294 17978
rect 8294 17926 8324 17978
rect 8348 17926 8358 17978
rect 8358 17926 8404 17978
rect 8108 17924 8164 17926
rect 8188 17924 8244 17926
rect 8268 17924 8324 17926
rect 8348 17924 8404 17926
rect 4256 17434 4312 17436
rect 4336 17434 4392 17436
rect 4416 17434 4472 17436
rect 4496 17434 4552 17436
rect 4256 17382 4302 17434
rect 4302 17382 4312 17434
rect 4336 17382 4366 17434
rect 4366 17382 4378 17434
rect 4378 17382 4392 17434
rect 4416 17382 4430 17434
rect 4430 17382 4442 17434
rect 4442 17382 4472 17434
rect 4496 17382 4506 17434
rect 4506 17382 4552 17434
rect 4256 17380 4312 17382
rect 4336 17380 4392 17382
rect 4416 17380 4472 17382
rect 4496 17380 4552 17382
rect 8108 16890 8164 16892
rect 8188 16890 8244 16892
rect 8268 16890 8324 16892
rect 8348 16890 8404 16892
rect 8108 16838 8154 16890
rect 8154 16838 8164 16890
rect 8188 16838 8218 16890
rect 8218 16838 8230 16890
rect 8230 16838 8244 16890
rect 8268 16838 8282 16890
rect 8282 16838 8294 16890
rect 8294 16838 8324 16890
rect 8348 16838 8358 16890
rect 8358 16838 8404 16890
rect 8108 16836 8164 16838
rect 8188 16836 8244 16838
rect 8268 16836 8324 16838
rect 8348 16836 8404 16838
rect 4256 16346 4312 16348
rect 4336 16346 4392 16348
rect 4416 16346 4472 16348
rect 4496 16346 4552 16348
rect 4256 16294 4302 16346
rect 4302 16294 4312 16346
rect 4336 16294 4366 16346
rect 4366 16294 4378 16346
rect 4378 16294 4392 16346
rect 4416 16294 4430 16346
rect 4430 16294 4442 16346
rect 4442 16294 4472 16346
rect 4496 16294 4506 16346
rect 4506 16294 4552 16346
rect 4256 16292 4312 16294
rect 4336 16292 4392 16294
rect 4416 16292 4472 16294
rect 4496 16292 4552 16294
rect 8108 15802 8164 15804
rect 8188 15802 8244 15804
rect 8268 15802 8324 15804
rect 8348 15802 8404 15804
rect 8108 15750 8154 15802
rect 8154 15750 8164 15802
rect 8188 15750 8218 15802
rect 8218 15750 8230 15802
rect 8230 15750 8244 15802
rect 8268 15750 8282 15802
rect 8282 15750 8294 15802
rect 8294 15750 8324 15802
rect 8348 15750 8358 15802
rect 8358 15750 8404 15802
rect 8108 15748 8164 15750
rect 8188 15748 8244 15750
rect 8268 15748 8324 15750
rect 8348 15748 8404 15750
rect 4256 15258 4312 15260
rect 4336 15258 4392 15260
rect 4416 15258 4472 15260
rect 4496 15258 4552 15260
rect 4256 15206 4302 15258
rect 4302 15206 4312 15258
rect 4336 15206 4366 15258
rect 4366 15206 4378 15258
rect 4378 15206 4392 15258
rect 4416 15206 4430 15258
rect 4430 15206 4442 15258
rect 4442 15206 4472 15258
rect 4496 15206 4506 15258
rect 4506 15206 4552 15258
rect 4256 15204 4312 15206
rect 4336 15204 4392 15206
rect 4416 15204 4472 15206
rect 4496 15204 4552 15206
rect 8108 14714 8164 14716
rect 8188 14714 8244 14716
rect 8268 14714 8324 14716
rect 8348 14714 8404 14716
rect 8108 14662 8154 14714
rect 8154 14662 8164 14714
rect 8188 14662 8218 14714
rect 8218 14662 8230 14714
rect 8230 14662 8244 14714
rect 8268 14662 8282 14714
rect 8282 14662 8294 14714
rect 8294 14662 8324 14714
rect 8348 14662 8358 14714
rect 8358 14662 8404 14714
rect 8108 14660 8164 14662
rect 8188 14660 8244 14662
rect 8268 14660 8324 14662
rect 8348 14660 8404 14662
rect 4256 14170 4312 14172
rect 4336 14170 4392 14172
rect 4416 14170 4472 14172
rect 4496 14170 4552 14172
rect 4256 14118 4302 14170
rect 4302 14118 4312 14170
rect 4336 14118 4366 14170
rect 4366 14118 4378 14170
rect 4378 14118 4392 14170
rect 4416 14118 4430 14170
rect 4430 14118 4442 14170
rect 4442 14118 4472 14170
rect 4496 14118 4506 14170
rect 4506 14118 4552 14170
rect 4256 14116 4312 14118
rect 4336 14116 4392 14118
rect 4416 14116 4472 14118
rect 4496 14116 4552 14118
rect 8108 13626 8164 13628
rect 8188 13626 8244 13628
rect 8268 13626 8324 13628
rect 8348 13626 8404 13628
rect 8108 13574 8154 13626
rect 8154 13574 8164 13626
rect 8188 13574 8218 13626
rect 8218 13574 8230 13626
rect 8230 13574 8244 13626
rect 8268 13574 8282 13626
rect 8282 13574 8294 13626
rect 8294 13574 8324 13626
rect 8348 13574 8358 13626
rect 8358 13574 8404 13626
rect 8108 13572 8164 13574
rect 8188 13572 8244 13574
rect 8268 13572 8324 13574
rect 8348 13572 8404 13574
rect 4256 13082 4312 13084
rect 4336 13082 4392 13084
rect 4416 13082 4472 13084
rect 4496 13082 4552 13084
rect 4256 13030 4302 13082
rect 4302 13030 4312 13082
rect 4336 13030 4366 13082
rect 4366 13030 4378 13082
rect 4378 13030 4392 13082
rect 4416 13030 4430 13082
rect 4430 13030 4442 13082
rect 4442 13030 4472 13082
rect 4496 13030 4506 13082
rect 4506 13030 4552 13082
rect 4256 13028 4312 13030
rect 4336 13028 4392 13030
rect 4416 13028 4472 13030
rect 4496 13028 4552 13030
rect 8108 12538 8164 12540
rect 8188 12538 8244 12540
rect 8268 12538 8324 12540
rect 8348 12538 8404 12540
rect 8108 12486 8154 12538
rect 8154 12486 8164 12538
rect 8188 12486 8218 12538
rect 8218 12486 8230 12538
rect 8230 12486 8244 12538
rect 8268 12486 8282 12538
rect 8282 12486 8294 12538
rect 8294 12486 8324 12538
rect 8348 12486 8358 12538
rect 8358 12486 8404 12538
rect 8108 12484 8164 12486
rect 8188 12484 8244 12486
rect 8268 12484 8324 12486
rect 8348 12484 8404 12486
rect 6918 12280 6974 12336
rect 4256 11994 4312 11996
rect 4336 11994 4392 11996
rect 4416 11994 4472 11996
rect 4496 11994 4552 11996
rect 4256 11942 4302 11994
rect 4302 11942 4312 11994
rect 4336 11942 4366 11994
rect 4366 11942 4378 11994
rect 4378 11942 4392 11994
rect 4416 11942 4430 11994
rect 4430 11942 4442 11994
rect 4442 11942 4472 11994
rect 4496 11942 4506 11994
rect 4506 11942 4552 11994
rect 4256 11940 4312 11942
rect 4336 11940 4392 11942
rect 4416 11940 4472 11942
rect 4496 11940 4552 11942
rect 6918 11600 6974 11656
rect 8108 11450 8164 11452
rect 8188 11450 8244 11452
rect 8268 11450 8324 11452
rect 8348 11450 8404 11452
rect 8108 11398 8154 11450
rect 8154 11398 8164 11450
rect 8188 11398 8218 11450
rect 8218 11398 8230 11450
rect 8230 11398 8244 11450
rect 8268 11398 8282 11450
rect 8282 11398 8294 11450
rect 8294 11398 8324 11450
rect 8348 11398 8358 11450
rect 8358 11398 8404 11450
rect 8108 11396 8164 11398
rect 8188 11396 8244 11398
rect 8268 11396 8324 11398
rect 8348 11396 8404 11398
rect 4256 10906 4312 10908
rect 4336 10906 4392 10908
rect 4416 10906 4472 10908
rect 4496 10906 4552 10908
rect 4256 10854 4302 10906
rect 4302 10854 4312 10906
rect 4336 10854 4366 10906
rect 4366 10854 4378 10906
rect 4378 10854 4392 10906
rect 4416 10854 4430 10906
rect 4430 10854 4442 10906
rect 4442 10854 4472 10906
rect 4496 10854 4506 10906
rect 4506 10854 4552 10906
rect 4256 10852 4312 10854
rect 4336 10852 4392 10854
rect 4416 10852 4472 10854
rect 4496 10852 4552 10854
rect 8108 10362 8164 10364
rect 8188 10362 8244 10364
rect 8268 10362 8324 10364
rect 8348 10362 8404 10364
rect 8108 10310 8154 10362
rect 8154 10310 8164 10362
rect 8188 10310 8218 10362
rect 8218 10310 8230 10362
rect 8230 10310 8244 10362
rect 8268 10310 8282 10362
rect 8282 10310 8294 10362
rect 8294 10310 8324 10362
rect 8348 10310 8358 10362
rect 8358 10310 8404 10362
rect 8108 10308 8164 10310
rect 8188 10308 8244 10310
rect 8268 10308 8324 10310
rect 8348 10308 8404 10310
rect 7102 10260 7158 10296
rect 7102 10240 7104 10260
rect 7104 10240 7156 10260
rect 7156 10240 7158 10260
rect 4256 9818 4312 9820
rect 4336 9818 4392 9820
rect 4416 9818 4472 9820
rect 4496 9818 4552 9820
rect 4256 9766 4302 9818
rect 4302 9766 4312 9818
rect 4336 9766 4366 9818
rect 4366 9766 4378 9818
rect 4378 9766 4392 9818
rect 4416 9766 4430 9818
rect 4430 9766 4442 9818
rect 4442 9766 4472 9818
rect 4496 9766 4506 9818
rect 4506 9766 4552 9818
rect 4256 9764 4312 9766
rect 4336 9764 4392 9766
rect 4416 9764 4472 9766
rect 4496 9764 4552 9766
rect 6734 8900 6790 8936
rect 6734 8880 6736 8900
rect 6736 8880 6788 8900
rect 6788 8880 6790 8900
rect 4256 8730 4312 8732
rect 4336 8730 4392 8732
rect 4416 8730 4472 8732
rect 4496 8730 4552 8732
rect 4256 8678 4302 8730
rect 4302 8678 4312 8730
rect 4336 8678 4366 8730
rect 4366 8678 4378 8730
rect 4378 8678 4392 8730
rect 4416 8678 4430 8730
rect 4430 8678 4442 8730
rect 4442 8678 4472 8730
rect 4496 8678 4506 8730
rect 4506 8678 4552 8730
rect 4256 8676 4312 8678
rect 4336 8676 4392 8678
rect 4416 8676 4472 8678
rect 4496 8676 4552 8678
rect 4256 7642 4312 7644
rect 4336 7642 4392 7644
rect 4416 7642 4472 7644
rect 4496 7642 4552 7644
rect 4256 7590 4302 7642
rect 4302 7590 4312 7642
rect 4336 7590 4366 7642
rect 4366 7590 4378 7642
rect 4378 7590 4392 7642
rect 4416 7590 4430 7642
rect 4430 7590 4442 7642
rect 4442 7590 4472 7642
rect 4496 7590 4506 7642
rect 4506 7590 4552 7642
rect 4256 7588 4312 7590
rect 4336 7588 4392 7590
rect 4416 7588 4472 7590
rect 4496 7588 4552 7590
rect 6642 6840 6698 6896
rect 4256 6554 4312 6556
rect 4336 6554 4392 6556
rect 4416 6554 4472 6556
rect 4496 6554 4552 6556
rect 4256 6502 4302 6554
rect 4302 6502 4312 6554
rect 4336 6502 4366 6554
rect 4366 6502 4378 6554
rect 4378 6502 4392 6554
rect 4416 6502 4430 6554
rect 4430 6502 4442 6554
rect 4442 6502 4472 6554
rect 4496 6502 4506 6554
rect 4506 6502 4552 6554
rect 4256 6500 4312 6502
rect 4336 6500 4392 6502
rect 4416 6500 4472 6502
rect 4496 6500 4552 6502
rect 4256 5466 4312 5468
rect 4336 5466 4392 5468
rect 4416 5466 4472 5468
rect 4496 5466 4552 5468
rect 4256 5414 4302 5466
rect 4302 5414 4312 5466
rect 4336 5414 4366 5466
rect 4366 5414 4378 5466
rect 4378 5414 4392 5466
rect 4416 5414 4430 5466
rect 4430 5414 4442 5466
rect 4442 5414 4472 5466
rect 4496 5414 4506 5466
rect 4506 5414 4552 5466
rect 4256 5412 4312 5414
rect 4336 5412 4392 5414
rect 4416 5412 4472 5414
rect 4496 5412 4552 5414
rect 4256 4378 4312 4380
rect 4336 4378 4392 4380
rect 4416 4378 4472 4380
rect 4496 4378 4552 4380
rect 4256 4326 4302 4378
rect 4302 4326 4312 4378
rect 4336 4326 4366 4378
rect 4366 4326 4378 4378
rect 4378 4326 4392 4378
rect 4416 4326 4430 4378
rect 4430 4326 4442 4378
rect 4442 4326 4472 4378
rect 4496 4326 4506 4378
rect 4506 4326 4552 4378
rect 4256 4324 4312 4326
rect 4336 4324 4392 4326
rect 4416 4324 4472 4326
rect 4496 4324 4552 4326
rect 4256 3290 4312 3292
rect 4336 3290 4392 3292
rect 4416 3290 4472 3292
rect 4496 3290 4552 3292
rect 4256 3238 4302 3290
rect 4302 3238 4312 3290
rect 4336 3238 4366 3290
rect 4366 3238 4378 3290
rect 4378 3238 4392 3290
rect 4416 3238 4430 3290
rect 4430 3238 4442 3290
rect 4442 3238 4472 3290
rect 4496 3238 4506 3290
rect 4506 3238 4552 3290
rect 4256 3236 4312 3238
rect 4336 3236 4392 3238
rect 4416 3236 4472 3238
rect 4496 3236 4552 3238
rect 9770 9596 9772 9616
rect 9772 9596 9824 9616
rect 9824 9596 9826 9616
rect 9770 9560 9826 9596
rect 8108 9274 8164 9276
rect 8188 9274 8244 9276
rect 8268 9274 8324 9276
rect 8348 9274 8404 9276
rect 8108 9222 8154 9274
rect 8154 9222 8164 9274
rect 8188 9222 8218 9274
rect 8218 9222 8230 9274
rect 8230 9222 8244 9274
rect 8268 9222 8282 9274
rect 8282 9222 8294 9274
rect 8294 9222 8324 9274
rect 8348 9222 8358 9274
rect 8358 9222 8404 9274
rect 8108 9220 8164 9222
rect 8188 9220 8244 9222
rect 8268 9220 8324 9222
rect 8348 9220 8404 9222
rect 8108 8186 8164 8188
rect 8188 8186 8244 8188
rect 8268 8186 8324 8188
rect 8348 8186 8404 8188
rect 8108 8134 8154 8186
rect 8154 8134 8164 8186
rect 8188 8134 8218 8186
rect 8218 8134 8230 8186
rect 8230 8134 8244 8186
rect 8268 8134 8282 8186
rect 8282 8134 8294 8186
rect 8294 8134 8324 8186
rect 8348 8134 8358 8186
rect 8358 8134 8404 8186
rect 8108 8132 8164 8134
rect 8188 8132 8244 8134
rect 8268 8132 8324 8134
rect 8348 8132 8404 8134
rect 9402 7928 9458 7984
rect 9310 7792 9366 7848
rect 11961 18522 12017 18524
rect 12041 18522 12097 18524
rect 12121 18522 12177 18524
rect 12201 18522 12257 18524
rect 11961 18470 12007 18522
rect 12007 18470 12017 18522
rect 12041 18470 12071 18522
rect 12071 18470 12083 18522
rect 12083 18470 12097 18522
rect 12121 18470 12135 18522
rect 12135 18470 12147 18522
rect 12147 18470 12177 18522
rect 12201 18470 12211 18522
rect 12211 18470 12257 18522
rect 11961 18468 12017 18470
rect 12041 18468 12097 18470
rect 12121 18468 12177 18470
rect 12201 18468 12257 18470
rect 11961 17434 12017 17436
rect 12041 17434 12097 17436
rect 12121 17434 12177 17436
rect 12201 17434 12257 17436
rect 11961 17382 12007 17434
rect 12007 17382 12017 17434
rect 12041 17382 12071 17434
rect 12071 17382 12083 17434
rect 12083 17382 12097 17434
rect 12121 17382 12135 17434
rect 12135 17382 12147 17434
rect 12147 17382 12177 17434
rect 12201 17382 12211 17434
rect 12211 17382 12257 17434
rect 11961 17380 12017 17382
rect 12041 17380 12097 17382
rect 12121 17380 12177 17382
rect 12201 17380 12257 17382
rect 11961 16346 12017 16348
rect 12041 16346 12097 16348
rect 12121 16346 12177 16348
rect 12201 16346 12257 16348
rect 11961 16294 12007 16346
rect 12007 16294 12017 16346
rect 12041 16294 12071 16346
rect 12071 16294 12083 16346
rect 12083 16294 12097 16346
rect 12121 16294 12135 16346
rect 12135 16294 12147 16346
rect 12147 16294 12177 16346
rect 12201 16294 12211 16346
rect 12211 16294 12257 16346
rect 11961 16292 12017 16294
rect 12041 16292 12097 16294
rect 12121 16292 12177 16294
rect 12201 16292 12257 16294
rect 11961 15258 12017 15260
rect 12041 15258 12097 15260
rect 12121 15258 12177 15260
rect 12201 15258 12257 15260
rect 11961 15206 12007 15258
rect 12007 15206 12017 15258
rect 12041 15206 12071 15258
rect 12071 15206 12083 15258
rect 12083 15206 12097 15258
rect 12121 15206 12135 15258
rect 12135 15206 12147 15258
rect 12147 15206 12177 15258
rect 12201 15206 12211 15258
rect 12211 15206 12257 15258
rect 11961 15204 12017 15206
rect 12041 15204 12097 15206
rect 12121 15204 12177 15206
rect 12201 15204 12257 15206
rect 11961 14170 12017 14172
rect 12041 14170 12097 14172
rect 12121 14170 12177 14172
rect 12201 14170 12257 14172
rect 11961 14118 12007 14170
rect 12007 14118 12017 14170
rect 12041 14118 12071 14170
rect 12071 14118 12083 14170
rect 12083 14118 12097 14170
rect 12121 14118 12135 14170
rect 12135 14118 12147 14170
rect 12147 14118 12177 14170
rect 12201 14118 12211 14170
rect 12211 14118 12257 14170
rect 11961 14116 12017 14118
rect 12041 14116 12097 14118
rect 12121 14116 12177 14118
rect 12201 14116 12257 14118
rect 11961 13082 12017 13084
rect 12041 13082 12097 13084
rect 12121 13082 12177 13084
rect 12201 13082 12257 13084
rect 11961 13030 12007 13082
rect 12007 13030 12017 13082
rect 12041 13030 12071 13082
rect 12071 13030 12083 13082
rect 12083 13030 12097 13082
rect 12121 13030 12135 13082
rect 12135 13030 12147 13082
rect 12147 13030 12177 13082
rect 12201 13030 12211 13082
rect 12211 13030 12257 13082
rect 11961 13028 12017 13030
rect 12041 13028 12097 13030
rect 12121 13028 12177 13030
rect 12201 13028 12257 13030
rect 11961 11994 12017 11996
rect 12041 11994 12097 11996
rect 12121 11994 12177 11996
rect 12201 11994 12257 11996
rect 11961 11942 12007 11994
rect 12007 11942 12017 11994
rect 12041 11942 12071 11994
rect 12071 11942 12083 11994
rect 12083 11942 12097 11994
rect 12121 11942 12135 11994
rect 12135 11942 12147 11994
rect 12147 11942 12177 11994
rect 12201 11942 12211 11994
rect 12211 11942 12257 11994
rect 11961 11940 12017 11942
rect 12041 11940 12097 11942
rect 12121 11940 12177 11942
rect 12201 11940 12257 11942
rect 15813 19066 15869 19068
rect 15893 19066 15949 19068
rect 15973 19066 16029 19068
rect 16053 19066 16109 19068
rect 15813 19014 15859 19066
rect 15859 19014 15869 19066
rect 15893 19014 15923 19066
rect 15923 19014 15935 19066
rect 15935 19014 15949 19066
rect 15973 19014 15987 19066
rect 15987 19014 15999 19066
rect 15999 19014 16029 19066
rect 16053 19014 16063 19066
rect 16063 19014 16109 19066
rect 15813 19012 15869 19014
rect 15893 19012 15949 19014
rect 15973 19012 16029 19014
rect 16053 19012 16109 19014
rect 15813 17978 15869 17980
rect 15893 17978 15949 17980
rect 15973 17978 16029 17980
rect 16053 17978 16109 17980
rect 15813 17926 15859 17978
rect 15859 17926 15869 17978
rect 15893 17926 15923 17978
rect 15923 17926 15935 17978
rect 15935 17926 15949 17978
rect 15973 17926 15987 17978
rect 15987 17926 15999 17978
rect 15999 17926 16029 17978
rect 16053 17926 16063 17978
rect 16063 17926 16109 17978
rect 15813 17924 15869 17926
rect 15893 17924 15949 17926
rect 15973 17924 16029 17926
rect 16053 17924 16109 17926
rect 15813 16890 15869 16892
rect 15893 16890 15949 16892
rect 15973 16890 16029 16892
rect 16053 16890 16109 16892
rect 15813 16838 15859 16890
rect 15859 16838 15869 16890
rect 15893 16838 15923 16890
rect 15923 16838 15935 16890
rect 15935 16838 15949 16890
rect 15973 16838 15987 16890
rect 15987 16838 15999 16890
rect 15999 16838 16029 16890
rect 16053 16838 16063 16890
rect 16063 16838 16109 16890
rect 15813 16836 15869 16838
rect 15893 16836 15949 16838
rect 15973 16836 16029 16838
rect 16053 16836 16109 16838
rect 15813 15802 15869 15804
rect 15893 15802 15949 15804
rect 15973 15802 16029 15804
rect 16053 15802 16109 15804
rect 15813 15750 15859 15802
rect 15859 15750 15869 15802
rect 15893 15750 15923 15802
rect 15923 15750 15935 15802
rect 15935 15750 15949 15802
rect 15973 15750 15987 15802
rect 15987 15750 15999 15802
rect 15999 15750 16029 15802
rect 16053 15750 16063 15802
rect 16063 15750 16109 15802
rect 15813 15748 15869 15750
rect 15893 15748 15949 15750
rect 15973 15748 16029 15750
rect 16053 15748 16109 15750
rect 15813 14714 15869 14716
rect 15893 14714 15949 14716
rect 15973 14714 16029 14716
rect 16053 14714 16109 14716
rect 15813 14662 15859 14714
rect 15859 14662 15869 14714
rect 15893 14662 15923 14714
rect 15923 14662 15935 14714
rect 15935 14662 15949 14714
rect 15973 14662 15987 14714
rect 15987 14662 15999 14714
rect 15999 14662 16029 14714
rect 16053 14662 16063 14714
rect 16063 14662 16109 14714
rect 15813 14660 15869 14662
rect 15893 14660 15949 14662
rect 15973 14660 16029 14662
rect 16053 14660 16109 14662
rect 15813 13626 15869 13628
rect 15893 13626 15949 13628
rect 15973 13626 16029 13628
rect 16053 13626 16109 13628
rect 15813 13574 15859 13626
rect 15859 13574 15869 13626
rect 15893 13574 15923 13626
rect 15923 13574 15935 13626
rect 15935 13574 15949 13626
rect 15973 13574 15987 13626
rect 15987 13574 15999 13626
rect 15999 13574 16029 13626
rect 16053 13574 16063 13626
rect 16063 13574 16109 13626
rect 15813 13572 15869 13574
rect 15893 13572 15949 13574
rect 15973 13572 16029 13574
rect 16053 13572 16109 13574
rect 15813 12538 15869 12540
rect 15893 12538 15949 12540
rect 15973 12538 16029 12540
rect 16053 12538 16109 12540
rect 15813 12486 15859 12538
rect 15859 12486 15869 12538
rect 15893 12486 15923 12538
rect 15923 12486 15935 12538
rect 15935 12486 15949 12538
rect 15973 12486 15987 12538
rect 15987 12486 15999 12538
rect 15999 12486 16029 12538
rect 16053 12486 16063 12538
rect 16063 12486 16109 12538
rect 15813 12484 15869 12486
rect 15893 12484 15949 12486
rect 15973 12484 16029 12486
rect 16053 12484 16109 12486
rect 15813 11450 15869 11452
rect 15893 11450 15949 11452
rect 15973 11450 16029 11452
rect 16053 11450 16109 11452
rect 15813 11398 15859 11450
rect 15859 11398 15869 11450
rect 15893 11398 15923 11450
rect 15923 11398 15935 11450
rect 15935 11398 15949 11450
rect 15973 11398 15987 11450
rect 15987 11398 15999 11450
rect 15999 11398 16029 11450
rect 16053 11398 16063 11450
rect 16063 11398 16109 11450
rect 15813 11396 15869 11398
rect 15893 11396 15949 11398
rect 15973 11396 16029 11398
rect 16053 11396 16109 11398
rect 11961 10906 12017 10908
rect 12041 10906 12097 10908
rect 12121 10906 12177 10908
rect 12201 10906 12257 10908
rect 11961 10854 12007 10906
rect 12007 10854 12017 10906
rect 12041 10854 12071 10906
rect 12071 10854 12083 10906
rect 12083 10854 12097 10906
rect 12121 10854 12135 10906
rect 12135 10854 12147 10906
rect 12147 10854 12177 10906
rect 12201 10854 12211 10906
rect 12211 10854 12257 10906
rect 11961 10852 12017 10854
rect 12041 10852 12097 10854
rect 12121 10852 12177 10854
rect 12201 10852 12257 10854
rect 11150 10804 11206 10840
rect 11150 10784 11152 10804
rect 11152 10784 11204 10804
rect 11204 10784 11206 10804
rect 11961 9818 12017 9820
rect 12041 9818 12097 9820
rect 12121 9818 12177 9820
rect 12201 9818 12257 9820
rect 11961 9766 12007 9818
rect 12007 9766 12017 9818
rect 12041 9766 12071 9818
rect 12071 9766 12083 9818
rect 12083 9766 12097 9818
rect 12121 9766 12135 9818
rect 12135 9766 12147 9818
rect 12147 9766 12177 9818
rect 12201 9766 12211 9818
rect 12211 9766 12257 9818
rect 11961 9764 12017 9766
rect 12041 9764 12097 9766
rect 12121 9764 12177 9766
rect 12201 9764 12257 9766
rect 8108 7098 8164 7100
rect 8188 7098 8244 7100
rect 8268 7098 8324 7100
rect 8348 7098 8404 7100
rect 8108 7046 8154 7098
rect 8154 7046 8164 7098
rect 8188 7046 8218 7098
rect 8218 7046 8230 7098
rect 8230 7046 8244 7098
rect 8268 7046 8282 7098
rect 8282 7046 8294 7098
rect 8294 7046 8324 7098
rect 8348 7046 8358 7098
rect 8358 7046 8404 7098
rect 8108 7044 8164 7046
rect 8188 7044 8244 7046
rect 8268 7044 8324 7046
rect 8348 7044 8404 7046
rect 7838 6160 7894 6216
rect 8108 6010 8164 6012
rect 8188 6010 8244 6012
rect 8268 6010 8324 6012
rect 8348 6010 8404 6012
rect 8108 5958 8154 6010
rect 8154 5958 8164 6010
rect 8188 5958 8218 6010
rect 8218 5958 8230 6010
rect 8230 5958 8244 6010
rect 8268 5958 8282 6010
rect 8282 5958 8294 6010
rect 8294 5958 8324 6010
rect 8348 5958 8358 6010
rect 8358 5958 8404 6010
rect 8108 5956 8164 5958
rect 8188 5956 8244 5958
rect 8268 5956 8324 5958
rect 8348 5956 8404 5958
rect 8108 4922 8164 4924
rect 8188 4922 8244 4924
rect 8268 4922 8324 4924
rect 8348 4922 8404 4924
rect 8108 4870 8154 4922
rect 8154 4870 8164 4922
rect 8188 4870 8218 4922
rect 8218 4870 8230 4922
rect 8230 4870 8244 4922
rect 8268 4870 8282 4922
rect 8282 4870 8294 4922
rect 8294 4870 8324 4922
rect 8348 4870 8358 4922
rect 8358 4870 8404 4922
rect 8108 4868 8164 4870
rect 8188 4868 8244 4870
rect 8268 4868 8324 4870
rect 8348 4868 8404 4870
rect 8108 3834 8164 3836
rect 8188 3834 8244 3836
rect 8268 3834 8324 3836
rect 8348 3834 8404 3836
rect 8108 3782 8154 3834
rect 8154 3782 8164 3834
rect 8188 3782 8218 3834
rect 8218 3782 8230 3834
rect 8230 3782 8244 3834
rect 8268 3782 8282 3834
rect 8282 3782 8294 3834
rect 8294 3782 8324 3834
rect 8348 3782 8358 3834
rect 8358 3782 8404 3834
rect 8108 3780 8164 3782
rect 8188 3780 8244 3782
rect 8268 3780 8324 3782
rect 8348 3780 8404 3782
rect 8108 2746 8164 2748
rect 8188 2746 8244 2748
rect 8268 2746 8324 2748
rect 8348 2746 8404 2748
rect 4256 2202 4312 2204
rect 4336 2202 4392 2204
rect 4416 2202 4472 2204
rect 4496 2202 4552 2204
rect 4256 2150 4302 2202
rect 4302 2150 4312 2202
rect 4336 2150 4366 2202
rect 4366 2150 4378 2202
rect 4378 2150 4392 2202
rect 4416 2150 4430 2202
rect 4430 2150 4442 2202
rect 4442 2150 4472 2202
rect 4496 2150 4506 2202
rect 4506 2150 4552 2202
rect 4256 2148 4312 2150
rect 4336 2148 4392 2150
rect 4416 2148 4472 2150
rect 4496 2148 4552 2150
rect 4256 1114 4312 1116
rect 4336 1114 4392 1116
rect 4416 1114 4472 1116
rect 4496 1114 4552 1116
rect 4256 1062 4302 1114
rect 4302 1062 4312 1114
rect 4336 1062 4366 1114
rect 4366 1062 4378 1114
rect 4378 1062 4392 1114
rect 4416 1062 4430 1114
rect 4430 1062 4442 1114
rect 4442 1062 4472 1114
rect 4496 1062 4506 1114
rect 4506 1062 4552 1114
rect 4256 1060 4312 1062
rect 4336 1060 4392 1062
rect 4416 1060 4472 1062
rect 4496 1060 4552 1062
rect 8108 2694 8154 2746
rect 8154 2694 8164 2746
rect 8188 2694 8218 2746
rect 8218 2694 8230 2746
rect 8230 2694 8244 2746
rect 8268 2694 8282 2746
rect 8282 2694 8294 2746
rect 8294 2694 8324 2746
rect 8348 2694 8358 2746
rect 8358 2694 8404 2746
rect 8108 2692 8164 2694
rect 8188 2692 8244 2694
rect 8268 2692 8324 2694
rect 8348 2692 8404 2694
rect 8108 1658 8164 1660
rect 8188 1658 8244 1660
rect 8268 1658 8324 1660
rect 8348 1658 8404 1660
rect 8108 1606 8154 1658
rect 8154 1606 8164 1658
rect 8188 1606 8218 1658
rect 8218 1606 8230 1658
rect 8230 1606 8244 1658
rect 8268 1606 8282 1658
rect 8282 1606 8294 1658
rect 8294 1606 8324 1658
rect 8348 1606 8358 1658
rect 8358 1606 8404 1658
rect 8108 1604 8164 1606
rect 8188 1604 8244 1606
rect 8268 1604 8324 1606
rect 8348 1604 8404 1606
rect 8108 570 8164 572
rect 8188 570 8244 572
rect 8268 570 8324 572
rect 8348 570 8404 572
rect 8108 518 8154 570
rect 8154 518 8164 570
rect 8188 518 8218 570
rect 8218 518 8230 570
rect 8230 518 8244 570
rect 8268 518 8282 570
rect 8282 518 8294 570
rect 8294 518 8324 570
rect 8348 518 8358 570
rect 8358 518 8404 570
rect 8108 516 8164 518
rect 8188 516 8244 518
rect 8268 516 8324 518
rect 8348 516 8404 518
rect 11961 8730 12017 8732
rect 12041 8730 12097 8732
rect 12121 8730 12177 8732
rect 12201 8730 12257 8732
rect 11961 8678 12007 8730
rect 12007 8678 12017 8730
rect 12041 8678 12071 8730
rect 12071 8678 12083 8730
rect 12083 8678 12097 8730
rect 12121 8678 12135 8730
rect 12135 8678 12147 8730
rect 12147 8678 12177 8730
rect 12201 8678 12211 8730
rect 12211 8678 12257 8730
rect 11961 8676 12017 8678
rect 12041 8676 12097 8678
rect 12121 8676 12177 8678
rect 12201 8676 12257 8678
rect 11961 7642 12017 7644
rect 12041 7642 12097 7644
rect 12121 7642 12177 7644
rect 12201 7642 12257 7644
rect 11961 7590 12007 7642
rect 12007 7590 12017 7642
rect 12041 7590 12071 7642
rect 12071 7590 12083 7642
rect 12083 7590 12097 7642
rect 12121 7590 12135 7642
rect 12135 7590 12147 7642
rect 12147 7590 12177 7642
rect 12201 7590 12211 7642
rect 12211 7590 12257 7642
rect 11961 7588 12017 7590
rect 12041 7588 12097 7590
rect 12121 7588 12177 7590
rect 12201 7588 12257 7590
rect 11961 6554 12017 6556
rect 12041 6554 12097 6556
rect 12121 6554 12177 6556
rect 12201 6554 12257 6556
rect 11961 6502 12007 6554
rect 12007 6502 12017 6554
rect 12041 6502 12071 6554
rect 12071 6502 12083 6554
rect 12083 6502 12097 6554
rect 12121 6502 12135 6554
rect 12135 6502 12147 6554
rect 12147 6502 12177 6554
rect 12201 6502 12211 6554
rect 12211 6502 12257 6554
rect 11961 6500 12017 6502
rect 12041 6500 12097 6502
rect 12121 6500 12177 6502
rect 12201 6500 12257 6502
rect 11961 5466 12017 5468
rect 12041 5466 12097 5468
rect 12121 5466 12177 5468
rect 12201 5466 12257 5468
rect 11961 5414 12007 5466
rect 12007 5414 12017 5466
rect 12041 5414 12071 5466
rect 12071 5414 12083 5466
rect 12083 5414 12097 5466
rect 12121 5414 12135 5466
rect 12135 5414 12147 5466
rect 12147 5414 12177 5466
rect 12201 5414 12211 5466
rect 12211 5414 12257 5466
rect 11961 5412 12017 5414
rect 12041 5412 12097 5414
rect 12121 5412 12177 5414
rect 12201 5412 12257 5414
rect 11961 4378 12017 4380
rect 12041 4378 12097 4380
rect 12121 4378 12177 4380
rect 12201 4378 12257 4380
rect 11961 4326 12007 4378
rect 12007 4326 12017 4378
rect 12041 4326 12071 4378
rect 12071 4326 12083 4378
rect 12083 4326 12097 4378
rect 12121 4326 12135 4378
rect 12135 4326 12147 4378
rect 12147 4326 12177 4378
rect 12201 4326 12211 4378
rect 12211 4326 12257 4378
rect 11961 4324 12017 4326
rect 12041 4324 12097 4326
rect 12121 4324 12177 4326
rect 12201 4324 12257 4326
rect 11961 3290 12017 3292
rect 12041 3290 12097 3292
rect 12121 3290 12177 3292
rect 12201 3290 12257 3292
rect 11961 3238 12007 3290
rect 12007 3238 12017 3290
rect 12041 3238 12071 3290
rect 12071 3238 12083 3290
rect 12083 3238 12097 3290
rect 12121 3238 12135 3290
rect 12135 3238 12147 3290
rect 12147 3238 12177 3290
rect 12201 3238 12211 3290
rect 12211 3238 12257 3290
rect 11961 3236 12017 3238
rect 12041 3236 12097 3238
rect 12121 3236 12177 3238
rect 12201 3236 12257 3238
rect 11961 2202 12017 2204
rect 12041 2202 12097 2204
rect 12121 2202 12177 2204
rect 12201 2202 12257 2204
rect 11961 2150 12007 2202
rect 12007 2150 12017 2202
rect 12041 2150 12071 2202
rect 12071 2150 12083 2202
rect 12083 2150 12097 2202
rect 12121 2150 12135 2202
rect 12135 2150 12147 2202
rect 12147 2150 12177 2202
rect 12201 2150 12211 2202
rect 12211 2150 12257 2202
rect 11961 2148 12017 2150
rect 12041 2148 12097 2150
rect 12121 2148 12177 2150
rect 12201 2148 12257 2150
rect 11961 1114 12017 1116
rect 12041 1114 12097 1116
rect 12121 1114 12177 1116
rect 12201 1114 12257 1116
rect 11961 1062 12007 1114
rect 12007 1062 12017 1114
rect 12041 1062 12071 1114
rect 12071 1062 12083 1114
rect 12083 1062 12097 1114
rect 12121 1062 12135 1114
rect 12135 1062 12147 1114
rect 12147 1062 12177 1114
rect 12201 1062 12211 1114
rect 12211 1062 12257 1114
rect 11961 1060 12017 1062
rect 12041 1060 12097 1062
rect 12121 1060 12177 1062
rect 12201 1060 12257 1062
rect 15813 10362 15869 10364
rect 15893 10362 15949 10364
rect 15973 10362 16029 10364
rect 16053 10362 16109 10364
rect 15813 10310 15859 10362
rect 15859 10310 15869 10362
rect 15893 10310 15923 10362
rect 15923 10310 15935 10362
rect 15935 10310 15949 10362
rect 15973 10310 15987 10362
rect 15987 10310 15999 10362
rect 15999 10310 16029 10362
rect 16053 10310 16063 10362
rect 16063 10310 16109 10362
rect 15813 10308 15869 10310
rect 15893 10308 15949 10310
rect 15973 10308 16029 10310
rect 16053 10308 16109 10310
rect 19666 18522 19722 18524
rect 19746 18522 19802 18524
rect 19826 18522 19882 18524
rect 19906 18522 19962 18524
rect 19666 18470 19712 18522
rect 19712 18470 19722 18522
rect 19746 18470 19776 18522
rect 19776 18470 19788 18522
rect 19788 18470 19802 18522
rect 19826 18470 19840 18522
rect 19840 18470 19852 18522
rect 19852 18470 19882 18522
rect 19906 18470 19916 18522
rect 19916 18470 19962 18522
rect 19666 18468 19722 18470
rect 19746 18468 19802 18470
rect 19826 18468 19882 18470
rect 19906 18468 19962 18470
rect 19666 17434 19722 17436
rect 19746 17434 19802 17436
rect 19826 17434 19882 17436
rect 19906 17434 19962 17436
rect 19666 17382 19712 17434
rect 19712 17382 19722 17434
rect 19746 17382 19776 17434
rect 19776 17382 19788 17434
rect 19788 17382 19802 17434
rect 19826 17382 19840 17434
rect 19840 17382 19852 17434
rect 19852 17382 19882 17434
rect 19906 17382 19916 17434
rect 19916 17382 19962 17434
rect 19666 17380 19722 17382
rect 19746 17380 19802 17382
rect 19826 17380 19882 17382
rect 19906 17380 19962 17382
rect 19666 16346 19722 16348
rect 19746 16346 19802 16348
rect 19826 16346 19882 16348
rect 19906 16346 19962 16348
rect 19666 16294 19712 16346
rect 19712 16294 19722 16346
rect 19746 16294 19776 16346
rect 19776 16294 19788 16346
rect 19788 16294 19802 16346
rect 19826 16294 19840 16346
rect 19840 16294 19852 16346
rect 19852 16294 19882 16346
rect 19906 16294 19916 16346
rect 19916 16294 19962 16346
rect 19666 16292 19722 16294
rect 19746 16292 19802 16294
rect 19826 16292 19882 16294
rect 19906 16292 19962 16294
rect 19666 15258 19722 15260
rect 19746 15258 19802 15260
rect 19826 15258 19882 15260
rect 19906 15258 19962 15260
rect 19666 15206 19712 15258
rect 19712 15206 19722 15258
rect 19746 15206 19776 15258
rect 19776 15206 19788 15258
rect 19788 15206 19802 15258
rect 19826 15206 19840 15258
rect 19840 15206 19852 15258
rect 19852 15206 19882 15258
rect 19906 15206 19916 15258
rect 19916 15206 19962 15258
rect 19666 15204 19722 15206
rect 19746 15204 19802 15206
rect 19826 15204 19882 15206
rect 19906 15204 19962 15206
rect 19666 14170 19722 14172
rect 19746 14170 19802 14172
rect 19826 14170 19882 14172
rect 19906 14170 19962 14172
rect 19666 14118 19712 14170
rect 19712 14118 19722 14170
rect 19746 14118 19776 14170
rect 19776 14118 19788 14170
rect 19788 14118 19802 14170
rect 19826 14118 19840 14170
rect 19840 14118 19852 14170
rect 19852 14118 19882 14170
rect 19906 14118 19916 14170
rect 19916 14118 19962 14170
rect 19666 14116 19722 14118
rect 19746 14116 19802 14118
rect 19826 14116 19882 14118
rect 19906 14116 19962 14118
rect 19666 13082 19722 13084
rect 19746 13082 19802 13084
rect 19826 13082 19882 13084
rect 19906 13082 19962 13084
rect 19666 13030 19712 13082
rect 19712 13030 19722 13082
rect 19746 13030 19776 13082
rect 19776 13030 19788 13082
rect 19788 13030 19802 13082
rect 19826 13030 19840 13082
rect 19840 13030 19852 13082
rect 19852 13030 19882 13082
rect 19906 13030 19916 13082
rect 19916 13030 19962 13082
rect 19666 13028 19722 13030
rect 19746 13028 19802 13030
rect 19826 13028 19882 13030
rect 19906 13028 19962 13030
rect 19666 11994 19722 11996
rect 19746 11994 19802 11996
rect 19826 11994 19882 11996
rect 19906 11994 19962 11996
rect 19666 11942 19712 11994
rect 19712 11942 19722 11994
rect 19746 11942 19776 11994
rect 19776 11942 19788 11994
rect 19788 11942 19802 11994
rect 19826 11942 19840 11994
rect 19840 11942 19852 11994
rect 19852 11942 19882 11994
rect 19906 11942 19916 11994
rect 19916 11942 19962 11994
rect 19666 11940 19722 11942
rect 19746 11940 19802 11942
rect 19826 11940 19882 11942
rect 19906 11940 19962 11942
rect 19666 10906 19722 10908
rect 19746 10906 19802 10908
rect 19826 10906 19882 10908
rect 19906 10906 19962 10908
rect 19666 10854 19712 10906
rect 19712 10854 19722 10906
rect 19746 10854 19776 10906
rect 19776 10854 19788 10906
rect 19788 10854 19802 10906
rect 19826 10854 19840 10906
rect 19840 10854 19852 10906
rect 19852 10854 19882 10906
rect 19906 10854 19916 10906
rect 19916 10854 19962 10906
rect 19666 10852 19722 10854
rect 19746 10852 19802 10854
rect 19826 10852 19882 10854
rect 19906 10852 19962 10854
rect 23518 19066 23574 19068
rect 23598 19066 23654 19068
rect 23678 19066 23734 19068
rect 23758 19066 23814 19068
rect 23518 19014 23564 19066
rect 23564 19014 23574 19066
rect 23598 19014 23628 19066
rect 23628 19014 23640 19066
rect 23640 19014 23654 19066
rect 23678 19014 23692 19066
rect 23692 19014 23704 19066
rect 23704 19014 23734 19066
rect 23758 19014 23768 19066
rect 23768 19014 23814 19066
rect 23518 19012 23574 19014
rect 23598 19012 23654 19014
rect 23678 19012 23734 19014
rect 23758 19012 23814 19014
rect 31223 19066 31279 19068
rect 31303 19066 31359 19068
rect 31383 19066 31439 19068
rect 31463 19066 31519 19068
rect 31223 19014 31269 19066
rect 31269 19014 31279 19066
rect 31303 19014 31333 19066
rect 31333 19014 31345 19066
rect 31345 19014 31359 19066
rect 31383 19014 31397 19066
rect 31397 19014 31409 19066
rect 31409 19014 31439 19066
rect 31463 19014 31473 19066
rect 31473 19014 31519 19066
rect 31223 19012 31279 19014
rect 31303 19012 31359 19014
rect 31383 19012 31439 19014
rect 31463 19012 31519 19014
rect 27371 18522 27427 18524
rect 27451 18522 27507 18524
rect 27531 18522 27587 18524
rect 27611 18522 27667 18524
rect 27371 18470 27417 18522
rect 27417 18470 27427 18522
rect 27451 18470 27481 18522
rect 27481 18470 27493 18522
rect 27493 18470 27507 18522
rect 27531 18470 27545 18522
rect 27545 18470 27557 18522
rect 27557 18470 27587 18522
rect 27611 18470 27621 18522
rect 27621 18470 27667 18522
rect 27371 18468 27427 18470
rect 27451 18468 27507 18470
rect 27531 18468 27587 18470
rect 27611 18468 27667 18470
rect 23518 17978 23574 17980
rect 23598 17978 23654 17980
rect 23678 17978 23734 17980
rect 23758 17978 23814 17980
rect 23518 17926 23564 17978
rect 23564 17926 23574 17978
rect 23598 17926 23628 17978
rect 23628 17926 23640 17978
rect 23640 17926 23654 17978
rect 23678 17926 23692 17978
rect 23692 17926 23704 17978
rect 23704 17926 23734 17978
rect 23758 17926 23768 17978
rect 23768 17926 23814 17978
rect 23518 17924 23574 17926
rect 23598 17924 23654 17926
rect 23678 17924 23734 17926
rect 23758 17924 23814 17926
rect 31223 17978 31279 17980
rect 31303 17978 31359 17980
rect 31383 17978 31439 17980
rect 31463 17978 31519 17980
rect 31223 17926 31269 17978
rect 31269 17926 31279 17978
rect 31303 17926 31333 17978
rect 31333 17926 31345 17978
rect 31345 17926 31359 17978
rect 31383 17926 31397 17978
rect 31397 17926 31409 17978
rect 31409 17926 31439 17978
rect 31463 17926 31473 17978
rect 31473 17926 31519 17978
rect 31223 17924 31279 17926
rect 31303 17924 31359 17926
rect 31383 17924 31439 17926
rect 31463 17924 31519 17926
rect 27371 17434 27427 17436
rect 27451 17434 27507 17436
rect 27531 17434 27587 17436
rect 27611 17434 27667 17436
rect 27371 17382 27417 17434
rect 27417 17382 27427 17434
rect 27451 17382 27481 17434
rect 27481 17382 27493 17434
rect 27493 17382 27507 17434
rect 27531 17382 27545 17434
rect 27545 17382 27557 17434
rect 27557 17382 27587 17434
rect 27611 17382 27621 17434
rect 27621 17382 27667 17434
rect 27371 17380 27427 17382
rect 27451 17380 27507 17382
rect 27531 17380 27587 17382
rect 27611 17380 27667 17382
rect 23518 16890 23574 16892
rect 23598 16890 23654 16892
rect 23678 16890 23734 16892
rect 23758 16890 23814 16892
rect 23518 16838 23564 16890
rect 23564 16838 23574 16890
rect 23598 16838 23628 16890
rect 23628 16838 23640 16890
rect 23640 16838 23654 16890
rect 23678 16838 23692 16890
rect 23692 16838 23704 16890
rect 23704 16838 23734 16890
rect 23758 16838 23768 16890
rect 23768 16838 23814 16890
rect 23518 16836 23574 16838
rect 23598 16836 23654 16838
rect 23678 16836 23734 16838
rect 23758 16836 23814 16838
rect 31223 16890 31279 16892
rect 31303 16890 31359 16892
rect 31383 16890 31439 16892
rect 31463 16890 31519 16892
rect 31223 16838 31269 16890
rect 31269 16838 31279 16890
rect 31303 16838 31333 16890
rect 31333 16838 31345 16890
rect 31345 16838 31359 16890
rect 31383 16838 31397 16890
rect 31397 16838 31409 16890
rect 31409 16838 31439 16890
rect 31463 16838 31473 16890
rect 31473 16838 31519 16890
rect 31223 16836 31279 16838
rect 31303 16836 31359 16838
rect 31383 16836 31439 16838
rect 31463 16836 31519 16838
rect 27371 16346 27427 16348
rect 27451 16346 27507 16348
rect 27531 16346 27587 16348
rect 27611 16346 27667 16348
rect 27371 16294 27417 16346
rect 27417 16294 27427 16346
rect 27451 16294 27481 16346
rect 27481 16294 27493 16346
rect 27493 16294 27507 16346
rect 27531 16294 27545 16346
rect 27545 16294 27557 16346
rect 27557 16294 27587 16346
rect 27611 16294 27621 16346
rect 27621 16294 27667 16346
rect 27371 16292 27427 16294
rect 27451 16292 27507 16294
rect 27531 16292 27587 16294
rect 27611 16292 27667 16294
rect 23518 15802 23574 15804
rect 23598 15802 23654 15804
rect 23678 15802 23734 15804
rect 23758 15802 23814 15804
rect 23518 15750 23564 15802
rect 23564 15750 23574 15802
rect 23598 15750 23628 15802
rect 23628 15750 23640 15802
rect 23640 15750 23654 15802
rect 23678 15750 23692 15802
rect 23692 15750 23704 15802
rect 23704 15750 23734 15802
rect 23758 15750 23768 15802
rect 23768 15750 23814 15802
rect 23518 15748 23574 15750
rect 23598 15748 23654 15750
rect 23678 15748 23734 15750
rect 23758 15748 23814 15750
rect 31223 15802 31279 15804
rect 31303 15802 31359 15804
rect 31383 15802 31439 15804
rect 31463 15802 31519 15804
rect 31223 15750 31269 15802
rect 31269 15750 31279 15802
rect 31303 15750 31333 15802
rect 31333 15750 31345 15802
rect 31345 15750 31359 15802
rect 31383 15750 31397 15802
rect 31397 15750 31409 15802
rect 31409 15750 31439 15802
rect 31463 15750 31473 15802
rect 31473 15750 31519 15802
rect 31223 15748 31279 15750
rect 31303 15748 31359 15750
rect 31383 15748 31439 15750
rect 31463 15748 31519 15750
rect 27371 15258 27427 15260
rect 27451 15258 27507 15260
rect 27531 15258 27587 15260
rect 27611 15258 27667 15260
rect 27371 15206 27417 15258
rect 27417 15206 27427 15258
rect 27451 15206 27481 15258
rect 27481 15206 27493 15258
rect 27493 15206 27507 15258
rect 27531 15206 27545 15258
rect 27545 15206 27557 15258
rect 27557 15206 27587 15258
rect 27611 15206 27621 15258
rect 27621 15206 27667 15258
rect 27371 15204 27427 15206
rect 27451 15204 27507 15206
rect 27531 15204 27587 15206
rect 27611 15204 27667 15206
rect 27986 15000 28042 15056
rect 23518 14714 23574 14716
rect 23598 14714 23654 14716
rect 23678 14714 23734 14716
rect 23758 14714 23814 14716
rect 23518 14662 23564 14714
rect 23564 14662 23574 14714
rect 23598 14662 23628 14714
rect 23628 14662 23640 14714
rect 23640 14662 23654 14714
rect 23678 14662 23692 14714
rect 23692 14662 23704 14714
rect 23704 14662 23734 14714
rect 23758 14662 23768 14714
rect 23768 14662 23814 14714
rect 23518 14660 23574 14662
rect 23598 14660 23654 14662
rect 23678 14660 23734 14662
rect 23758 14660 23814 14662
rect 27371 14170 27427 14172
rect 27451 14170 27507 14172
rect 27531 14170 27587 14172
rect 27611 14170 27667 14172
rect 27371 14118 27417 14170
rect 27417 14118 27427 14170
rect 27451 14118 27481 14170
rect 27481 14118 27493 14170
rect 27493 14118 27507 14170
rect 27531 14118 27545 14170
rect 27545 14118 27557 14170
rect 27557 14118 27587 14170
rect 27611 14118 27621 14170
rect 27621 14118 27667 14170
rect 27371 14116 27427 14118
rect 27451 14116 27507 14118
rect 27531 14116 27587 14118
rect 27611 14116 27667 14118
rect 23518 13626 23574 13628
rect 23598 13626 23654 13628
rect 23678 13626 23734 13628
rect 23758 13626 23814 13628
rect 23518 13574 23564 13626
rect 23564 13574 23574 13626
rect 23598 13574 23628 13626
rect 23628 13574 23640 13626
rect 23640 13574 23654 13626
rect 23678 13574 23692 13626
rect 23692 13574 23704 13626
rect 23704 13574 23734 13626
rect 23758 13574 23768 13626
rect 23768 13574 23814 13626
rect 23518 13572 23574 13574
rect 23598 13572 23654 13574
rect 23678 13572 23734 13574
rect 23758 13572 23814 13574
rect 27371 13082 27427 13084
rect 27451 13082 27507 13084
rect 27531 13082 27587 13084
rect 27611 13082 27667 13084
rect 27371 13030 27417 13082
rect 27417 13030 27427 13082
rect 27451 13030 27481 13082
rect 27481 13030 27493 13082
rect 27493 13030 27507 13082
rect 27531 13030 27545 13082
rect 27545 13030 27557 13082
rect 27557 13030 27587 13082
rect 27611 13030 27621 13082
rect 27621 13030 27667 13082
rect 27371 13028 27427 13030
rect 27451 13028 27507 13030
rect 27531 13028 27587 13030
rect 27611 13028 27667 13030
rect 31223 14714 31279 14716
rect 31303 14714 31359 14716
rect 31383 14714 31439 14716
rect 31463 14714 31519 14716
rect 31223 14662 31269 14714
rect 31269 14662 31279 14714
rect 31303 14662 31333 14714
rect 31333 14662 31345 14714
rect 31345 14662 31359 14714
rect 31383 14662 31397 14714
rect 31397 14662 31409 14714
rect 31409 14662 31439 14714
rect 31463 14662 31473 14714
rect 31473 14662 31519 14714
rect 31223 14660 31279 14662
rect 31303 14660 31359 14662
rect 31383 14660 31439 14662
rect 31463 14660 31519 14662
rect 28446 14320 28502 14376
rect 28262 12980 28318 13016
rect 28262 12960 28264 12980
rect 28264 12960 28316 12980
rect 28316 12960 28318 12980
rect 23518 12538 23574 12540
rect 23598 12538 23654 12540
rect 23678 12538 23734 12540
rect 23758 12538 23814 12540
rect 23518 12486 23564 12538
rect 23564 12486 23574 12538
rect 23598 12486 23628 12538
rect 23628 12486 23640 12538
rect 23640 12486 23654 12538
rect 23678 12486 23692 12538
rect 23692 12486 23704 12538
rect 23704 12486 23734 12538
rect 23758 12486 23768 12538
rect 23768 12486 23814 12538
rect 23518 12484 23574 12486
rect 23598 12484 23654 12486
rect 23678 12484 23734 12486
rect 23758 12484 23814 12486
rect 31666 13640 31722 13696
rect 31223 13626 31279 13628
rect 31303 13626 31359 13628
rect 31383 13626 31439 13628
rect 31463 13626 31519 13628
rect 31223 13574 31269 13626
rect 31269 13574 31279 13626
rect 31303 13574 31333 13626
rect 31333 13574 31345 13626
rect 31345 13574 31359 13626
rect 31383 13574 31397 13626
rect 31397 13574 31409 13626
rect 31409 13574 31439 13626
rect 31463 13574 31473 13626
rect 31473 13574 31519 13626
rect 31223 13572 31279 13574
rect 31303 13572 31359 13574
rect 31383 13572 31439 13574
rect 31463 13572 31519 13574
rect 15813 9274 15869 9276
rect 15893 9274 15949 9276
rect 15973 9274 16029 9276
rect 16053 9274 16109 9276
rect 15813 9222 15859 9274
rect 15859 9222 15869 9274
rect 15893 9222 15923 9274
rect 15923 9222 15935 9274
rect 15935 9222 15949 9274
rect 15973 9222 15987 9274
rect 15987 9222 15999 9274
rect 15999 9222 16029 9274
rect 16053 9222 16063 9274
rect 16063 9222 16109 9274
rect 15813 9220 15869 9222
rect 15893 9220 15949 9222
rect 15973 9220 16029 9222
rect 16053 9220 16109 9222
rect 15813 8186 15869 8188
rect 15893 8186 15949 8188
rect 15973 8186 16029 8188
rect 16053 8186 16109 8188
rect 15813 8134 15859 8186
rect 15859 8134 15869 8186
rect 15893 8134 15923 8186
rect 15923 8134 15935 8186
rect 15935 8134 15949 8186
rect 15973 8134 15987 8186
rect 15987 8134 15999 8186
rect 15999 8134 16029 8186
rect 16053 8134 16063 8186
rect 16063 8134 16109 8186
rect 15813 8132 15869 8134
rect 15893 8132 15949 8134
rect 15973 8132 16029 8134
rect 16053 8132 16109 8134
rect 19666 9818 19722 9820
rect 19746 9818 19802 9820
rect 19826 9818 19882 9820
rect 19906 9818 19962 9820
rect 19666 9766 19712 9818
rect 19712 9766 19722 9818
rect 19746 9766 19776 9818
rect 19776 9766 19788 9818
rect 19788 9766 19802 9818
rect 19826 9766 19840 9818
rect 19840 9766 19852 9818
rect 19852 9766 19882 9818
rect 19906 9766 19916 9818
rect 19916 9766 19962 9818
rect 19666 9764 19722 9766
rect 19746 9764 19802 9766
rect 19826 9764 19882 9766
rect 19906 9764 19962 9766
rect 15813 7098 15869 7100
rect 15893 7098 15949 7100
rect 15973 7098 16029 7100
rect 16053 7098 16109 7100
rect 15813 7046 15859 7098
rect 15859 7046 15869 7098
rect 15893 7046 15923 7098
rect 15923 7046 15935 7098
rect 15935 7046 15949 7098
rect 15973 7046 15987 7098
rect 15987 7046 15999 7098
rect 15999 7046 16029 7098
rect 16053 7046 16063 7098
rect 16063 7046 16109 7098
rect 15813 7044 15869 7046
rect 15893 7044 15949 7046
rect 15973 7044 16029 7046
rect 16053 7044 16109 7046
rect 15813 6010 15869 6012
rect 15893 6010 15949 6012
rect 15973 6010 16029 6012
rect 16053 6010 16109 6012
rect 15813 5958 15859 6010
rect 15859 5958 15869 6010
rect 15893 5958 15923 6010
rect 15923 5958 15935 6010
rect 15935 5958 15949 6010
rect 15973 5958 15987 6010
rect 15987 5958 15999 6010
rect 15999 5958 16029 6010
rect 16053 5958 16063 6010
rect 16063 5958 16109 6010
rect 15813 5956 15869 5958
rect 15893 5956 15949 5958
rect 15973 5956 16029 5958
rect 16053 5956 16109 5958
rect 15813 4922 15869 4924
rect 15893 4922 15949 4924
rect 15973 4922 16029 4924
rect 16053 4922 16109 4924
rect 15813 4870 15859 4922
rect 15859 4870 15869 4922
rect 15893 4870 15923 4922
rect 15923 4870 15935 4922
rect 15935 4870 15949 4922
rect 15973 4870 15987 4922
rect 15987 4870 15999 4922
rect 15999 4870 16029 4922
rect 16053 4870 16063 4922
rect 16063 4870 16109 4922
rect 15813 4868 15869 4870
rect 15893 4868 15949 4870
rect 15973 4868 16029 4870
rect 16053 4868 16109 4870
rect 15813 3834 15869 3836
rect 15893 3834 15949 3836
rect 15973 3834 16029 3836
rect 16053 3834 16109 3836
rect 15813 3782 15859 3834
rect 15859 3782 15869 3834
rect 15893 3782 15923 3834
rect 15923 3782 15935 3834
rect 15935 3782 15949 3834
rect 15973 3782 15987 3834
rect 15987 3782 15999 3834
rect 15999 3782 16029 3834
rect 16053 3782 16063 3834
rect 16063 3782 16109 3834
rect 15813 3780 15869 3782
rect 15893 3780 15949 3782
rect 15973 3780 16029 3782
rect 16053 3780 16109 3782
rect 15813 2746 15869 2748
rect 15893 2746 15949 2748
rect 15973 2746 16029 2748
rect 16053 2746 16109 2748
rect 15813 2694 15859 2746
rect 15859 2694 15869 2746
rect 15893 2694 15923 2746
rect 15923 2694 15935 2746
rect 15935 2694 15949 2746
rect 15973 2694 15987 2746
rect 15987 2694 15999 2746
rect 15999 2694 16029 2746
rect 16053 2694 16063 2746
rect 16063 2694 16109 2746
rect 15813 2692 15869 2694
rect 15893 2692 15949 2694
rect 15973 2692 16029 2694
rect 16053 2692 16109 2694
rect 15813 1658 15869 1660
rect 15893 1658 15949 1660
rect 15973 1658 16029 1660
rect 16053 1658 16109 1660
rect 15813 1606 15859 1658
rect 15859 1606 15869 1658
rect 15893 1606 15923 1658
rect 15923 1606 15935 1658
rect 15935 1606 15949 1658
rect 15973 1606 15987 1658
rect 15987 1606 15999 1658
rect 15999 1606 16029 1658
rect 16053 1606 16063 1658
rect 16063 1606 16109 1658
rect 15813 1604 15869 1606
rect 15893 1604 15949 1606
rect 15973 1604 16029 1606
rect 16053 1604 16109 1606
rect 15813 570 15869 572
rect 15893 570 15949 572
rect 15973 570 16029 572
rect 16053 570 16109 572
rect 15813 518 15859 570
rect 15859 518 15869 570
rect 15893 518 15923 570
rect 15923 518 15935 570
rect 15935 518 15949 570
rect 15973 518 15987 570
rect 15987 518 15999 570
rect 15999 518 16029 570
rect 16053 518 16063 570
rect 16063 518 16109 570
rect 15813 516 15869 518
rect 15893 516 15949 518
rect 15973 516 16029 518
rect 16053 516 16109 518
rect 19666 8730 19722 8732
rect 19746 8730 19802 8732
rect 19826 8730 19882 8732
rect 19906 8730 19962 8732
rect 19666 8678 19712 8730
rect 19712 8678 19722 8730
rect 19746 8678 19776 8730
rect 19776 8678 19788 8730
rect 19788 8678 19802 8730
rect 19826 8678 19840 8730
rect 19840 8678 19852 8730
rect 19852 8678 19882 8730
rect 19906 8678 19916 8730
rect 19916 8678 19962 8730
rect 19666 8676 19722 8678
rect 19746 8676 19802 8678
rect 19826 8676 19882 8678
rect 19906 8676 19962 8678
rect 19666 7642 19722 7644
rect 19746 7642 19802 7644
rect 19826 7642 19882 7644
rect 19906 7642 19962 7644
rect 19666 7590 19712 7642
rect 19712 7590 19722 7642
rect 19746 7590 19776 7642
rect 19776 7590 19788 7642
rect 19788 7590 19802 7642
rect 19826 7590 19840 7642
rect 19840 7590 19852 7642
rect 19852 7590 19882 7642
rect 19906 7590 19916 7642
rect 19916 7590 19962 7642
rect 19666 7588 19722 7590
rect 19746 7588 19802 7590
rect 19826 7588 19882 7590
rect 19906 7588 19962 7590
rect 19666 6554 19722 6556
rect 19746 6554 19802 6556
rect 19826 6554 19882 6556
rect 19906 6554 19962 6556
rect 19666 6502 19712 6554
rect 19712 6502 19722 6554
rect 19746 6502 19776 6554
rect 19776 6502 19788 6554
rect 19788 6502 19802 6554
rect 19826 6502 19840 6554
rect 19840 6502 19852 6554
rect 19852 6502 19882 6554
rect 19906 6502 19916 6554
rect 19916 6502 19962 6554
rect 19666 6500 19722 6502
rect 19746 6500 19802 6502
rect 19826 6500 19882 6502
rect 19906 6500 19962 6502
rect 19666 5466 19722 5468
rect 19746 5466 19802 5468
rect 19826 5466 19882 5468
rect 19906 5466 19962 5468
rect 19666 5414 19712 5466
rect 19712 5414 19722 5466
rect 19746 5414 19776 5466
rect 19776 5414 19788 5466
rect 19788 5414 19802 5466
rect 19826 5414 19840 5466
rect 19840 5414 19852 5466
rect 19852 5414 19882 5466
rect 19906 5414 19916 5466
rect 19916 5414 19962 5466
rect 19666 5412 19722 5414
rect 19746 5412 19802 5414
rect 19826 5412 19882 5414
rect 19906 5412 19962 5414
rect 19666 4378 19722 4380
rect 19746 4378 19802 4380
rect 19826 4378 19882 4380
rect 19906 4378 19962 4380
rect 19666 4326 19712 4378
rect 19712 4326 19722 4378
rect 19746 4326 19776 4378
rect 19776 4326 19788 4378
rect 19788 4326 19802 4378
rect 19826 4326 19840 4378
rect 19840 4326 19852 4378
rect 19852 4326 19882 4378
rect 19906 4326 19916 4378
rect 19916 4326 19962 4378
rect 19666 4324 19722 4326
rect 19746 4324 19802 4326
rect 19826 4324 19882 4326
rect 19906 4324 19962 4326
rect 19666 3290 19722 3292
rect 19746 3290 19802 3292
rect 19826 3290 19882 3292
rect 19906 3290 19962 3292
rect 19666 3238 19712 3290
rect 19712 3238 19722 3290
rect 19746 3238 19776 3290
rect 19776 3238 19788 3290
rect 19788 3238 19802 3290
rect 19826 3238 19840 3290
rect 19840 3238 19852 3290
rect 19852 3238 19882 3290
rect 19906 3238 19916 3290
rect 19916 3238 19962 3290
rect 19666 3236 19722 3238
rect 19746 3236 19802 3238
rect 19826 3236 19882 3238
rect 19906 3236 19962 3238
rect 19666 2202 19722 2204
rect 19746 2202 19802 2204
rect 19826 2202 19882 2204
rect 19906 2202 19962 2204
rect 19666 2150 19712 2202
rect 19712 2150 19722 2202
rect 19746 2150 19776 2202
rect 19776 2150 19788 2202
rect 19788 2150 19802 2202
rect 19826 2150 19840 2202
rect 19840 2150 19852 2202
rect 19852 2150 19882 2202
rect 19906 2150 19916 2202
rect 19916 2150 19962 2202
rect 19666 2148 19722 2150
rect 19746 2148 19802 2150
rect 19826 2148 19882 2150
rect 19906 2148 19962 2150
rect 19666 1114 19722 1116
rect 19746 1114 19802 1116
rect 19826 1114 19882 1116
rect 19906 1114 19962 1116
rect 19666 1062 19712 1114
rect 19712 1062 19722 1114
rect 19746 1062 19776 1114
rect 19776 1062 19788 1114
rect 19788 1062 19802 1114
rect 19826 1062 19840 1114
rect 19840 1062 19852 1114
rect 19852 1062 19882 1114
rect 19906 1062 19916 1114
rect 19916 1062 19962 1114
rect 19666 1060 19722 1062
rect 19746 1060 19802 1062
rect 19826 1060 19882 1062
rect 19906 1060 19962 1062
rect 28262 12280 28318 12336
rect 27371 11994 27427 11996
rect 27451 11994 27507 11996
rect 27531 11994 27587 11996
rect 27611 11994 27667 11996
rect 27371 11942 27417 11994
rect 27417 11942 27427 11994
rect 27451 11942 27481 11994
rect 27481 11942 27493 11994
rect 27493 11942 27507 11994
rect 27531 11942 27545 11994
rect 27545 11942 27557 11994
rect 27557 11942 27587 11994
rect 27611 11942 27621 11994
rect 27621 11942 27667 11994
rect 27371 11940 27427 11942
rect 27451 11940 27507 11942
rect 27531 11940 27587 11942
rect 27611 11940 27667 11942
rect 31223 12538 31279 12540
rect 31303 12538 31359 12540
rect 31383 12538 31439 12540
rect 31463 12538 31519 12540
rect 31223 12486 31269 12538
rect 31269 12486 31279 12538
rect 31303 12486 31333 12538
rect 31333 12486 31345 12538
rect 31345 12486 31359 12538
rect 31383 12486 31397 12538
rect 31397 12486 31409 12538
rect 31409 12486 31439 12538
rect 31463 12486 31473 12538
rect 31473 12486 31519 12538
rect 31223 12484 31279 12486
rect 31303 12484 31359 12486
rect 31383 12484 31439 12486
rect 31463 12484 31519 12486
rect 28262 11600 28318 11656
rect 23518 11450 23574 11452
rect 23598 11450 23654 11452
rect 23678 11450 23734 11452
rect 23758 11450 23814 11452
rect 23518 11398 23564 11450
rect 23564 11398 23574 11450
rect 23598 11398 23628 11450
rect 23628 11398 23640 11450
rect 23640 11398 23654 11450
rect 23678 11398 23692 11450
rect 23692 11398 23704 11450
rect 23704 11398 23734 11450
rect 23758 11398 23768 11450
rect 23768 11398 23814 11450
rect 23518 11396 23574 11398
rect 23598 11396 23654 11398
rect 23678 11396 23734 11398
rect 23758 11396 23814 11398
rect 31223 11450 31279 11452
rect 31303 11450 31359 11452
rect 31383 11450 31439 11452
rect 31463 11450 31519 11452
rect 31223 11398 31269 11450
rect 31269 11398 31279 11450
rect 31303 11398 31333 11450
rect 31333 11398 31345 11450
rect 31345 11398 31359 11450
rect 31383 11398 31397 11450
rect 31397 11398 31409 11450
rect 31409 11398 31439 11450
rect 31463 11398 31473 11450
rect 31473 11398 31519 11450
rect 31223 11396 31279 11398
rect 31303 11396 31359 11398
rect 31383 11396 31439 11398
rect 31463 11396 31519 11398
rect 28262 10920 28318 10976
rect 27371 10906 27427 10908
rect 27451 10906 27507 10908
rect 27531 10906 27587 10908
rect 27611 10906 27667 10908
rect 27371 10854 27417 10906
rect 27417 10854 27427 10906
rect 27451 10854 27481 10906
rect 27481 10854 27493 10906
rect 27493 10854 27507 10906
rect 27531 10854 27545 10906
rect 27545 10854 27557 10906
rect 27557 10854 27587 10906
rect 27611 10854 27621 10906
rect 27621 10854 27667 10906
rect 27371 10852 27427 10854
rect 27451 10852 27507 10854
rect 27531 10852 27587 10854
rect 27611 10852 27667 10854
rect 23518 10362 23574 10364
rect 23598 10362 23654 10364
rect 23678 10362 23734 10364
rect 23758 10362 23814 10364
rect 23518 10310 23564 10362
rect 23564 10310 23574 10362
rect 23598 10310 23628 10362
rect 23628 10310 23640 10362
rect 23640 10310 23654 10362
rect 23678 10310 23692 10362
rect 23692 10310 23704 10362
rect 23704 10310 23734 10362
rect 23758 10310 23768 10362
rect 23768 10310 23814 10362
rect 23518 10308 23574 10310
rect 23598 10308 23654 10310
rect 23678 10308 23734 10310
rect 23758 10308 23814 10310
rect 31223 10362 31279 10364
rect 31303 10362 31359 10364
rect 31383 10362 31439 10364
rect 31463 10362 31519 10364
rect 31223 10310 31269 10362
rect 31269 10310 31279 10362
rect 31303 10310 31333 10362
rect 31333 10310 31345 10362
rect 31345 10310 31359 10362
rect 31383 10310 31397 10362
rect 31397 10310 31409 10362
rect 31409 10310 31439 10362
rect 31463 10310 31473 10362
rect 31473 10310 31519 10362
rect 31223 10308 31279 10310
rect 31303 10308 31359 10310
rect 31383 10308 31439 10310
rect 31463 10308 31519 10310
rect 31666 10240 31722 10296
rect 27371 9818 27427 9820
rect 27451 9818 27507 9820
rect 27531 9818 27587 9820
rect 27611 9818 27667 9820
rect 27371 9766 27417 9818
rect 27417 9766 27427 9818
rect 27451 9766 27481 9818
rect 27481 9766 27493 9818
rect 27493 9766 27507 9818
rect 27531 9766 27545 9818
rect 27545 9766 27557 9818
rect 27557 9766 27587 9818
rect 27611 9766 27621 9818
rect 27621 9766 27667 9818
rect 27371 9764 27427 9766
rect 27451 9764 27507 9766
rect 27531 9764 27587 9766
rect 27611 9764 27667 9766
rect 28262 9560 28318 9616
rect 23518 9274 23574 9276
rect 23598 9274 23654 9276
rect 23678 9274 23734 9276
rect 23758 9274 23814 9276
rect 23518 9222 23564 9274
rect 23564 9222 23574 9274
rect 23598 9222 23628 9274
rect 23628 9222 23640 9274
rect 23640 9222 23654 9274
rect 23678 9222 23692 9274
rect 23692 9222 23704 9274
rect 23704 9222 23734 9274
rect 23758 9222 23768 9274
rect 23768 9222 23814 9274
rect 23518 9220 23574 9222
rect 23598 9220 23654 9222
rect 23678 9220 23734 9222
rect 23758 9220 23814 9222
rect 31223 9274 31279 9276
rect 31303 9274 31359 9276
rect 31383 9274 31439 9276
rect 31463 9274 31519 9276
rect 31223 9222 31269 9274
rect 31269 9222 31279 9274
rect 31303 9222 31333 9274
rect 31333 9222 31345 9274
rect 31345 9222 31359 9274
rect 31383 9222 31397 9274
rect 31397 9222 31409 9274
rect 31409 9222 31439 9274
rect 31463 9222 31473 9274
rect 31473 9222 31519 9274
rect 31223 9220 31279 9222
rect 31303 9220 31359 9222
rect 31383 9220 31439 9222
rect 31463 9220 31519 9222
rect 28262 8880 28318 8936
rect 27371 8730 27427 8732
rect 27451 8730 27507 8732
rect 27531 8730 27587 8732
rect 27611 8730 27667 8732
rect 27371 8678 27417 8730
rect 27417 8678 27427 8730
rect 27451 8678 27481 8730
rect 27481 8678 27493 8730
rect 27493 8678 27507 8730
rect 27531 8678 27545 8730
rect 27545 8678 27557 8730
rect 27557 8678 27587 8730
rect 27611 8678 27621 8730
rect 27621 8678 27667 8730
rect 27371 8676 27427 8678
rect 27451 8676 27507 8678
rect 27531 8676 27587 8678
rect 27611 8676 27667 8678
rect 23386 8472 23442 8528
rect 23518 8186 23574 8188
rect 23598 8186 23654 8188
rect 23678 8186 23734 8188
rect 23758 8186 23814 8188
rect 23518 8134 23564 8186
rect 23564 8134 23574 8186
rect 23598 8134 23628 8186
rect 23628 8134 23640 8186
rect 23640 8134 23654 8186
rect 23678 8134 23692 8186
rect 23692 8134 23704 8186
rect 23704 8134 23734 8186
rect 23758 8134 23768 8186
rect 23768 8134 23814 8186
rect 23518 8132 23574 8134
rect 23598 8132 23654 8134
rect 23678 8132 23734 8134
rect 23758 8132 23814 8134
rect 27371 7642 27427 7644
rect 27451 7642 27507 7644
rect 27531 7642 27587 7644
rect 27611 7642 27667 7644
rect 27371 7590 27417 7642
rect 27417 7590 27427 7642
rect 27451 7590 27481 7642
rect 27481 7590 27493 7642
rect 27493 7590 27507 7642
rect 27531 7590 27545 7642
rect 27545 7590 27557 7642
rect 27557 7590 27587 7642
rect 27611 7590 27621 7642
rect 27621 7590 27667 7642
rect 27371 7588 27427 7590
rect 27451 7588 27507 7590
rect 27531 7588 27587 7590
rect 27611 7588 27667 7590
rect 28262 7520 28318 7576
rect 23518 7098 23574 7100
rect 23598 7098 23654 7100
rect 23678 7098 23734 7100
rect 23758 7098 23814 7100
rect 23518 7046 23564 7098
rect 23564 7046 23574 7098
rect 23598 7046 23628 7098
rect 23628 7046 23640 7098
rect 23640 7046 23654 7098
rect 23678 7046 23692 7098
rect 23692 7046 23704 7098
rect 23704 7046 23734 7098
rect 23758 7046 23768 7098
rect 23768 7046 23814 7098
rect 23518 7044 23574 7046
rect 23598 7044 23654 7046
rect 23678 7044 23734 7046
rect 23758 7044 23814 7046
rect 28262 6840 28318 6896
rect 27371 6554 27427 6556
rect 27451 6554 27507 6556
rect 27531 6554 27587 6556
rect 27611 6554 27667 6556
rect 27371 6502 27417 6554
rect 27417 6502 27427 6554
rect 27451 6502 27481 6554
rect 27481 6502 27493 6554
rect 27493 6502 27507 6554
rect 27531 6502 27545 6554
rect 27545 6502 27557 6554
rect 27557 6502 27587 6554
rect 27611 6502 27621 6554
rect 27621 6502 27667 6554
rect 27371 6500 27427 6502
rect 27451 6500 27507 6502
rect 27531 6500 27587 6502
rect 27611 6500 27667 6502
rect 28262 6160 28318 6216
rect 23518 6010 23574 6012
rect 23598 6010 23654 6012
rect 23678 6010 23734 6012
rect 23758 6010 23814 6012
rect 23518 5958 23564 6010
rect 23564 5958 23574 6010
rect 23598 5958 23628 6010
rect 23628 5958 23640 6010
rect 23640 5958 23654 6010
rect 23678 5958 23692 6010
rect 23692 5958 23704 6010
rect 23704 5958 23734 6010
rect 23758 5958 23768 6010
rect 23768 5958 23814 6010
rect 23518 5956 23574 5958
rect 23598 5956 23654 5958
rect 23678 5956 23734 5958
rect 23758 5956 23814 5958
rect 31666 8472 31722 8528
rect 31666 8200 31722 8256
rect 31223 8186 31279 8188
rect 31303 8186 31359 8188
rect 31383 8186 31439 8188
rect 31463 8186 31519 8188
rect 31223 8134 31269 8186
rect 31269 8134 31279 8186
rect 31303 8134 31333 8186
rect 31333 8134 31345 8186
rect 31345 8134 31359 8186
rect 31383 8134 31397 8186
rect 31397 8134 31409 8186
rect 31409 8134 31439 8186
rect 31463 8134 31473 8186
rect 31473 8134 31519 8186
rect 31223 8132 31279 8134
rect 31303 8132 31359 8134
rect 31383 8132 31439 8134
rect 31463 8132 31519 8134
rect 31223 7098 31279 7100
rect 31303 7098 31359 7100
rect 31383 7098 31439 7100
rect 31463 7098 31519 7100
rect 31223 7046 31269 7098
rect 31269 7046 31279 7098
rect 31303 7046 31333 7098
rect 31333 7046 31345 7098
rect 31345 7046 31359 7098
rect 31383 7046 31397 7098
rect 31397 7046 31409 7098
rect 31409 7046 31439 7098
rect 31463 7046 31473 7098
rect 31473 7046 31519 7098
rect 31223 7044 31279 7046
rect 31303 7044 31359 7046
rect 31383 7044 31439 7046
rect 31463 7044 31519 7046
rect 31223 6010 31279 6012
rect 31303 6010 31359 6012
rect 31383 6010 31439 6012
rect 31463 6010 31519 6012
rect 31223 5958 31269 6010
rect 31269 5958 31279 6010
rect 31303 5958 31333 6010
rect 31333 5958 31345 6010
rect 31345 5958 31359 6010
rect 31383 5958 31397 6010
rect 31397 5958 31409 6010
rect 31409 5958 31439 6010
rect 31463 5958 31473 6010
rect 31473 5958 31519 6010
rect 31223 5956 31279 5958
rect 31303 5956 31359 5958
rect 31383 5956 31439 5958
rect 31463 5956 31519 5958
rect 28446 5480 28502 5536
rect 27371 5466 27427 5468
rect 27451 5466 27507 5468
rect 27531 5466 27587 5468
rect 27611 5466 27667 5468
rect 27371 5414 27417 5466
rect 27417 5414 27427 5466
rect 27451 5414 27481 5466
rect 27481 5414 27493 5466
rect 27493 5414 27507 5466
rect 27531 5414 27545 5466
rect 27545 5414 27557 5466
rect 27557 5414 27587 5466
rect 27611 5414 27621 5466
rect 27621 5414 27667 5466
rect 27371 5412 27427 5414
rect 27451 5412 27507 5414
rect 27531 5412 27587 5414
rect 27611 5412 27667 5414
rect 23518 4922 23574 4924
rect 23598 4922 23654 4924
rect 23678 4922 23734 4924
rect 23758 4922 23814 4924
rect 23518 4870 23564 4922
rect 23564 4870 23574 4922
rect 23598 4870 23628 4922
rect 23628 4870 23640 4922
rect 23640 4870 23654 4922
rect 23678 4870 23692 4922
rect 23692 4870 23704 4922
rect 23704 4870 23734 4922
rect 23758 4870 23768 4922
rect 23768 4870 23814 4922
rect 23518 4868 23574 4870
rect 23598 4868 23654 4870
rect 23678 4868 23734 4870
rect 23758 4868 23814 4870
rect 31223 4922 31279 4924
rect 31303 4922 31359 4924
rect 31383 4922 31439 4924
rect 31463 4922 31519 4924
rect 31223 4870 31269 4922
rect 31269 4870 31279 4922
rect 31303 4870 31333 4922
rect 31333 4870 31345 4922
rect 31345 4870 31359 4922
rect 31383 4870 31397 4922
rect 31397 4870 31409 4922
rect 31409 4870 31439 4922
rect 31463 4870 31473 4922
rect 31473 4870 31519 4922
rect 31223 4868 31279 4870
rect 31303 4868 31359 4870
rect 31383 4868 31439 4870
rect 31463 4868 31519 4870
rect 27371 4378 27427 4380
rect 27451 4378 27507 4380
rect 27531 4378 27587 4380
rect 27611 4378 27667 4380
rect 27371 4326 27417 4378
rect 27417 4326 27427 4378
rect 27451 4326 27481 4378
rect 27481 4326 27493 4378
rect 27493 4326 27507 4378
rect 27531 4326 27545 4378
rect 27545 4326 27557 4378
rect 27557 4326 27587 4378
rect 27611 4326 27621 4378
rect 27621 4326 27667 4378
rect 27371 4324 27427 4326
rect 27451 4324 27507 4326
rect 27531 4324 27587 4326
rect 27611 4324 27667 4326
rect 23518 3834 23574 3836
rect 23598 3834 23654 3836
rect 23678 3834 23734 3836
rect 23758 3834 23814 3836
rect 23518 3782 23564 3834
rect 23564 3782 23574 3834
rect 23598 3782 23628 3834
rect 23628 3782 23640 3834
rect 23640 3782 23654 3834
rect 23678 3782 23692 3834
rect 23692 3782 23704 3834
rect 23704 3782 23734 3834
rect 23758 3782 23768 3834
rect 23768 3782 23814 3834
rect 23518 3780 23574 3782
rect 23598 3780 23654 3782
rect 23678 3780 23734 3782
rect 23758 3780 23814 3782
rect 31223 3834 31279 3836
rect 31303 3834 31359 3836
rect 31383 3834 31439 3836
rect 31463 3834 31519 3836
rect 31223 3782 31269 3834
rect 31269 3782 31279 3834
rect 31303 3782 31333 3834
rect 31333 3782 31345 3834
rect 31345 3782 31359 3834
rect 31383 3782 31397 3834
rect 31397 3782 31409 3834
rect 31409 3782 31439 3834
rect 31463 3782 31473 3834
rect 31473 3782 31519 3834
rect 31223 3780 31279 3782
rect 31303 3780 31359 3782
rect 31383 3780 31439 3782
rect 31463 3780 31519 3782
rect 27371 3290 27427 3292
rect 27451 3290 27507 3292
rect 27531 3290 27587 3292
rect 27611 3290 27667 3292
rect 27371 3238 27417 3290
rect 27417 3238 27427 3290
rect 27451 3238 27481 3290
rect 27481 3238 27493 3290
rect 27493 3238 27507 3290
rect 27531 3238 27545 3290
rect 27545 3238 27557 3290
rect 27557 3238 27587 3290
rect 27611 3238 27621 3290
rect 27621 3238 27667 3290
rect 27371 3236 27427 3238
rect 27451 3236 27507 3238
rect 27531 3236 27587 3238
rect 27611 3236 27667 3238
rect 23518 2746 23574 2748
rect 23598 2746 23654 2748
rect 23678 2746 23734 2748
rect 23758 2746 23814 2748
rect 23518 2694 23564 2746
rect 23564 2694 23574 2746
rect 23598 2694 23628 2746
rect 23628 2694 23640 2746
rect 23640 2694 23654 2746
rect 23678 2694 23692 2746
rect 23692 2694 23704 2746
rect 23704 2694 23734 2746
rect 23758 2694 23768 2746
rect 23768 2694 23814 2746
rect 23518 2692 23574 2694
rect 23598 2692 23654 2694
rect 23678 2692 23734 2694
rect 23758 2692 23814 2694
rect 31223 2746 31279 2748
rect 31303 2746 31359 2748
rect 31383 2746 31439 2748
rect 31463 2746 31519 2748
rect 31223 2694 31269 2746
rect 31269 2694 31279 2746
rect 31303 2694 31333 2746
rect 31333 2694 31345 2746
rect 31345 2694 31359 2746
rect 31383 2694 31397 2746
rect 31397 2694 31409 2746
rect 31409 2694 31439 2746
rect 31463 2694 31473 2746
rect 31473 2694 31519 2746
rect 31223 2692 31279 2694
rect 31303 2692 31359 2694
rect 31383 2692 31439 2694
rect 31463 2692 31519 2694
rect 27371 2202 27427 2204
rect 27451 2202 27507 2204
rect 27531 2202 27587 2204
rect 27611 2202 27667 2204
rect 27371 2150 27417 2202
rect 27417 2150 27427 2202
rect 27451 2150 27481 2202
rect 27481 2150 27493 2202
rect 27493 2150 27507 2202
rect 27531 2150 27545 2202
rect 27545 2150 27557 2202
rect 27557 2150 27587 2202
rect 27611 2150 27621 2202
rect 27621 2150 27667 2202
rect 27371 2148 27427 2150
rect 27451 2148 27507 2150
rect 27531 2148 27587 2150
rect 27611 2148 27667 2150
rect 23518 1658 23574 1660
rect 23598 1658 23654 1660
rect 23678 1658 23734 1660
rect 23758 1658 23814 1660
rect 23518 1606 23564 1658
rect 23564 1606 23574 1658
rect 23598 1606 23628 1658
rect 23628 1606 23640 1658
rect 23640 1606 23654 1658
rect 23678 1606 23692 1658
rect 23692 1606 23704 1658
rect 23704 1606 23734 1658
rect 23758 1606 23768 1658
rect 23768 1606 23814 1658
rect 23518 1604 23574 1606
rect 23598 1604 23654 1606
rect 23678 1604 23734 1606
rect 23758 1604 23814 1606
rect 31223 1658 31279 1660
rect 31303 1658 31359 1660
rect 31383 1658 31439 1660
rect 31463 1658 31519 1660
rect 31223 1606 31269 1658
rect 31269 1606 31279 1658
rect 31303 1606 31333 1658
rect 31333 1606 31345 1658
rect 31345 1606 31359 1658
rect 31383 1606 31397 1658
rect 31397 1606 31409 1658
rect 31409 1606 31439 1658
rect 31463 1606 31473 1658
rect 31473 1606 31519 1658
rect 31223 1604 31279 1606
rect 31303 1604 31359 1606
rect 31383 1604 31439 1606
rect 31463 1604 31519 1606
rect 27371 1114 27427 1116
rect 27451 1114 27507 1116
rect 27531 1114 27587 1116
rect 27611 1114 27667 1116
rect 27371 1062 27417 1114
rect 27417 1062 27427 1114
rect 27451 1062 27481 1114
rect 27481 1062 27493 1114
rect 27493 1062 27507 1114
rect 27531 1062 27545 1114
rect 27545 1062 27557 1114
rect 27557 1062 27587 1114
rect 27611 1062 27621 1114
rect 27621 1062 27667 1114
rect 27371 1060 27427 1062
rect 27451 1060 27507 1062
rect 27531 1060 27587 1062
rect 27611 1060 27667 1062
rect 23518 570 23574 572
rect 23598 570 23654 572
rect 23678 570 23734 572
rect 23758 570 23814 572
rect 23518 518 23564 570
rect 23564 518 23574 570
rect 23598 518 23628 570
rect 23628 518 23640 570
rect 23640 518 23654 570
rect 23678 518 23692 570
rect 23692 518 23704 570
rect 23704 518 23734 570
rect 23758 518 23768 570
rect 23768 518 23814 570
rect 23518 516 23574 518
rect 23598 516 23654 518
rect 23678 516 23734 518
rect 23758 516 23814 518
rect 31223 570 31279 572
rect 31303 570 31359 572
rect 31383 570 31439 572
rect 31463 570 31519 572
rect 31223 518 31269 570
rect 31269 518 31279 570
rect 31303 518 31333 570
rect 31333 518 31345 570
rect 31345 518 31359 570
rect 31383 518 31397 570
rect 31397 518 31409 570
rect 31409 518 31439 570
rect 31463 518 31473 570
rect 31473 518 31519 570
rect 31223 516 31279 518
rect 31303 516 31359 518
rect 31383 516 31439 518
rect 31463 516 31519 518
<< metal3 >>
rect 8098 19072 8414 19073
rect 8098 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8414 19072
rect 8098 19007 8414 19008
rect 15803 19072 16119 19073
rect 15803 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16119 19072
rect 15803 19007 16119 19008
rect 23508 19072 23824 19073
rect 23508 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23824 19072
rect 23508 19007 23824 19008
rect 31213 19072 31529 19073
rect 31213 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31529 19072
rect 31213 19007 31529 19008
rect 4246 18528 4562 18529
rect 4246 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4562 18528
rect 4246 18463 4562 18464
rect 11951 18528 12267 18529
rect 11951 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12267 18528
rect 11951 18463 12267 18464
rect 19656 18528 19972 18529
rect 19656 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19972 18528
rect 19656 18463 19972 18464
rect 27361 18528 27677 18529
rect 27361 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27677 18528
rect 27361 18463 27677 18464
rect 8098 17984 8414 17985
rect 8098 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8414 17984
rect 8098 17919 8414 17920
rect 15803 17984 16119 17985
rect 15803 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16119 17984
rect 15803 17919 16119 17920
rect 23508 17984 23824 17985
rect 23508 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23824 17984
rect 23508 17919 23824 17920
rect 31213 17984 31529 17985
rect 31213 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31529 17984
rect 31213 17919 31529 17920
rect 4246 17440 4562 17441
rect 4246 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4562 17440
rect 4246 17375 4562 17376
rect 11951 17440 12267 17441
rect 11951 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12267 17440
rect 11951 17375 12267 17376
rect 19656 17440 19972 17441
rect 19656 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19972 17440
rect 19656 17375 19972 17376
rect 27361 17440 27677 17441
rect 27361 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27677 17440
rect 27361 17375 27677 17376
rect 8098 16896 8414 16897
rect 8098 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8414 16896
rect 8098 16831 8414 16832
rect 15803 16896 16119 16897
rect 15803 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16119 16896
rect 15803 16831 16119 16832
rect 23508 16896 23824 16897
rect 23508 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23824 16896
rect 23508 16831 23824 16832
rect 31213 16896 31529 16897
rect 31213 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31529 16896
rect 31213 16831 31529 16832
rect 4246 16352 4562 16353
rect 4246 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4562 16352
rect 4246 16287 4562 16288
rect 11951 16352 12267 16353
rect 11951 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12267 16352
rect 11951 16287 12267 16288
rect 19656 16352 19972 16353
rect 19656 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19972 16352
rect 19656 16287 19972 16288
rect 27361 16352 27677 16353
rect 27361 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27677 16352
rect 27361 16287 27677 16288
rect 8098 15808 8414 15809
rect 8098 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8414 15808
rect 8098 15743 8414 15744
rect 15803 15808 16119 15809
rect 15803 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16119 15808
rect 15803 15743 16119 15744
rect 23508 15808 23824 15809
rect 23508 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23824 15808
rect 23508 15743 23824 15744
rect 31213 15808 31529 15809
rect 31213 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31529 15808
rect 31213 15743 31529 15744
rect 4246 15264 4562 15265
rect 4246 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4562 15264
rect 4246 15199 4562 15200
rect 11951 15264 12267 15265
rect 11951 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12267 15264
rect 11951 15199 12267 15200
rect 19656 15264 19972 15265
rect 19656 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19972 15264
rect 19656 15199 19972 15200
rect 27361 15264 27677 15265
rect 27361 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27677 15264
rect 27361 15199 27677 15200
rect 27981 15058 28047 15061
rect 31600 15058 32000 15088
rect 27981 15056 32000 15058
rect 27981 15000 27986 15056
rect 28042 15000 32000 15056
rect 27981 14998 32000 15000
rect 27981 14995 28047 14998
rect 31600 14968 32000 14998
rect 8098 14720 8414 14721
rect 8098 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8414 14720
rect 8098 14655 8414 14656
rect 15803 14720 16119 14721
rect 15803 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16119 14720
rect 15803 14655 16119 14656
rect 23508 14720 23824 14721
rect 23508 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23824 14720
rect 23508 14655 23824 14656
rect 31213 14720 31529 14721
rect 31213 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31529 14720
rect 31213 14655 31529 14656
rect 28441 14378 28507 14381
rect 31600 14378 32000 14408
rect 28441 14376 32000 14378
rect 28441 14320 28446 14376
rect 28502 14320 32000 14376
rect 28441 14318 32000 14320
rect 28441 14315 28507 14318
rect 31600 14288 32000 14318
rect 4246 14176 4562 14177
rect 4246 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4562 14176
rect 4246 14111 4562 14112
rect 11951 14176 12267 14177
rect 11951 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12267 14176
rect 11951 14111 12267 14112
rect 19656 14176 19972 14177
rect 19656 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19972 14176
rect 19656 14111 19972 14112
rect 27361 14176 27677 14177
rect 27361 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27677 14176
rect 27361 14111 27677 14112
rect 31600 13696 32000 13728
rect 31600 13640 31666 13696
rect 31722 13640 32000 13696
rect 8098 13632 8414 13633
rect 8098 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8414 13632
rect 8098 13567 8414 13568
rect 15803 13632 16119 13633
rect 15803 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16119 13632
rect 15803 13567 16119 13568
rect 23508 13632 23824 13633
rect 23508 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23824 13632
rect 23508 13567 23824 13568
rect 31213 13632 31529 13633
rect 31213 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31529 13632
rect 31600 13608 32000 13640
rect 31213 13567 31529 13568
rect 4246 13088 4562 13089
rect 4246 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4562 13088
rect 4246 13023 4562 13024
rect 11951 13088 12267 13089
rect 11951 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12267 13088
rect 11951 13023 12267 13024
rect 19656 13088 19972 13089
rect 19656 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19972 13088
rect 19656 13023 19972 13024
rect 27361 13088 27677 13089
rect 27361 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27677 13088
rect 27361 13023 27677 13024
rect 28257 13018 28323 13021
rect 31600 13018 32000 13048
rect 28257 13016 32000 13018
rect 28257 12960 28262 13016
rect 28318 12960 32000 13016
rect 28257 12958 32000 12960
rect 28257 12955 28323 12958
rect 31600 12928 32000 12958
rect 8098 12544 8414 12545
rect 8098 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8414 12544
rect 8098 12479 8414 12480
rect 15803 12544 16119 12545
rect 15803 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16119 12544
rect 15803 12479 16119 12480
rect 23508 12544 23824 12545
rect 23508 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23824 12544
rect 23508 12479 23824 12480
rect 31213 12544 31529 12545
rect 31213 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31529 12544
rect 31213 12479 31529 12480
rect 0 12338 400 12368
rect 6913 12338 6979 12341
rect 0 12336 6979 12338
rect 0 12280 6918 12336
rect 6974 12280 6979 12336
rect 0 12278 6979 12280
rect 0 12248 400 12278
rect 6913 12275 6979 12278
rect 28257 12338 28323 12341
rect 31600 12338 32000 12368
rect 28257 12336 32000 12338
rect 28257 12280 28262 12336
rect 28318 12280 32000 12336
rect 28257 12278 32000 12280
rect 28257 12275 28323 12278
rect 31600 12248 32000 12278
rect 4246 12000 4562 12001
rect 4246 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4562 12000
rect 4246 11935 4562 11936
rect 11951 12000 12267 12001
rect 11951 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12267 12000
rect 11951 11935 12267 11936
rect 19656 12000 19972 12001
rect 19656 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19972 12000
rect 19656 11935 19972 11936
rect 27361 12000 27677 12001
rect 27361 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27677 12000
rect 27361 11935 27677 11936
rect 0 11658 400 11688
rect 6913 11658 6979 11661
rect 0 11656 6979 11658
rect 0 11600 6918 11656
rect 6974 11600 6979 11656
rect 0 11598 6979 11600
rect 0 11568 400 11598
rect 6913 11595 6979 11598
rect 28257 11658 28323 11661
rect 31600 11658 32000 11688
rect 28257 11656 32000 11658
rect 28257 11600 28262 11656
rect 28318 11600 32000 11656
rect 28257 11598 32000 11600
rect 28257 11595 28323 11598
rect 31600 11568 32000 11598
rect 8098 11456 8414 11457
rect 8098 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8414 11456
rect 8098 11391 8414 11392
rect 15803 11456 16119 11457
rect 15803 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16119 11456
rect 15803 11391 16119 11392
rect 23508 11456 23824 11457
rect 23508 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23824 11456
rect 23508 11391 23824 11392
rect 31213 11456 31529 11457
rect 31213 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31529 11456
rect 31213 11391 31529 11392
rect 0 10978 400 11008
rect 28257 10978 28323 10981
rect 31600 10978 32000 11008
rect 0 10918 2790 10978
rect 0 10888 400 10918
rect 2730 10706 2790 10918
rect 28257 10976 32000 10978
rect 28257 10920 28262 10976
rect 28318 10920 32000 10976
rect 28257 10918 32000 10920
rect 28257 10915 28323 10918
rect 4246 10912 4562 10913
rect 4246 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4562 10912
rect 4246 10847 4562 10848
rect 11951 10912 12267 10913
rect 11951 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12267 10912
rect 11951 10847 12267 10848
rect 19656 10912 19972 10913
rect 19656 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19972 10912
rect 19656 10847 19972 10848
rect 27361 10912 27677 10913
rect 27361 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27677 10912
rect 31600 10888 32000 10918
rect 27361 10847 27677 10848
rect 11145 10842 11211 10845
rect 4662 10840 11211 10842
rect 4662 10784 11150 10840
rect 11206 10784 11211 10840
rect 4662 10782 11211 10784
rect 4662 10706 4722 10782
rect 11145 10779 11211 10782
rect 2730 10646 4722 10706
rect 8098 10368 8414 10369
rect 0 10298 400 10328
rect 8098 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8414 10368
rect 8098 10303 8414 10304
rect 15803 10368 16119 10369
rect 15803 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16119 10368
rect 15803 10303 16119 10304
rect 23508 10368 23824 10369
rect 23508 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23824 10368
rect 23508 10303 23824 10304
rect 31213 10368 31529 10369
rect 31213 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31529 10368
rect 31213 10303 31529 10304
rect 7097 10298 7163 10301
rect 0 10296 7163 10298
rect 0 10240 7102 10296
rect 7158 10240 7163 10296
rect 0 10238 7163 10240
rect 0 10208 400 10238
rect 7097 10235 7163 10238
rect 31600 10296 32000 10328
rect 31600 10240 31666 10296
rect 31722 10240 32000 10296
rect 31600 10208 32000 10240
rect 4246 9824 4562 9825
rect 4246 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4562 9824
rect 4246 9759 4562 9760
rect 11951 9824 12267 9825
rect 11951 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12267 9824
rect 11951 9759 12267 9760
rect 19656 9824 19972 9825
rect 19656 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19972 9824
rect 19656 9759 19972 9760
rect 27361 9824 27677 9825
rect 27361 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27677 9824
rect 27361 9759 27677 9760
rect 0 9618 400 9648
rect 9765 9618 9831 9621
rect 0 9616 9831 9618
rect 0 9560 9770 9616
rect 9826 9560 9831 9616
rect 0 9558 9831 9560
rect 0 9528 400 9558
rect 9765 9555 9831 9558
rect 28257 9618 28323 9621
rect 31600 9618 32000 9648
rect 28257 9616 32000 9618
rect 28257 9560 28262 9616
rect 28318 9560 32000 9616
rect 28257 9558 32000 9560
rect 28257 9555 28323 9558
rect 31600 9528 32000 9558
rect 8098 9280 8414 9281
rect 8098 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8414 9280
rect 8098 9215 8414 9216
rect 15803 9280 16119 9281
rect 15803 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16119 9280
rect 15803 9215 16119 9216
rect 23508 9280 23824 9281
rect 23508 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23824 9280
rect 23508 9215 23824 9216
rect 31213 9280 31529 9281
rect 31213 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31529 9280
rect 31213 9215 31529 9216
rect 0 8938 400 8968
rect 6729 8938 6795 8941
rect 0 8936 6795 8938
rect 0 8880 6734 8936
rect 6790 8880 6795 8936
rect 0 8878 6795 8880
rect 0 8848 400 8878
rect 6729 8875 6795 8878
rect 28257 8938 28323 8941
rect 31600 8938 32000 8968
rect 28257 8936 32000 8938
rect 28257 8880 28262 8936
rect 28318 8880 32000 8936
rect 28257 8878 32000 8880
rect 28257 8875 28323 8878
rect 31600 8848 32000 8878
rect 4246 8736 4562 8737
rect 4246 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4562 8736
rect 4246 8671 4562 8672
rect 11951 8736 12267 8737
rect 11951 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12267 8736
rect 11951 8671 12267 8672
rect 19656 8736 19972 8737
rect 19656 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19972 8736
rect 19656 8671 19972 8672
rect 27361 8736 27677 8737
rect 27361 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27677 8736
rect 27361 8671 27677 8672
rect 23381 8530 23447 8533
rect 31661 8530 31727 8533
rect 23381 8528 31727 8530
rect 23381 8472 23386 8528
rect 23442 8472 31666 8528
rect 31722 8472 31727 8528
rect 23381 8470 31727 8472
rect 23381 8467 23447 8470
rect 31661 8467 31727 8470
rect 0 8258 400 8288
rect 0 8198 2790 8258
rect 0 8168 400 8198
rect 2730 7986 2790 8198
rect 31600 8256 32000 8288
rect 31600 8200 31666 8256
rect 31722 8200 32000 8256
rect 8098 8192 8414 8193
rect 8098 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8414 8192
rect 8098 8127 8414 8128
rect 15803 8192 16119 8193
rect 15803 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16119 8192
rect 15803 8127 16119 8128
rect 23508 8192 23824 8193
rect 23508 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23824 8192
rect 23508 8127 23824 8128
rect 31213 8192 31529 8193
rect 31213 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31529 8192
rect 31600 8168 32000 8200
rect 31213 8127 31529 8128
rect 9397 7986 9463 7989
rect 2730 7984 9463 7986
rect 2730 7928 9402 7984
rect 9458 7928 9463 7984
rect 2730 7926 9463 7928
rect 9397 7923 9463 7926
rect 9305 7850 9371 7853
rect 2730 7848 9371 7850
rect 2730 7792 9310 7848
rect 9366 7792 9371 7848
rect 2730 7790 9371 7792
rect 0 7578 400 7608
rect 2730 7578 2790 7790
rect 9305 7787 9371 7790
rect 4246 7648 4562 7649
rect 4246 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4562 7648
rect 4246 7583 4562 7584
rect 11951 7648 12267 7649
rect 11951 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12267 7648
rect 11951 7583 12267 7584
rect 19656 7648 19972 7649
rect 19656 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19972 7648
rect 19656 7583 19972 7584
rect 27361 7648 27677 7649
rect 27361 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27677 7648
rect 27361 7583 27677 7584
rect 0 7518 2790 7578
rect 28257 7578 28323 7581
rect 31600 7578 32000 7608
rect 28257 7576 32000 7578
rect 28257 7520 28262 7576
rect 28318 7520 32000 7576
rect 28257 7518 32000 7520
rect 0 7488 400 7518
rect 28257 7515 28323 7518
rect 31600 7488 32000 7518
rect 8098 7104 8414 7105
rect 8098 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8414 7104
rect 8098 7039 8414 7040
rect 15803 7104 16119 7105
rect 15803 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16119 7104
rect 15803 7039 16119 7040
rect 23508 7104 23824 7105
rect 23508 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23824 7104
rect 23508 7039 23824 7040
rect 31213 7104 31529 7105
rect 31213 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31529 7104
rect 31213 7039 31529 7040
rect 0 6898 400 6928
rect 6637 6898 6703 6901
rect 0 6896 6703 6898
rect 0 6840 6642 6896
rect 6698 6840 6703 6896
rect 0 6838 6703 6840
rect 0 6808 400 6838
rect 6637 6835 6703 6838
rect 28257 6898 28323 6901
rect 31600 6898 32000 6928
rect 28257 6896 32000 6898
rect 28257 6840 28262 6896
rect 28318 6840 32000 6896
rect 28257 6838 32000 6840
rect 28257 6835 28323 6838
rect 31600 6808 32000 6838
rect 4246 6560 4562 6561
rect 4246 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4562 6560
rect 4246 6495 4562 6496
rect 11951 6560 12267 6561
rect 11951 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12267 6560
rect 11951 6495 12267 6496
rect 19656 6560 19972 6561
rect 19656 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19972 6560
rect 19656 6495 19972 6496
rect 27361 6560 27677 6561
rect 27361 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27677 6560
rect 27361 6495 27677 6496
rect 0 6218 400 6248
rect 7833 6218 7899 6221
rect 0 6216 7899 6218
rect 0 6160 7838 6216
rect 7894 6160 7899 6216
rect 0 6158 7899 6160
rect 0 6128 400 6158
rect 7833 6155 7899 6158
rect 28257 6218 28323 6221
rect 31600 6218 32000 6248
rect 28257 6216 32000 6218
rect 28257 6160 28262 6216
rect 28318 6160 32000 6216
rect 28257 6158 32000 6160
rect 28257 6155 28323 6158
rect 31600 6128 32000 6158
rect 8098 6016 8414 6017
rect 8098 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8414 6016
rect 8098 5951 8414 5952
rect 15803 6016 16119 6017
rect 15803 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16119 6016
rect 15803 5951 16119 5952
rect 23508 6016 23824 6017
rect 23508 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23824 6016
rect 23508 5951 23824 5952
rect 31213 6016 31529 6017
rect 31213 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31529 6016
rect 31213 5951 31529 5952
rect 28441 5538 28507 5541
rect 31600 5538 32000 5568
rect 28441 5536 32000 5538
rect 28441 5480 28446 5536
rect 28502 5480 32000 5536
rect 28441 5478 32000 5480
rect 28441 5475 28507 5478
rect 4246 5472 4562 5473
rect 4246 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4562 5472
rect 4246 5407 4562 5408
rect 11951 5472 12267 5473
rect 11951 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12267 5472
rect 11951 5407 12267 5408
rect 19656 5472 19972 5473
rect 19656 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19972 5472
rect 19656 5407 19972 5408
rect 27361 5472 27677 5473
rect 27361 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27677 5472
rect 31600 5448 32000 5478
rect 27361 5407 27677 5408
rect 8098 4928 8414 4929
rect 8098 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8414 4928
rect 8098 4863 8414 4864
rect 15803 4928 16119 4929
rect 15803 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16119 4928
rect 15803 4863 16119 4864
rect 23508 4928 23824 4929
rect 23508 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23824 4928
rect 23508 4863 23824 4864
rect 31213 4928 31529 4929
rect 31213 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31529 4928
rect 31213 4863 31529 4864
rect 4246 4384 4562 4385
rect 4246 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4562 4384
rect 4246 4319 4562 4320
rect 11951 4384 12267 4385
rect 11951 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12267 4384
rect 11951 4319 12267 4320
rect 19656 4384 19972 4385
rect 19656 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19972 4384
rect 19656 4319 19972 4320
rect 27361 4384 27677 4385
rect 27361 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27677 4384
rect 27361 4319 27677 4320
rect 8098 3840 8414 3841
rect 8098 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8414 3840
rect 8098 3775 8414 3776
rect 15803 3840 16119 3841
rect 15803 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16119 3840
rect 15803 3775 16119 3776
rect 23508 3840 23824 3841
rect 23508 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23824 3840
rect 23508 3775 23824 3776
rect 31213 3840 31529 3841
rect 31213 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31529 3840
rect 31213 3775 31529 3776
rect 4246 3296 4562 3297
rect 4246 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4562 3296
rect 4246 3231 4562 3232
rect 11951 3296 12267 3297
rect 11951 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12267 3296
rect 11951 3231 12267 3232
rect 19656 3296 19972 3297
rect 19656 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19972 3296
rect 19656 3231 19972 3232
rect 27361 3296 27677 3297
rect 27361 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27677 3296
rect 27361 3231 27677 3232
rect 8098 2752 8414 2753
rect 8098 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8414 2752
rect 8098 2687 8414 2688
rect 15803 2752 16119 2753
rect 15803 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16119 2752
rect 15803 2687 16119 2688
rect 23508 2752 23824 2753
rect 23508 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23824 2752
rect 23508 2687 23824 2688
rect 31213 2752 31529 2753
rect 31213 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31529 2752
rect 31213 2687 31529 2688
rect 4246 2208 4562 2209
rect 4246 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4562 2208
rect 4246 2143 4562 2144
rect 11951 2208 12267 2209
rect 11951 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12267 2208
rect 11951 2143 12267 2144
rect 19656 2208 19972 2209
rect 19656 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19972 2208
rect 19656 2143 19972 2144
rect 27361 2208 27677 2209
rect 27361 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27677 2208
rect 27361 2143 27677 2144
rect 8098 1664 8414 1665
rect 8098 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8414 1664
rect 8098 1599 8414 1600
rect 15803 1664 16119 1665
rect 15803 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16119 1664
rect 15803 1599 16119 1600
rect 23508 1664 23824 1665
rect 23508 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23824 1664
rect 23508 1599 23824 1600
rect 31213 1664 31529 1665
rect 31213 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31529 1664
rect 31213 1599 31529 1600
rect 4246 1120 4562 1121
rect 4246 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4562 1120
rect 4246 1055 4562 1056
rect 11951 1120 12267 1121
rect 11951 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12267 1120
rect 11951 1055 12267 1056
rect 19656 1120 19972 1121
rect 19656 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19972 1120
rect 19656 1055 19972 1056
rect 27361 1120 27677 1121
rect 27361 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27677 1120
rect 27361 1055 27677 1056
rect 8098 576 8414 577
rect 8098 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8414 576
rect 8098 511 8414 512
rect 15803 576 16119 577
rect 15803 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16119 576
rect 15803 511 16119 512
rect 23508 576 23824 577
rect 23508 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23824 576
rect 23508 511 23824 512
rect 31213 576 31529 577
rect 31213 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31529 576
rect 31213 511 31529 512
<< via3 >>
rect 8104 19068 8168 19072
rect 8104 19012 8108 19068
rect 8108 19012 8164 19068
rect 8164 19012 8168 19068
rect 8104 19008 8168 19012
rect 8184 19068 8248 19072
rect 8184 19012 8188 19068
rect 8188 19012 8244 19068
rect 8244 19012 8248 19068
rect 8184 19008 8248 19012
rect 8264 19068 8328 19072
rect 8264 19012 8268 19068
rect 8268 19012 8324 19068
rect 8324 19012 8328 19068
rect 8264 19008 8328 19012
rect 8344 19068 8408 19072
rect 8344 19012 8348 19068
rect 8348 19012 8404 19068
rect 8404 19012 8408 19068
rect 8344 19008 8408 19012
rect 15809 19068 15873 19072
rect 15809 19012 15813 19068
rect 15813 19012 15869 19068
rect 15869 19012 15873 19068
rect 15809 19008 15873 19012
rect 15889 19068 15953 19072
rect 15889 19012 15893 19068
rect 15893 19012 15949 19068
rect 15949 19012 15953 19068
rect 15889 19008 15953 19012
rect 15969 19068 16033 19072
rect 15969 19012 15973 19068
rect 15973 19012 16029 19068
rect 16029 19012 16033 19068
rect 15969 19008 16033 19012
rect 16049 19068 16113 19072
rect 16049 19012 16053 19068
rect 16053 19012 16109 19068
rect 16109 19012 16113 19068
rect 16049 19008 16113 19012
rect 23514 19068 23578 19072
rect 23514 19012 23518 19068
rect 23518 19012 23574 19068
rect 23574 19012 23578 19068
rect 23514 19008 23578 19012
rect 23594 19068 23658 19072
rect 23594 19012 23598 19068
rect 23598 19012 23654 19068
rect 23654 19012 23658 19068
rect 23594 19008 23658 19012
rect 23674 19068 23738 19072
rect 23674 19012 23678 19068
rect 23678 19012 23734 19068
rect 23734 19012 23738 19068
rect 23674 19008 23738 19012
rect 23754 19068 23818 19072
rect 23754 19012 23758 19068
rect 23758 19012 23814 19068
rect 23814 19012 23818 19068
rect 23754 19008 23818 19012
rect 31219 19068 31283 19072
rect 31219 19012 31223 19068
rect 31223 19012 31279 19068
rect 31279 19012 31283 19068
rect 31219 19008 31283 19012
rect 31299 19068 31363 19072
rect 31299 19012 31303 19068
rect 31303 19012 31359 19068
rect 31359 19012 31363 19068
rect 31299 19008 31363 19012
rect 31379 19068 31443 19072
rect 31379 19012 31383 19068
rect 31383 19012 31439 19068
rect 31439 19012 31443 19068
rect 31379 19008 31443 19012
rect 31459 19068 31523 19072
rect 31459 19012 31463 19068
rect 31463 19012 31519 19068
rect 31519 19012 31523 19068
rect 31459 19008 31523 19012
rect 4252 18524 4316 18528
rect 4252 18468 4256 18524
rect 4256 18468 4312 18524
rect 4312 18468 4316 18524
rect 4252 18464 4316 18468
rect 4332 18524 4396 18528
rect 4332 18468 4336 18524
rect 4336 18468 4392 18524
rect 4392 18468 4396 18524
rect 4332 18464 4396 18468
rect 4412 18524 4476 18528
rect 4412 18468 4416 18524
rect 4416 18468 4472 18524
rect 4472 18468 4476 18524
rect 4412 18464 4476 18468
rect 4492 18524 4556 18528
rect 4492 18468 4496 18524
rect 4496 18468 4552 18524
rect 4552 18468 4556 18524
rect 4492 18464 4556 18468
rect 11957 18524 12021 18528
rect 11957 18468 11961 18524
rect 11961 18468 12017 18524
rect 12017 18468 12021 18524
rect 11957 18464 12021 18468
rect 12037 18524 12101 18528
rect 12037 18468 12041 18524
rect 12041 18468 12097 18524
rect 12097 18468 12101 18524
rect 12037 18464 12101 18468
rect 12117 18524 12181 18528
rect 12117 18468 12121 18524
rect 12121 18468 12177 18524
rect 12177 18468 12181 18524
rect 12117 18464 12181 18468
rect 12197 18524 12261 18528
rect 12197 18468 12201 18524
rect 12201 18468 12257 18524
rect 12257 18468 12261 18524
rect 12197 18464 12261 18468
rect 19662 18524 19726 18528
rect 19662 18468 19666 18524
rect 19666 18468 19722 18524
rect 19722 18468 19726 18524
rect 19662 18464 19726 18468
rect 19742 18524 19806 18528
rect 19742 18468 19746 18524
rect 19746 18468 19802 18524
rect 19802 18468 19806 18524
rect 19742 18464 19806 18468
rect 19822 18524 19886 18528
rect 19822 18468 19826 18524
rect 19826 18468 19882 18524
rect 19882 18468 19886 18524
rect 19822 18464 19886 18468
rect 19902 18524 19966 18528
rect 19902 18468 19906 18524
rect 19906 18468 19962 18524
rect 19962 18468 19966 18524
rect 19902 18464 19966 18468
rect 27367 18524 27431 18528
rect 27367 18468 27371 18524
rect 27371 18468 27427 18524
rect 27427 18468 27431 18524
rect 27367 18464 27431 18468
rect 27447 18524 27511 18528
rect 27447 18468 27451 18524
rect 27451 18468 27507 18524
rect 27507 18468 27511 18524
rect 27447 18464 27511 18468
rect 27527 18524 27591 18528
rect 27527 18468 27531 18524
rect 27531 18468 27587 18524
rect 27587 18468 27591 18524
rect 27527 18464 27591 18468
rect 27607 18524 27671 18528
rect 27607 18468 27611 18524
rect 27611 18468 27667 18524
rect 27667 18468 27671 18524
rect 27607 18464 27671 18468
rect 8104 17980 8168 17984
rect 8104 17924 8108 17980
rect 8108 17924 8164 17980
rect 8164 17924 8168 17980
rect 8104 17920 8168 17924
rect 8184 17980 8248 17984
rect 8184 17924 8188 17980
rect 8188 17924 8244 17980
rect 8244 17924 8248 17980
rect 8184 17920 8248 17924
rect 8264 17980 8328 17984
rect 8264 17924 8268 17980
rect 8268 17924 8324 17980
rect 8324 17924 8328 17980
rect 8264 17920 8328 17924
rect 8344 17980 8408 17984
rect 8344 17924 8348 17980
rect 8348 17924 8404 17980
rect 8404 17924 8408 17980
rect 8344 17920 8408 17924
rect 15809 17980 15873 17984
rect 15809 17924 15813 17980
rect 15813 17924 15869 17980
rect 15869 17924 15873 17980
rect 15809 17920 15873 17924
rect 15889 17980 15953 17984
rect 15889 17924 15893 17980
rect 15893 17924 15949 17980
rect 15949 17924 15953 17980
rect 15889 17920 15953 17924
rect 15969 17980 16033 17984
rect 15969 17924 15973 17980
rect 15973 17924 16029 17980
rect 16029 17924 16033 17980
rect 15969 17920 16033 17924
rect 16049 17980 16113 17984
rect 16049 17924 16053 17980
rect 16053 17924 16109 17980
rect 16109 17924 16113 17980
rect 16049 17920 16113 17924
rect 23514 17980 23578 17984
rect 23514 17924 23518 17980
rect 23518 17924 23574 17980
rect 23574 17924 23578 17980
rect 23514 17920 23578 17924
rect 23594 17980 23658 17984
rect 23594 17924 23598 17980
rect 23598 17924 23654 17980
rect 23654 17924 23658 17980
rect 23594 17920 23658 17924
rect 23674 17980 23738 17984
rect 23674 17924 23678 17980
rect 23678 17924 23734 17980
rect 23734 17924 23738 17980
rect 23674 17920 23738 17924
rect 23754 17980 23818 17984
rect 23754 17924 23758 17980
rect 23758 17924 23814 17980
rect 23814 17924 23818 17980
rect 23754 17920 23818 17924
rect 31219 17980 31283 17984
rect 31219 17924 31223 17980
rect 31223 17924 31279 17980
rect 31279 17924 31283 17980
rect 31219 17920 31283 17924
rect 31299 17980 31363 17984
rect 31299 17924 31303 17980
rect 31303 17924 31359 17980
rect 31359 17924 31363 17980
rect 31299 17920 31363 17924
rect 31379 17980 31443 17984
rect 31379 17924 31383 17980
rect 31383 17924 31439 17980
rect 31439 17924 31443 17980
rect 31379 17920 31443 17924
rect 31459 17980 31523 17984
rect 31459 17924 31463 17980
rect 31463 17924 31519 17980
rect 31519 17924 31523 17980
rect 31459 17920 31523 17924
rect 4252 17436 4316 17440
rect 4252 17380 4256 17436
rect 4256 17380 4312 17436
rect 4312 17380 4316 17436
rect 4252 17376 4316 17380
rect 4332 17436 4396 17440
rect 4332 17380 4336 17436
rect 4336 17380 4392 17436
rect 4392 17380 4396 17436
rect 4332 17376 4396 17380
rect 4412 17436 4476 17440
rect 4412 17380 4416 17436
rect 4416 17380 4472 17436
rect 4472 17380 4476 17436
rect 4412 17376 4476 17380
rect 4492 17436 4556 17440
rect 4492 17380 4496 17436
rect 4496 17380 4552 17436
rect 4552 17380 4556 17436
rect 4492 17376 4556 17380
rect 11957 17436 12021 17440
rect 11957 17380 11961 17436
rect 11961 17380 12017 17436
rect 12017 17380 12021 17436
rect 11957 17376 12021 17380
rect 12037 17436 12101 17440
rect 12037 17380 12041 17436
rect 12041 17380 12097 17436
rect 12097 17380 12101 17436
rect 12037 17376 12101 17380
rect 12117 17436 12181 17440
rect 12117 17380 12121 17436
rect 12121 17380 12177 17436
rect 12177 17380 12181 17436
rect 12117 17376 12181 17380
rect 12197 17436 12261 17440
rect 12197 17380 12201 17436
rect 12201 17380 12257 17436
rect 12257 17380 12261 17436
rect 12197 17376 12261 17380
rect 19662 17436 19726 17440
rect 19662 17380 19666 17436
rect 19666 17380 19722 17436
rect 19722 17380 19726 17436
rect 19662 17376 19726 17380
rect 19742 17436 19806 17440
rect 19742 17380 19746 17436
rect 19746 17380 19802 17436
rect 19802 17380 19806 17436
rect 19742 17376 19806 17380
rect 19822 17436 19886 17440
rect 19822 17380 19826 17436
rect 19826 17380 19882 17436
rect 19882 17380 19886 17436
rect 19822 17376 19886 17380
rect 19902 17436 19966 17440
rect 19902 17380 19906 17436
rect 19906 17380 19962 17436
rect 19962 17380 19966 17436
rect 19902 17376 19966 17380
rect 27367 17436 27431 17440
rect 27367 17380 27371 17436
rect 27371 17380 27427 17436
rect 27427 17380 27431 17436
rect 27367 17376 27431 17380
rect 27447 17436 27511 17440
rect 27447 17380 27451 17436
rect 27451 17380 27507 17436
rect 27507 17380 27511 17436
rect 27447 17376 27511 17380
rect 27527 17436 27591 17440
rect 27527 17380 27531 17436
rect 27531 17380 27587 17436
rect 27587 17380 27591 17436
rect 27527 17376 27591 17380
rect 27607 17436 27671 17440
rect 27607 17380 27611 17436
rect 27611 17380 27667 17436
rect 27667 17380 27671 17436
rect 27607 17376 27671 17380
rect 8104 16892 8168 16896
rect 8104 16836 8108 16892
rect 8108 16836 8164 16892
rect 8164 16836 8168 16892
rect 8104 16832 8168 16836
rect 8184 16892 8248 16896
rect 8184 16836 8188 16892
rect 8188 16836 8244 16892
rect 8244 16836 8248 16892
rect 8184 16832 8248 16836
rect 8264 16892 8328 16896
rect 8264 16836 8268 16892
rect 8268 16836 8324 16892
rect 8324 16836 8328 16892
rect 8264 16832 8328 16836
rect 8344 16892 8408 16896
rect 8344 16836 8348 16892
rect 8348 16836 8404 16892
rect 8404 16836 8408 16892
rect 8344 16832 8408 16836
rect 15809 16892 15873 16896
rect 15809 16836 15813 16892
rect 15813 16836 15869 16892
rect 15869 16836 15873 16892
rect 15809 16832 15873 16836
rect 15889 16892 15953 16896
rect 15889 16836 15893 16892
rect 15893 16836 15949 16892
rect 15949 16836 15953 16892
rect 15889 16832 15953 16836
rect 15969 16892 16033 16896
rect 15969 16836 15973 16892
rect 15973 16836 16029 16892
rect 16029 16836 16033 16892
rect 15969 16832 16033 16836
rect 16049 16892 16113 16896
rect 16049 16836 16053 16892
rect 16053 16836 16109 16892
rect 16109 16836 16113 16892
rect 16049 16832 16113 16836
rect 23514 16892 23578 16896
rect 23514 16836 23518 16892
rect 23518 16836 23574 16892
rect 23574 16836 23578 16892
rect 23514 16832 23578 16836
rect 23594 16892 23658 16896
rect 23594 16836 23598 16892
rect 23598 16836 23654 16892
rect 23654 16836 23658 16892
rect 23594 16832 23658 16836
rect 23674 16892 23738 16896
rect 23674 16836 23678 16892
rect 23678 16836 23734 16892
rect 23734 16836 23738 16892
rect 23674 16832 23738 16836
rect 23754 16892 23818 16896
rect 23754 16836 23758 16892
rect 23758 16836 23814 16892
rect 23814 16836 23818 16892
rect 23754 16832 23818 16836
rect 31219 16892 31283 16896
rect 31219 16836 31223 16892
rect 31223 16836 31279 16892
rect 31279 16836 31283 16892
rect 31219 16832 31283 16836
rect 31299 16892 31363 16896
rect 31299 16836 31303 16892
rect 31303 16836 31359 16892
rect 31359 16836 31363 16892
rect 31299 16832 31363 16836
rect 31379 16892 31443 16896
rect 31379 16836 31383 16892
rect 31383 16836 31439 16892
rect 31439 16836 31443 16892
rect 31379 16832 31443 16836
rect 31459 16892 31523 16896
rect 31459 16836 31463 16892
rect 31463 16836 31519 16892
rect 31519 16836 31523 16892
rect 31459 16832 31523 16836
rect 4252 16348 4316 16352
rect 4252 16292 4256 16348
rect 4256 16292 4312 16348
rect 4312 16292 4316 16348
rect 4252 16288 4316 16292
rect 4332 16348 4396 16352
rect 4332 16292 4336 16348
rect 4336 16292 4392 16348
rect 4392 16292 4396 16348
rect 4332 16288 4396 16292
rect 4412 16348 4476 16352
rect 4412 16292 4416 16348
rect 4416 16292 4472 16348
rect 4472 16292 4476 16348
rect 4412 16288 4476 16292
rect 4492 16348 4556 16352
rect 4492 16292 4496 16348
rect 4496 16292 4552 16348
rect 4552 16292 4556 16348
rect 4492 16288 4556 16292
rect 11957 16348 12021 16352
rect 11957 16292 11961 16348
rect 11961 16292 12017 16348
rect 12017 16292 12021 16348
rect 11957 16288 12021 16292
rect 12037 16348 12101 16352
rect 12037 16292 12041 16348
rect 12041 16292 12097 16348
rect 12097 16292 12101 16348
rect 12037 16288 12101 16292
rect 12117 16348 12181 16352
rect 12117 16292 12121 16348
rect 12121 16292 12177 16348
rect 12177 16292 12181 16348
rect 12117 16288 12181 16292
rect 12197 16348 12261 16352
rect 12197 16292 12201 16348
rect 12201 16292 12257 16348
rect 12257 16292 12261 16348
rect 12197 16288 12261 16292
rect 19662 16348 19726 16352
rect 19662 16292 19666 16348
rect 19666 16292 19722 16348
rect 19722 16292 19726 16348
rect 19662 16288 19726 16292
rect 19742 16348 19806 16352
rect 19742 16292 19746 16348
rect 19746 16292 19802 16348
rect 19802 16292 19806 16348
rect 19742 16288 19806 16292
rect 19822 16348 19886 16352
rect 19822 16292 19826 16348
rect 19826 16292 19882 16348
rect 19882 16292 19886 16348
rect 19822 16288 19886 16292
rect 19902 16348 19966 16352
rect 19902 16292 19906 16348
rect 19906 16292 19962 16348
rect 19962 16292 19966 16348
rect 19902 16288 19966 16292
rect 27367 16348 27431 16352
rect 27367 16292 27371 16348
rect 27371 16292 27427 16348
rect 27427 16292 27431 16348
rect 27367 16288 27431 16292
rect 27447 16348 27511 16352
rect 27447 16292 27451 16348
rect 27451 16292 27507 16348
rect 27507 16292 27511 16348
rect 27447 16288 27511 16292
rect 27527 16348 27591 16352
rect 27527 16292 27531 16348
rect 27531 16292 27587 16348
rect 27587 16292 27591 16348
rect 27527 16288 27591 16292
rect 27607 16348 27671 16352
rect 27607 16292 27611 16348
rect 27611 16292 27667 16348
rect 27667 16292 27671 16348
rect 27607 16288 27671 16292
rect 8104 15804 8168 15808
rect 8104 15748 8108 15804
rect 8108 15748 8164 15804
rect 8164 15748 8168 15804
rect 8104 15744 8168 15748
rect 8184 15804 8248 15808
rect 8184 15748 8188 15804
rect 8188 15748 8244 15804
rect 8244 15748 8248 15804
rect 8184 15744 8248 15748
rect 8264 15804 8328 15808
rect 8264 15748 8268 15804
rect 8268 15748 8324 15804
rect 8324 15748 8328 15804
rect 8264 15744 8328 15748
rect 8344 15804 8408 15808
rect 8344 15748 8348 15804
rect 8348 15748 8404 15804
rect 8404 15748 8408 15804
rect 8344 15744 8408 15748
rect 15809 15804 15873 15808
rect 15809 15748 15813 15804
rect 15813 15748 15869 15804
rect 15869 15748 15873 15804
rect 15809 15744 15873 15748
rect 15889 15804 15953 15808
rect 15889 15748 15893 15804
rect 15893 15748 15949 15804
rect 15949 15748 15953 15804
rect 15889 15744 15953 15748
rect 15969 15804 16033 15808
rect 15969 15748 15973 15804
rect 15973 15748 16029 15804
rect 16029 15748 16033 15804
rect 15969 15744 16033 15748
rect 16049 15804 16113 15808
rect 16049 15748 16053 15804
rect 16053 15748 16109 15804
rect 16109 15748 16113 15804
rect 16049 15744 16113 15748
rect 23514 15804 23578 15808
rect 23514 15748 23518 15804
rect 23518 15748 23574 15804
rect 23574 15748 23578 15804
rect 23514 15744 23578 15748
rect 23594 15804 23658 15808
rect 23594 15748 23598 15804
rect 23598 15748 23654 15804
rect 23654 15748 23658 15804
rect 23594 15744 23658 15748
rect 23674 15804 23738 15808
rect 23674 15748 23678 15804
rect 23678 15748 23734 15804
rect 23734 15748 23738 15804
rect 23674 15744 23738 15748
rect 23754 15804 23818 15808
rect 23754 15748 23758 15804
rect 23758 15748 23814 15804
rect 23814 15748 23818 15804
rect 23754 15744 23818 15748
rect 31219 15804 31283 15808
rect 31219 15748 31223 15804
rect 31223 15748 31279 15804
rect 31279 15748 31283 15804
rect 31219 15744 31283 15748
rect 31299 15804 31363 15808
rect 31299 15748 31303 15804
rect 31303 15748 31359 15804
rect 31359 15748 31363 15804
rect 31299 15744 31363 15748
rect 31379 15804 31443 15808
rect 31379 15748 31383 15804
rect 31383 15748 31439 15804
rect 31439 15748 31443 15804
rect 31379 15744 31443 15748
rect 31459 15804 31523 15808
rect 31459 15748 31463 15804
rect 31463 15748 31519 15804
rect 31519 15748 31523 15804
rect 31459 15744 31523 15748
rect 4252 15260 4316 15264
rect 4252 15204 4256 15260
rect 4256 15204 4312 15260
rect 4312 15204 4316 15260
rect 4252 15200 4316 15204
rect 4332 15260 4396 15264
rect 4332 15204 4336 15260
rect 4336 15204 4392 15260
rect 4392 15204 4396 15260
rect 4332 15200 4396 15204
rect 4412 15260 4476 15264
rect 4412 15204 4416 15260
rect 4416 15204 4472 15260
rect 4472 15204 4476 15260
rect 4412 15200 4476 15204
rect 4492 15260 4556 15264
rect 4492 15204 4496 15260
rect 4496 15204 4552 15260
rect 4552 15204 4556 15260
rect 4492 15200 4556 15204
rect 11957 15260 12021 15264
rect 11957 15204 11961 15260
rect 11961 15204 12017 15260
rect 12017 15204 12021 15260
rect 11957 15200 12021 15204
rect 12037 15260 12101 15264
rect 12037 15204 12041 15260
rect 12041 15204 12097 15260
rect 12097 15204 12101 15260
rect 12037 15200 12101 15204
rect 12117 15260 12181 15264
rect 12117 15204 12121 15260
rect 12121 15204 12177 15260
rect 12177 15204 12181 15260
rect 12117 15200 12181 15204
rect 12197 15260 12261 15264
rect 12197 15204 12201 15260
rect 12201 15204 12257 15260
rect 12257 15204 12261 15260
rect 12197 15200 12261 15204
rect 19662 15260 19726 15264
rect 19662 15204 19666 15260
rect 19666 15204 19722 15260
rect 19722 15204 19726 15260
rect 19662 15200 19726 15204
rect 19742 15260 19806 15264
rect 19742 15204 19746 15260
rect 19746 15204 19802 15260
rect 19802 15204 19806 15260
rect 19742 15200 19806 15204
rect 19822 15260 19886 15264
rect 19822 15204 19826 15260
rect 19826 15204 19882 15260
rect 19882 15204 19886 15260
rect 19822 15200 19886 15204
rect 19902 15260 19966 15264
rect 19902 15204 19906 15260
rect 19906 15204 19962 15260
rect 19962 15204 19966 15260
rect 19902 15200 19966 15204
rect 27367 15260 27431 15264
rect 27367 15204 27371 15260
rect 27371 15204 27427 15260
rect 27427 15204 27431 15260
rect 27367 15200 27431 15204
rect 27447 15260 27511 15264
rect 27447 15204 27451 15260
rect 27451 15204 27507 15260
rect 27507 15204 27511 15260
rect 27447 15200 27511 15204
rect 27527 15260 27591 15264
rect 27527 15204 27531 15260
rect 27531 15204 27587 15260
rect 27587 15204 27591 15260
rect 27527 15200 27591 15204
rect 27607 15260 27671 15264
rect 27607 15204 27611 15260
rect 27611 15204 27667 15260
rect 27667 15204 27671 15260
rect 27607 15200 27671 15204
rect 8104 14716 8168 14720
rect 8104 14660 8108 14716
rect 8108 14660 8164 14716
rect 8164 14660 8168 14716
rect 8104 14656 8168 14660
rect 8184 14716 8248 14720
rect 8184 14660 8188 14716
rect 8188 14660 8244 14716
rect 8244 14660 8248 14716
rect 8184 14656 8248 14660
rect 8264 14716 8328 14720
rect 8264 14660 8268 14716
rect 8268 14660 8324 14716
rect 8324 14660 8328 14716
rect 8264 14656 8328 14660
rect 8344 14716 8408 14720
rect 8344 14660 8348 14716
rect 8348 14660 8404 14716
rect 8404 14660 8408 14716
rect 8344 14656 8408 14660
rect 15809 14716 15873 14720
rect 15809 14660 15813 14716
rect 15813 14660 15869 14716
rect 15869 14660 15873 14716
rect 15809 14656 15873 14660
rect 15889 14716 15953 14720
rect 15889 14660 15893 14716
rect 15893 14660 15949 14716
rect 15949 14660 15953 14716
rect 15889 14656 15953 14660
rect 15969 14716 16033 14720
rect 15969 14660 15973 14716
rect 15973 14660 16029 14716
rect 16029 14660 16033 14716
rect 15969 14656 16033 14660
rect 16049 14716 16113 14720
rect 16049 14660 16053 14716
rect 16053 14660 16109 14716
rect 16109 14660 16113 14716
rect 16049 14656 16113 14660
rect 23514 14716 23578 14720
rect 23514 14660 23518 14716
rect 23518 14660 23574 14716
rect 23574 14660 23578 14716
rect 23514 14656 23578 14660
rect 23594 14716 23658 14720
rect 23594 14660 23598 14716
rect 23598 14660 23654 14716
rect 23654 14660 23658 14716
rect 23594 14656 23658 14660
rect 23674 14716 23738 14720
rect 23674 14660 23678 14716
rect 23678 14660 23734 14716
rect 23734 14660 23738 14716
rect 23674 14656 23738 14660
rect 23754 14716 23818 14720
rect 23754 14660 23758 14716
rect 23758 14660 23814 14716
rect 23814 14660 23818 14716
rect 23754 14656 23818 14660
rect 31219 14716 31283 14720
rect 31219 14660 31223 14716
rect 31223 14660 31279 14716
rect 31279 14660 31283 14716
rect 31219 14656 31283 14660
rect 31299 14716 31363 14720
rect 31299 14660 31303 14716
rect 31303 14660 31359 14716
rect 31359 14660 31363 14716
rect 31299 14656 31363 14660
rect 31379 14716 31443 14720
rect 31379 14660 31383 14716
rect 31383 14660 31439 14716
rect 31439 14660 31443 14716
rect 31379 14656 31443 14660
rect 31459 14716 31523 14720
rect 31459 14660 31463 14716
rect 31463 14660 31519 14716
rect 31519 14660 31523 14716
rect 31459 14656 31523 14660
rect 4252 14172 4316 14176
rect 4252 14116 4256 14172
rect 4256 14116 4312 14172
rect 4312 14116 4316 14172
rect 4252 14112 4316 14116
rect 4332 14172 4396 14176
rect 4332 14116 4336 14172
rect 4336 14116 4392 14172
rect 4392 14116 4396 14172
rect 4332 14112 4396 14116
rect 4412 14172 4476 14176
rect 4412 14116 4416 14172
rect 4416 14116 4472 14172
rect 4472 14116 4476 14172
rect 4412 14112 4476 14116
rect 4492 14172 4556 14176
rect 4492 14116 4496 14172
rect 4496 14116 4552 14172
rect 4552 14116 4556 14172
rect 4492 14112 4556 14116
rect 11957 14172 12021 14176
rect 11957 14116 11961 14172
rect 11961 14116 12017 14172
rect 12017 14116 12021 14172
rect 11957 14112 12021 14116
rect 12037 14172 12101 14176
rect 12037 14116 12041 14172
rect 12041 14116 12097 14172
rect 12097 14116 12101 14172
rect 12037 14112 12101 14116
rect 12117 14172 12181 14176
rect 12117 14116 12121 14172
rect 12121 14116 12177 14172
rect 12177 14116 12181 14172
rect 12117 14112 12181 14116
rect 12197 14172 12261 14176
rect 12197 14116 12201 14172
rect 12201 14116 12257 14172
rect 12257 14116 12261 14172
rect 12197 14112 12261 14116
rect 19662 14172 19726 14176
rect 19662 14116 19666 14172
rect 19666 14116 19722 14172
rect 19722 14116 19726 14172
rect 19662 14112 19726 14116
rect 19742 14172 19806 14176
rect 19742 14116 19746 14172
rect 19746 14116 19802 14172
rect 19802 14116 19806 14172
rect 19742 14112 19806 14116
rect 19822 14172 19886 14176
rect 19822 14116 19826 14172
rect 19826 14116 19882 14172
rect 19882 14116 19886 14172
rect 19822 14112 19886 14116
rect 19902 14172 19966 14176
rect 19902 14116 19906 14172
rect 19906 14116 19962 14172
rect 19962 14116 19966 14172
rect 19902 14112 19966 14116
rect 27367 14172 27431 14176
rect 27367 14116 27371 14172
rect 27371 14116 27427 14172
rect 27427 14116 27431 14172
rect 27367 14112 27431 14116
rect 27447 14172 27511 14176
rect 27447 14116 27451 14172
rect 27451 14116 27507 14172
rect 27507 14116 27511 14172
rect 27447 14112 27511 14116
rect 27527 14172 27591 14176
rect 27527 14116 27531 14172
rect 27531 14116 27587 14172
rect 27587 14116 27591 14172
rect 27527 14112 27591 14116
rect 27607 14172 27671 14176
rect 27607 14116 27611 14172
rect 27611 14116 27667 14172
rect 27667 14116 27671 14172
rect 27607 14112 27671 14116
rect 8104 13628 8168 13632
rect 8104 13572 8108 13628
rect 8108 13572 8164 13628
rect 8164 13572 8168 13628
rect 8104 13568 8168 13572
rect 8184 13628 8248 13632
rect 8184 13572 8188 13628
rect 8188 13572 8244 13628
rect 8244 13572 8248 13628
rect 8184 13568 8248 13572
rect 8264 13628 8328 13632
rect 8264 13572 8268 13628
rect 8268 13572 8324 13628
rect 8324 13572 8328 13628
rect 8264 13568 8328 13572
rect 8344 13628 8408 13632
rect 8344 13572 8348 13628
rect 8348 13572 8404 13628
rect 8404 13572 8408 13628
rect 8344 13568 8408 13572
rect 15809 13628 15873 13632
rect 15809 13572 15813 13628
rect 15813 13572 15869 13628
rect 15869 13572 15873 13628
rect 15809 13568 15873 13572
rect 15889 13628 15953 13632
rect 15889 13572 15893 13628
rect 15893 13572 15949 13628
rect 15949 13572 15953 13628
rect 15889 13568 15953 13572
rect 15969 13628 16033 13632
rect 15969 13572 15973 13628
rect 15973 13572 16029 13628
rect 16029 13572 16033 13628
rect 15969 13568 16033 13572
rect 16049 13628 16113 13632
rect 16049 13572 16053 13628
rect 16053 13572 16109 13628
rect 16109 13572 16113 13628
rect 16049 13568 16113 13572
rect 23514 13628 23578 13632
rect 23514 13572 23518 13628
rect 23518 13572 23574 13628
rect 23574 13572 23578 13628
rect 23514 13568 23578 13572
rect 23594 13628 23658 13632
rect 23594 13572 23598 13628
rect 23598 13572 23654 13628
rect 23654 13572 23658 13628
rect 23594 13568 23658 13572
rect 23674 13628 23738 13632
rect 23674 13572 23678 13628
rect 23678 13572 23734 13628
rect 23734 13572 23738 13628
rect 23674 13568 23738 13572
rect 23754 13628 23818 13632
rect 23754 13572 23758 13628
rect 23758 13572 23814 13628
rect 23814 13572 23818 13628
rect 23754 13568 23818 13572
rect 31219 13628 31283 13632
rect 31219 13572 31223 13628
rect 31223 13572 31279 13628
rect 31279 13572 31283 13628
rect 31219 13568 31283 13572
rect 31299 13628 31363 13632
rect 31299 13572 31303 13628
rect 31303 13572 31359 13628
rect 31359 13572 31363 13628
rect 31299 13568 31363 13572
rect 31379 13628 31443 13632
rect 31379 13572 31383 13628
rect 31383 13572 31439 13628
rect 31439 13572 31443 13628
rect 31379 13568 31443 13572
rect 31459 13628 31523 13632
rect 31459 13572 31463 13628
rect 31463 13572 31519 13628
rect 31519 13572 31523 13628
rect 31459 13568 31523 13572
rect 4252 13084 4316 13088
rect 4252 13028 4256 13084
rect 4256 13028 4312 13084
rect 4312 13028 4316 13084
rect 4252 13024 4316 13028
rect 4332 13084 4396 13088
rect 4332 13028 4336 13084
rect 4336 13028 4392 13084
rect 4392 13028 4396 13084
rect 4332 13024 4396 13028
rect 4412 13084 4476 13088
rect 4412 13028 4416 13084
rect 4416 13028 4472 13084
rect 4472 13028 4476 13084
rect 4412 13024 4476 13028
rect 4492 13084 4556 13088
rect 4492 13028 4496 13084
rect 4496 13028 4552 13084
rect 4552 13028 4556 13084
rect 4492 13024 4556 13028
rect 11957 13084 12021 13088
rect 11957 13028 11961 13084
rect 11961 13028 12017 13084
rect 12017 13028 12021 13084
rect 11957 13024 12021 13028
rect 12037 13084 12101 13088
rect 12037 13028 12041 13084
rect 12041 13028 12097 13084
rect 12097 13028 12101 13084
rect 12037 13024 12101 13028
rect 12117 13084 12181 13088
rect 12117 13028 12121 13084
rect 12121 13028 12177 13084
rect 12177 13028 12181 13084
rect 12117 13024 12181 13028
rect 12197 13084 12261 13088
rect 12197 13028 12201 13084
rect 12201 13028 12257 13084
rect 12257 13028 12261 13084
rect 12197 13024 12261 13028
rect 19662 13084 19726 13088
rect 19662 13028 19666 13084
rect 19666 13028 19722 13084
rect 19722 13028 19726 13084
rect 19662 13024 19726 13028
rect 19742 13084 19806 13088
rect 19742 13028 19746 13084
rect 19746 13028 19802 13084
rect 19802 13028 19806 13084
rect 19742 13024 19806 13028
rect 19822 13084 19886 13088
rect 19822 13028 19826 13084
rect 19826 13028 19882 13084
rect 19882 13028 19886 13084
rect 19822 13024 19886 13028
rect 19902 13084 19966 13088
rect 19902 13028 19906 13084
rect 19906 13028 19962 13084
rect 19962 13028 19966 13084
rect 19902 13024 19966 13028
rect 27367 13084 27431 13088
rect 27367 13028 27371 13084
rect 27371 13028 27427 13084
rect 27427 13028 27431 13084
rect 27367 13024 27431 13028
rect 27447 13084 27511 13088
rect 27447 13028 27451 13084
rect 27451 13028 27507 13084
rect 27507 13028 27511 13084
rect 27447 13024 27511 13028
rect 27527 13084 27591 13088
rect 27527 13028 27531 13084
rect 27531 13028 27587 13084
rect 27587 13028 27591 13084
rect 27527 13024 27591 13028
rect 27607 13084 27671 13088
rect 27607 13028 27611 13084
rect 27611 13028 27667 13084
rect 27667 13028 27671 13084
rect 27607 13024 27671 13028
rect 8104 12540 8168 12544
rect 8104 12484 8108 12540
rect 8108 12484 8164 12540
rect 8164 12484 8168 12540
rect 8104 12480 8168 12484
rect 8184 12540 8248 12544
rect 8184 12484 8188 12540
rect 8188 12484 8244 12540
rect 8244 12484 8248 12540
rect 8184 12480 8248 12484
rect 8264 12540 8328 12544
rect 8264 12484 8268 12540
rect 8268 12484 8324 12540
rect 8324 12484 8328 12540
rect 8264 12480 8328 12484
rect 8344 12540 8408 12544
rect 8344 12484 8348 12540
rect 8348 12484 8404 12540
rect 8404 12484 8408 12540
rect 8344 12480 8408 12484
rect 15809 12540 15873 12544
rect 15809 12484 15813 12540
rect 15813 12484 15869 12540
rect 15869 12484 15873 12540
rect 15809 12480 15873 12484
rect 15889 12540 15953 12544
rect 15889 12484 15893 12540
rect 15893 12484 15949 12540
rect 15949 12484 15953 12540
rect 15889 12480 15953 12484
rect 15969 12540 16033 12544
rect 15969 12484 15973 12540
rect 15973 12484 16029 12540
rect 16029 12484 16033 12540
rect 15969 12480 16033 12484
rect 16049 12540 16113 12544
rect 16049 12484 16053 12540
rect 16053 12484 16109 12540
rect 16109 12484 16113 12540
rect 16049 12480 16113 12484
rect 23514 12540 23578 12544
rect 23514 12484 23518 12540
rect 23518 12484 23574 12540
rect 23574 12484 23578 12540
rect 23514 12480 23578 12484
rect 23594 12540 23658 12544
rect 23594 12484 23598 12540
rect 23598 12484 23654 12540
rect 23654 12484 23658 12540
rect 23594 12480 23658 12484
rect 23674 12540 23738 12544
rect 23674 12484 23678 12540
rect 23678 12484 23734 12540
rect 23734 12484 23738 12540
rect 23674 12480 23738 12484
rect 23754 12540 23818 12544
rect 23754 12484 23758 12540
rect 23758 12484 23814 12540
rect 23814 12484 23818 12540
rect 23754 12480 23818 12484
rect 31219 12540 31283 12544
rect 31219 12484 31223 12540
rect 31223 12484 31279 12540
rect 31279 12484 31283 12540
rect 31219 12480 31283 12484
rect 31299 12540 31363 12544
rect 31299 12484 31303 12540
rect 31303 12484 31359 12540
rect 31359 12484 31363 12540
rect 31299 12480 31363 12484
rect 31379 12540 31443 12544
rect 31379 12484 31383 12540
rect 31383 12484 31439 12540
rect 31439 12484 31443 12540
rect 31379 12480 31443 12484
rect 31459 12540 31523 12544
rect 31459 12484 31463 12540
rect 31463 12484 31519 12540
rect 31519 12484 31523 12540
rect 31459 12480 31523 12484
rect 4252 11996 4316 12000
rect 4252 11940 4256 11996
rect 4256 11940 4312 11996
rect 4312 11940 4316 11996
rect 4252 11936 4316 11940
rect 4332 11996 4396 12000
rect 4332 11940 4336 11996
rect 4336 11940 4392 11996
rect 4392 11940 4396 11996
rect 4332 11936 4396 11940
rect 4412 11996 4476 12000
rect 4412 11940 4416 11996
rect 4416 11940 4472 11996
rect 4472 11940 4476 11996
rect 4412 11936 4476 11940
rect 4492 11996 4556 12000
rect 4492 11940 4496 11996
rect 4496 11940 4552 11996
rect 4552 11940 4556 11996
rect 4492 11936 4556 11940
rect 11957 11996 12021 12000
rect 11957 11940 11961 11996
rect 11961 11940 12017 11996
rect 12017 11940 12021 11996
rect 11957 11936 12021 11940
rect 12037 11996 12101 12000
rect 12037 11940 12041 11996
rect 12041 11940 12097 11996
rect 12097 11940 12101 11996
rect 12037 11936 12101 11940
rect 12117 11996 12181 12000
rect 12117 11940 12121 11996
rect 12121 11940 12177 11996
rect 12177 11940 12181 11996
rect 12117 11936 12181 11940
rect 12197 11996 12261 12000
rect 12197 11940 12201 11996
rect 12201 11940 12257 11996
rect 12257 11940 12261 11996
rect 12197 11936 12261 11940
rect 19662 11996 19726 12000
rect 19662 11940 19666 11996
rect 19666 11940 19722 11996
rect 19722 11940 19726 11996
rect 19662 11936 19726 11940
rect 19742 11996 19806 12000
rect 19742 11940 19746 11996
rect 19746 11940 19802 11996
rect 19802 11940 19806 11996
rect 19742 11936 19806 11940
rect 19822 11996 19886 12000
rect 19822 11940 19826 11996
rect 19826 11940 19882 11996
rect 19882 11940 19886 11996
rect 19822 11936 19886 11940
rect 19902 11996 19966 12000
rect 19902 11940 19906 11996
rect 19906 11940 19962 11996
rect 19962 11940 19966 11996
rect 19902 11936 19966 11940
rect 27367 11996 27431 12000
rect 27367 11940 27371 11996
rect 27371 11940 27427 11996
rect 27427 11940 27431 11996
rect 27367 11936 27431 11940
rect 27447 11996 27511 12000
rect 27447 11940 27451 11996
rect 27451 11940 27507 11996
rect 27507 11940 27511 11996
rect 27447 11936 27511 11940
rect 27527 11996 27591 12000
rect 27527 11940 27531 11996
rect 27531 11940 27587 11996
rect 27587 11940 27591 11996
rect 27527 11936 27591 11940
rect 27607 11996 27671 12000
rect 27607 11940 27611 11996
rect 27611 11940 27667 11996
rect 27667 11940 27671 11996
rect 27607 11936 27671 11940
rect 8104 11452 8168 11456
rect 8104 11396 8108 11452
rect 8108 11396 8164 11452
rect 8164 11396 8168 11452
rect 8104 11392 8168 11396
rect 8184 11452 8248 11456
rect 8184 11396 8188 11452
rect 8188 11396 8244 11452
rect 8244 11396 8248 11452
rect 8184 11392 8248 11396
rect 8264 11452 8328 11456
rect 8264 11396 8268 11452
rect 8268 11396 8324 11452
rect 8324 11396 8328 11452
rect 8264 11392 8328 11396
rect 8344 11452 8408 11456
rect 8344 11396 8348 11452
rect 8348 11396 8404 11452
rect 8404 11396 8408 11452
rect 8344 11392 8408 11396
rect 15809 11452 15873 11456
rect 15809 11396 15813 11452
rect 15813 11396 15869 11452
rect 15869 11396 15873 11452
rect 15809 11392 15873 11396
rect 15889 11452 15953 11456
rect 15889 11396 15893 11452
rect 15893 11396 15949 11452
rect 15949 11396 15953 11452
rect 15889 11392 15953 11396
rect 15969 11452 16033 11456
rect 15969 11396 15973 11452
rect 15973 11396 16029 11452
rect 16029 11396 16033 11452
rect 15969 11392 16033 11396
rect 16049 11452 16113 11456
rect 16049 11396 16053 11452
rect 16053 11396 16109 11452
rect 16109 11396 16113 11452
rect 16049 11392 16113 11396
rect 23514 11452 23578 11456
rect 23514 11396 23518 11452
rect 23518 11396 23574 11452
rect 23574 11396 23578 11452
rect 23514 11392 23578 11396
rect 23594 11452 23658 11456
rect 23594 11396 23598 11452
rect 23598 11396 23654 11452
rect 23654 11396 23658 11452
rect 23594 11392 23658 11396
rect 23674 11452 23738 11456
rect 23674 11396 23678 11452
rect 23678 11396 23734 11452
rect 23734 11396 23738 11452
rect 23674 11392 23738 11396
rect 23754 11452 23818 11456
rect 23754 11396 23758 11452
rect 23758 11396 23814 11452
rect 23814 11396 23818 11452
rect 23754 11392 23818 11396
rect 31219 11452 31283 11456
rect 31219 11396 31223 11452
rect 31223 11396 31279 11452
rect 31279 11396 31283 11452
rect 31219 11392 31283 11396
rect 31299 11452 31363 11456
rect 31299 11396 31303 11452
rect 31303 11396 31359 11452
rect 31359 11396 31363 11452
rect 31299 11392 31363 11396
rect 31379 11452 31443 11456
rect 31379 11396 31383 11452
rect 31383 11396 31439 11452
rect 31439 11396 31443 11452
rect 31379 11392 31443 11396
rect 31459 11452 31523 11456
rect 31459 11396 31463 11452
rect 31463 11396 31519 11452
rect 31519 11396 31523 11452
rect 31459 11392 31523 11396
rect 4252 10908 4316 10912
rect 4252 10852 4256 10908
rect 4256 10852 4312 10908
rect 4312 10852 4316 10908
rect 4252 10848 4316 10852
rect 4332 10908 4396 10912
rect 4332 10852 4336 10908
rect 4336 10852 4392 10908
rect 4392 10852 4396 10908
rect 4332 10848 4396 10852
rect 4412 10908 4476 10912
rect 4412 10852 4416 10908
rect 4416 10852 4472 10908
rect 4472 10852 4476 10908
rect 4412 10848 4476 10852
rect 4492 10908 4556 10912
rect 4492 10852 4496 10908
rect 4496 10852 4552 10908
rect 4552 10852 4556 10908
rect 4492 10848 4556 10852
rect 11957 10908 12021 10912
rect 11957 10852 11961 10908
rect 11961 10852 12017 10908
rect 12017 10852 12021 10908
rect 11957 10848 12021 10852
rect 12037 10908 12101 10912
rect 12037 10852 12041 10908
rect 12041 10852 12097 10908
rect 12097 10852 12101 10908
rect 12037 10848 12101 10852
rect 12117 10908 12181 10912
rect 12117 10852 12121 10908
rect 12121 10852 12177 10908
rect 12177 10852 12181 10908
rect 12117 10848 12181 10852
rect 12197 10908 12261 10912
rect 12197 10852 12201 10908
rect 12201 10852 12257 10908
rect 12257 10852 12261 10908
rect 12197 10848 12261 10852
rect 19662 10908 19726 10912
rect 19662 10852 19666 10908
rect 19666 10852 19722 10908
rect 19722 10852 19726 10908
rect 19662 10848 19726 10852
rect 19742 10908 19806 10912
rect 19742 10852 19746 10908
rect 19746 10852 19802 10908
rect 19802 10852 19806 10908
rect 19742 10848 19806 10852
rect 19822 10908 19886 10912
rect 19822 10852 19826 10908
rect 19826 10852 19882 10908
rect 19882 10852 19886 10908
rect 19822 10848 19886 10852
rect 19902 10908 19966 10912
rect 19902 10852 19906 10908
rect 19906 10852 19962 10908
rect 19962 10852 19966 10908
rect 19902 10848 19966 10852
rect 27367 10908 27431 10912
rect 27367 10852 27371 10908
rect 27371 10852 27427 10908
rect 27427 10852 27431 10908
rect 27367 10848 27431 10852
rect 27447 10908 27511 10912
rect 27447 10852 27451 10908
rect 27451 10852 27507 10908
rect 27507 10852 27511 10908
rect 27447 10848 27511 10852
rect 27527 10908 27591 10912
rect 27527 10852 27531 10908
rect 27531 10852 27587 10908
rect 27587 10852 27591 10908
rect 27527 10848 27591 10852
rect 27607 10908 27671 10912
rect 27607 10852 27611 10908
rect 27611 10852 27667 10908
rect 27667 10852 27671 10908
rect 27607 10848 27671 10852
rect 8104 10364 8168 10368
rect 8104 10308 8108 10364
rect 8108 10308 8164 10364
rect 8164 10308 8168 10364
rect 8104 10304 8168 10308
rect 8184 10364 8248 10368
rect 8184 10308 8188 10364
rect 8188 10308 8244 10364
rect 8244 10308 8248 10364
rect 8184 10304 8248 10308
rect 8264 10364 8328 10368
rect 8264 10308 8268 10364
rect 8268 10308 8324 10364
rect 8324 10308 8328 10364
rect 8264 10304 8328 10308
rect 8344 10364 8408 10368
rect 8344 10308 8348 10364
rect 8348 10308 8404 10364
rect 8404 10308 8408 10364
rect 8344 10304 8408 10308
rect 15809 10364 15873 10368
rect 15809 10308 15813 10364
rect 15813 10308 15869 10364
rect 15869 10308 15873 10364
rect 15809 10304 15873 10308
rect 15889 10364 15953 10368
rect 15889 10308 15893 10364
rect 15893 10308 15949 10364
rect 15949 10308 15953 10364
rect 15889 10304 15953 10308
rect 15969 10364 16033 10368
rect 15969 10308 15973 10364
rect 15973 10308 16029 10364
rect 16029 10308 16033 10364
rect 15969 10304 16033 10308
rect 16049 10364 16113 10368
rect 16049 10308 16053 10364
rect 16053 10308 16109 10364
rect 16109 10308 16113 10364
rect 16049 10304 16113 10308
rect 23514 10364 23578 10368
rect 23514 10308 23518 10364
rect 23518 10308 23574 10364
rect 23574 10308 23578 10364
rect 23514 10304 23578 10308
rect 23594 10364 23658 10368
rect 23594 10308 23598 10364
rect 23598 10308 23654 10364
rect 23654 10308 23658 10364
rect 23594 10304 23658 10308
rect 23674 10364 23738 10368
rect 23674 10308 23678 10364
rect 23678 10308 23734 10364
rect 23734 10308 23738 10364
rect 23674 10304 23738 10308
rect 23754 10364 23818 10368
rect 23754 10308 23758 10364
rect 23758 10308 23814 10364
rect 23814 10308 23818 10364
rect 23754 10304 23818 10308
rect 31219 10364 31283 10368
rect 31219 10308 31223 10364
rect 31223 10308 31279 10364
rect 31279 10308 31283 10364
rect 31219 10304 31283 10308
rect 31299 10364 31363 10368
rect 31299 10308 31303 10364
rect 31303 10308 31359 10364
rect 31359 10308 31363 10364
rect 31299 10304 31363 10308
rect 31379 10364 31443 10368
rect 31379 10308 31383 10364
rect 31383 10308 31439 10364
rect 31439 10308 31443 10364
rect 31379 10304 31443 10308
rect 31459 10364 31523 10368
rect 31459 10308 31463 10364
rect 31463 10308 31519 10364
rect 31519 10308 31523 10364
rect 31459 10304 31523 10308
rect 4252 9820 4316 9824
rect 4252 9764 4256 9820
rect 4256 9764 4312 9820
rect 4312 9764 4316 9820
rect 4252 9760 4316 9764
rect 4332 9820 4396 9824
rect 4332 9764 4336 9820
rect 4336 9764 4392 9820
rect 4392 9764 4396 9820
rect 4332 9760 4396 9764
rect 4412 9820 4476 9824
rect 4412 9764 4416 9820
rect 4416 9764 4472 9820
rect 4472 9764 4476 9820
rect 4412 9760 4476 9764
rect 4492 9820 4556 9824
rect 4492 9764 4496 9820
rect 4496 9764 4552 9820
rect 4552 9764 4556 9820
rect 4492 9760 4556 9764
rect 11957 9820 12021 9824
rect 11957 9764 11961 9820
rect 11961 9764 12017 9820
rect 12017 9764 12021 9820
rect 11957 9760 12021 9764
rect 12037 9820 12101 9824
rect 12037 9764 12041 9820
rect 12041 9764 12097 9820
rect 12097 9764 12101 9820
rect 12037 9760 12101 9764
rect 12117 9820 12181 9824
rect 12117 9764 12121 9820
rect 12121 9764 12177 9820
rect 12177 9764 12181 9820
rect 12117 9760 12181 9764
rect 12197 9820 12261 9824
rect 12197 9764 12201 9820
rect 12201 9764 12257 9820
rect 12257 9764 12261 9820
rect 12197 9760 12261 9764
rect 19662 9820 19726 9824
rect 19662 9764 19666 9820
rect 19666 9764 19722 9820
rect 19722 9764 19726 9820
rect 19662 9760 19726 9764
rect 19742 9820 19806 9824
rect 19742 9764 19746 9820
rect 19746 9764 19802 9820
rect 19802 9764 19806 9820
rect 19742 9760 19806 9764
rect 19822 9820 19886 9824
rect 19822 9764 19826 9820
rect 19826 9764 19882 9820
rect 19882 9764 19886 9820
rect 19822 9760 19886 9764
rect 19902 9820 19966 9824
rect 19902 9764 19906 9820
rect 19906 9764 19962 9820
rect 19962 9764 19966 9820
rect 19902 9760 19966 9764
rect 27367 9820 27431 9824
rect 27367 9764 27371 9820
rect 27371 9764 27427 9820
rect 27427 9764 27431 9820
rect 27367 9760 27431 9764
rect 27447 9820 27511 9824
rect 27447 9764 27451 9820
rect 27451 9764 27507 9820
rect 27507 9764 27511 9820
rect 27447 9760 27511 9764
rect 27527 9820 27591 9824
rect 27527 9764 27531 9820
rect 27531 9764 27587 9820
rect 27587 9764 27591 9820
rect 27527 9760 27591 9764
rect 27607 9820 27671 9824
rect 27607 9764 27611 9820
rect 27611 9764 27667 9820
rect 27667 9764 27671 9820
rect 27607 9760 27671 9764
rect 8104 9276 8168 9280
rect 8104 9220 8108 9276
rect 8108 9220 8164 9276
rect 8164 9220 8168 9276
rect 8104 9216 8168 9220
rect 8184 9276 8248 9280
rect 8184 9220 8188 9276
rect 8188 9220 8244 9276
rect 8244 9220 8248 9276
rect 8184 9216 8248 9220
rect 8264 9276 8328 9280
rect 8264 9220 8268 9276
rect 8268 9220 8324 9276
rect 8324 9220 8328 9276
rect 8264 9216 8328 9220
rect 8344 9276 8408 9280
rect 8344 9220 8348 9276
rect 8348 9220 8404 9276
rect 8404 9220 8408 9276
rect 8344 9216 8408 9220
rect 15809 9276 15873 9280
rect 15809 9220 15813 9276
rect 15813 9220 15869 9276
rect 15869 9220 15873 9276
rect 15809 9216 15873 9220
rect 15889 9276 15953 9280
rect 15889 9220 15893 9276
rect 15893 9220 15949 9276
rect 15949 9220 15953 9276
rect 15889 9216 15953 9220
rect 15969 9276 16033 9280
rect 15969 9220 15973 9276
rect 15973 9220 16029 9276
rect 16029 9220 16033 9276
rect 15969 9216 16033 9220
rect 16049 9276 16113 9280
rect 16049 9220 16053 9276
rect 16053 9220 16109 9276
rect 16109 9220 16113 9276
rect 16049 9216 16113 9220
rect 23514 9276 23578 9280
rect 23514 9220 23518 9276
rect 23518 9220 23574 9276
rect 23574 9220 23578 9276
rect 23514 9216 23578 9220
rect 23594 9276 23658 9280
rect 23594 9220 23598 9276
rect 23598 9220 23654 9276
rect 23654 9220 23658 9276
rect 23594 9216 23658 9220
rect 23674 9276 23738 9280
rect 23674 9220 23678 9276
rect 23678 9220 23734 9276
rect 23734 9220 23738 9276
rect 23674 9216 23738 9220
rect 23754 9276 23818 9280
rect 23754 9220 23758 9276
rect 23758 9220 23814 9276
rect 23814 9220 23818 9276
rect 23754 9216 23818 9220
rect 31219 9276 31283 9280
rect 31219 9220 31223 9276
rect 31223 9220 31279 9276
rect 31279 9220 31283 9276
rect 31219 9216 31283 9220
rect 31299 9276 31363 9280
rect 31299 9220 31303 9276
rect 31303 9220 31359 9276
rect 31359 9220 31363 9276
rect 31299 9216 31363 9220
rect 31379 9276 31443 9280
rect 31379 9220 31383 9276
rect 31383 9220 31439 9276
rect 31439 9220 31443 9276
rect 31379 9216 31443 9220
rect 31459 9276 31523 9280
rect 31459 9220 31463 9276
rect 31463 9220 31519 9276
rect 31519 9220 31523 9276
rect 31459 9216 31523 9220
rect 4252 8732 4316 8736
rect 4252 8676 4256 8732
rect 4256 8676 4312 8732
rect 4312 8676 4316 8732
rect 4252 8672 4316 8676
rect 4332 8732 4396 8736
rect 4332 8676 4336 8732
rect 4336 8676 4392 8732
rect 4392 8676 4396 8732
rect 4332 8672 4396 8676
rect 4412 8732 4476 8736
rect 4412 8676 4416 8732
rect 4416 8676 4472 8732
rect 4472 8676 4476 8732
rect 4412 8672 4476 8676
rect 4492 8732 4556 8736
rect 4492 8676 4496 8732
rect 4496 8676 4552 8732
rect 4552 8676 4556 8732
rect 4492 8672 4556 8676
rect 11957 8732 12021 8736
rect 11957 8676 11961 8732
rect 11961 8676 12017 8732
rect 12017 8676 12021 8732
rect 11957 8672 12021 8676
rect 12037 8732 12101 8736
rect 12037 8676 12041 8732
rect 12041 8676 12097 8732
rect 12097 8676 12101 8732
rect 12037 8672 12101 8676
rect 12117 8732 12181 8736
rect 12117 8676 12121 8732
rect 12121 8676 12177 8732
rect 12177 8676 12181 8732
rect 12117 8672 12181 8676
rect 12197 8732 12261 8736
rect 12197 8676 12201 8732
rect 12201 8676 12257 8732
rect 12257 8676 12261 8732
rect 12197 8672 12261 8676
rect 19662 8732 19726 8736
rect 19662 8676 19666 8732
rect 19666 8676 19722 8732
rect 19722 8676 19726 8732
rect 19662 8672 19726 8676
rect 19742 8732 19806 8736
rect 19742 8676 19746 8732
rect 19746 8676 19802 8732
rect 19802 8676 19806 8732
rect 19742 8672 19806 8676
rect 19822 8732 19886 8736
rect 19822 8676 19826 8732
rect 19826 8676 19882 8732
rect 19882 8676 19886 8732
rect 19822 8672 19886 8676
rect 19902 8732 19966 8736
rect 19902 8676 19906 8732
rect 19906 8676 19962 8732
rect 19962 8676 19966 8732
rect 19902 8672 19966 8676
rect 27367 8732 27431 8736
rect 27367 8676 27371 8732
rect 27371 8676 27427 8732
rect 27427 8676 27431 8732
rect 27367 8672 27431 8676
rect 27447 8732 27511 8736
rect 27447 8676 27451 8732
rect 27451 8676 27507 8732
rect 27507 8676 27511 8732
rect 27447 8672 27511 8676
rect 27527 8732 27591 8736
rect 27527 8676 27531 8732
rect 27531 8676 27587 8732
rect 27587 8676 27591 8732
rect 27527 8672 27591 8676
rect 27607 8732 27671 8736
rect 27607 8676 27611 8732
rect 27611 8676 27667 8732
rect 27667 8676 27671 8732
rect 27607 8672 27671 8676
rect 8104 8188 8168 8192
rect 8104 8132 8108 8188
rect 8108 8132 8164 8188
rect 8164 8132 8168 8188
rect 8104 8128 8168 8132
rect 8184 8188 8248 8192
rect 8184 8132 8188 8188
rect 8188 8132 8244 8188
rect 8244 8132 8248 8188
rect 8184 8128 8248 8132
rect 8264 8188 8328 8192
rect 8264 8132 8268 8188
rect 8268 8132 8324 8188
rect 8324 8132 8328 8188
rect 8264 8128 8328 8132
rect 8344 8188 8408 8192
rect 8344 8132 8348 8188
rect 8348 8132 8404 8188
rect 8404 8132 8408 8188
rect 8344 8128 8408 8132
rect 15809 8188 15873 8192
rect 15809 8132 15813 8188
rect 15813 8132 15869 8188
rect 15869 8132 15873 8188
rect 15809 8128 15873 8132
rect 15889 8188 15953 8192
rect 15889 8132 15893 8188
rect 15893 8132 15949 8188
rect 15949 8132 15953 8188
rect 15889 8128 15953 8132
rect 15969 8188 16033 8192
rect 15969 8132 15973 8188
rect 15973 8132 16029 8188
rect 16029 8132 16033 8188
rect 15969 8128 16033 8132
rect 16049 8188 16113 8192
rect 16049 8132 16053 8188
rect 16053 8132 16109 8188
rect 16109 8132 16113 8188
rect 16049 8128 16113 8132
rect 23514 8188 23578 8192
rect 23514 8132 23518 8188
rect 23518 8132 23574 8188
rect 23574 8132 23578 8188
rect 23514 8128 23578 8132
rect 23594 8188 23658 8192
rect 23594 8132 23598 8188
rect 23598 8132 23654 8188
rect 23654 8132 23658 8188
rect 23594 8128 23658 8132
rect 23674 8188 23738 8192
rect 23674 8132 23678 8188
rect 23678 8132 23734 8188
rect 23734 8132 23738 8188
rect 23674 8128 23738 8132
rect 23754 8188 23818 8192
rect 23754 8132 23758 8188
rect 23758 8132 23814 8188
rect 23814 8132 23818 8188
rect 23754 8128 23818 8132
rect 31219 8188 31283 8192
rect 31219 8132 31223 8188
rect 31223 8132 31279 8188
rect 31279 8132 31283 8188
rect 31219 8128 31283 8132
rect 31299 8188 31363 8192
rect 31299 8132 31303 8188
rect 31303 8132 31359 8188
rect 31359 8132 31363 8188
rect 31299 8128 31363 8132
rect 31379 8188 31443 8192
rect 31379 8132 31383 8188
rect 31383 8132 31439 8188
rect 31439 8132 31443 8188
rect 31379 8128 31443 8132
rect 31459 8188 31523 8192
rect 31459 8132 31463 8188
rect 31463 8132 31519 8188
rect 31519 8132 31523 8188
rect 31459 8128 31523 8132
rect 4252 7644 4316 7648
rect 4252 7588 4256 7644
rect 4256 7588 4312 7644
rect 4312 7588 4316 7644
rect 4252 7584 4316 7588
rect 4332 7644 4396 7648
rect 4332 7588 4336 7644
rect 4336 7588 4392 7644
rect 4392 7588 4396 7644
rect 4332 7584 4396 7588
rect 4412 7644 4476 7648
rect 4412 7588 4416 7644
rect 4416 7588 4472 7644
rect 4472 7588 4476 7644
rect 4412 7584 4476 7588
rect 4492 7644 4556 7648
rect 4492 7588 4496 7644
rect 4496 7588 4552 7644
rect 4552 7588 4556 7644
rect 4492 7584 4556 7588
rect 11957 7644 12021 7648
rect 11957 7588 11961 7644
rect 11961 7588 12017 7644
rect 12017 7588 12021 7644
rect 11957 7584 12021 7588
rect 12037 7644 12101 7648
rect 12037 7588 12041 7644
rect 12041 7588 12097 7644
rect 12097 7588 12101 7644
rect 12037 7584 12101 7588
rect 12117 7644 12181 7648
rect 12117 7588 12121 7644
rect 12121 7588 12177 7644
rect 12177 7588 12181 7644
rect 12117 7584 12181 7588
rect 12197 7644 12261 7648
rect 12197 7588 12201 7644
rect 12201 7588 12257 7644
rect 12257 7588 12261 7644
rect 12197 7584 12261 7588
rect 19662 7644 19726 7648
rect 19662 7588 19666 7644
rect 19666 7588 19722 7644
rect 19722 7588 19726 7644
rect 19662 7584 19726 7588
rect 19742 7644 19806 7648
rect 19742 7588 19746 7644
rect 19746 7588 19802 7644
rect 19802 7588 19806 7644
rect 19742 7584 19806 7588
rect 19822 7644 19886 7648
rect 19822 7588 19826 7644
rect 19826 7588 19882 7644
rect 19882 7588 19886 7644
rect 19822 7584 19886 7588
rect 19902 7644 19966 7648
rect 19902 7588 19906 7644
rect 19906 7588 19962 7644
rect 19962 7588 19966 7644
rect 19902 7584 19966 7588
rect 27367 7644 27431 7648
rect 27367 7588 27371 7644
rect 27371 7588 27427 7644
rect 27427 7588 27431 7644
rect 27367 7584 27431 7588
rect 27447 7644 27511 7648
rect 27447 7588 27451 7644
rect 27451 7588 27507 7644
rect 27507 7588 27511 7644
rect 27447 7584 27511 7588
rect 27527 7644 27591 7648
rect 27527 7588 27531 7644
rect 27531 7588 27587 7644
rect 27587 7588 27591 7644
rect 27527 7584 27591 7588
rect 27607 7644 27671 7648
rect 27607 7588 27611 7644
rect 27611 7588 27667 7644
rect 27667 7588 27671 7644
rect 27607 7584 27671 7588
rect 8104 7100 8168 7104
rect 8104 7044 8108 7100
rect 8108 7044 8164 7100
rect 8164 7044 8168 7100
rect 8104 7040 8168 7044
rect 8184 7100 8248 7104
rect 8184 7044 8188 7100
rect 8188 7044 8244 7100
rect 8244 7044 8248 7100
rect 8184 7040 8248 7044
rect 8264 7100 8328 7104
rect 8264 7044 8268 7100
rect 8268 7044 8324 7100
rect 8324 7044 8328 7100
rect 8264 7040 8328 7044
rect 8344 7100 8408 7104
rect 8344 7044 8348 7100
rect 8348 7044 8404 7100
rect 8404 7044 8408 7100
rect 8344 7040 8408 7044
rect 15809 7100 15873 7104
rect 15809 7044 15813 7100
rect 15813 7044 15869 7100
rect 15869 7044 15873 7100
rect 15809 7040 15873 7044
rect 15889 7100 15953 7104
rect 15889 7044 15893 7100
rect 15893 7044 15949 7100
rect 15949 7044 15953 7100
rect 15889 7040 15953 7044
rect 15969 7100 16033 7104
rect 15969 7044 15973 7100
rect 15973 7044 16029 7100
rect 16029 7044 16033 7100
rect 15969 7040 16033 7044
rect 16049 7100 16113 7104
rect 16049 7044 16053 7100
rect 16053 7044 16109 7100
rect 16109 7044 16113 7100
rect 16049 7040 16113 7044
rect 23514 7100 23578 7104
rect 23514 7044 23518 7100
rect 23518 7044 23574 7100
rect 23574 7044 23578 7100
rect 23514 7040 23578 7044
rect 23594 7100 23658 7104
rect 23594 7044 23598 7100
rect 23598 7044 23654 7100
rect 23654 7044 23658 7100
rect 23594 7040 23658 7044
rect 23674 7100 23738 7104
rect 23674 7044 23678 7100
rect 23678 7044 23734 7100
rect 23734 7044 23738 7100
rect 23674 7040 23738 7044
rect 23754 7100 23818 7104
rect 23754 7044 23758 7100
rect 23758 7044 23814 7100
rect 23814 7044 23818 7100
rect 23754 7040 23818 7044
rect 31219 7100 31283 7104
rect 31219 7044 31223 7100
rect 31223 7044 31279 7100
rect 31279 7044 31283 7100
rect 31219 7040 31283 7044
rect 31299 7100 31363 7104
rect 31299 7044 31303 7100
rect 31303 7044 31359 7100
rect 31359 7044 31363 7100
rect 31299 7040 31363 7044
rect 31379 7100 31443 7104
rect 31379 7044 31383 7100
rect 31383 7044 31439 7100
rect 31439 7044 31443 7100
rect 31379 7040 31443 7044
rect 31459 7100 31523 7104
rect 31459 7044 31463 7100
rect 31463 7044 31519 7100
rect 31519 7044 31523 7100
rect 31459 7040 31523 7044
rect 4252 6556 4316 6560
rect 4252 6500 4256 6556
rect 4256 6500 4312 6556
rect 4312 6500 4316 6556
rect 4252 6496 4316 6500
rect 4332 6556 4396 6560
rect 4332 6500 4336 6556
rect 4336 6500 4392 6556
rect 4392 6500 4396 6556
rect 4332 6496 4396 6500
rect 4412 6556 4476 6560
rect 4412 6500 4416 6556
rect 4416 6500 4472 6556
rect 4472 6500 4476 6556
rect 4412 6496 4476 6500
rect 4492 6556 4556 6560
rect 4492 6500 4496 6556
rect 4496 6500 4552 6556
rect 4552 6500 4556 6556
rect 4492 6496 4556 6500
rect 11957 6556 12021 6560
rect 11957 6500 11961 6556
rect 11961 6500 12017 6556
rect 12017 6500 12021 6556
rect 11957 6496 12021 6500
rect 12037 6556 12101 6560
rect 12037 6500 12041 6556
rect 12041 6500 12097 6556
rect 12097 6500 12101 6556
rect 12037 6496 12101 6500
rect 12117 6556 12181 6560
rect 12117 6500 12121 6556
rect 12121 6500 12177 6556
rect 12177 6500 12181 6556
rect 12117 6496 12181 6500
rect 12197 6556 12261 6560
rect 12197 6500 12201 6556
rect 12201 6500 12257 6556
rect 12257 6500 12261 6556
rect 12197 6496 12261 6500
rect 19662 6556 19726 6560
rect 19662 6500 19666 6556
rect 19666 6500 19722 6556
rect 19722 6500 19726 6556
rect 19662 6496 19726 6500
rect 19742 6556 19806 6560
rect 19742 6500 19746 6556
rect 19746 6500 19802 6556
rect 19802 6500 19806 6556
rect 19742 6496 19806 6500
rect 19822 6556 19886 6560
rect 19822 6500 19826 6556
rect 19826 6500 19882 6556
rect 19882 6500 19886 6556
rect 19822 6496 19886 6500
rect 19902 6556 19966 6560
rect 19902 6500 19906 6556
rect 19906 6500 19962 6556
rect 19962 6500 19966 6556
rect 19902 6496 19966 6500
rect 27367 6556 27431 6560
rect 27367 6500 27371 6556
rect 27371 6500 27427 6556
rect 27427 6500 27431 6556
rect 27367 6496 27431 6500
rect 27447 6556 27511 6560
rect 27447 6500 27451 6556
rect 27451 6500 27507 6556
rect 27507 6500 27511 6556
rect 27447 6496 27511 6500
rect 27527 6556 27591 6560
rect 27527 6500 27531 6556
rect 27531 6500 27587 6556
rect 27587 6500 27591 6556
rect 27527 6496 27591 6500
rect 27607 6556 27671 6560
rect 27607 6500 27611 6556
rect 27611 6500 27667 6556
rect 27667 6500 27671 6556
rect 27607 6496 27671 6500
rect 8104 6012 8168 6016
rect 8104 5956 8108 6012
rect 8108 5956 8164 6012
rect 8164 5956 8168 6012
rect 8104 5952 8168 5956
rect 8184 6012 8248 6016
rect 8184 5956 8188 6012
rect 8188 5956 8244 6012
rect 8244 5956 8248 6012
rect 8184 5952 8248 5956
rect 8264 6012 8328 6016
rect 8264 5956 8268 6012
rect 8268 5956 8324 6012
rect 8324 5956 8328 6012
rect 8264 5952 8328 5956
rect 8344 6012 8408 6016
rect 8344 5956 8348 6012
rect 8348 5956 8404 6012
rect 8404 5956 8408 6012
rect 8344 5952 8408 5956
rect 15809 6012 15873 6016
rect 15809 5956 15813 6012
rect 15813 5956 15869 6012
rect 15869 5956 15873 6012
rect 15809 5952 15873 5956
rect 15889 6012 15953 6016
rect 15889 5956 15893 6012
rect 15893 5956 15949 6012
rect 15949 5956 15953 6012
rect 15889 5952 15953 5956
rect 15969 6012 16033 6016
rect 15969 5956 15973 6012
rect 15973 5956 16029 6012
rect 16029 5956 16033 6012
rect 15969 5952 16033 5956
rect 16049 6012 16113 6016
rect 16049 5956 16053 6012
rect 16053 5956 16109 6012
rect 16109 5956 16113 6012
rect 16049 5952 16113 5956
rect 23514 6012 23578 6016
rect 23514 5956 23518 6012
rect 23518 5956 23574 6012
rect 23574 5956 23578 6012
rect 23514 5952 23578 5956
rect 23594 6012 23658 6016
rect 23594 5956 23598 6012
rect 23598 5956 23654 6012
rect 23654 5956 23658 6012
rect 23594 5952 23658 5956
rect 23674 6012 23738 6016
rect 23674 5956 23678 6012
rect 23678 5956 23734 6012
rect 23734 5956 23738 6012
rect 23674 5952 23738 5956
rect 23754 6012 23818 6016
rect 23754 5956 23758 6012
rect 23758 5956 23814 6012
rect 23814 5956 23818 6012
rect 23754 5952 23818 5956
rect 31219 6012 31283 6016
rect 31219 5956 31223 6012
rect 31223 5956 31279 6012
rect 31279 5956 31283 6012
rect 31219 5952 31283 5956
rect 31299 6012 31363 6016
rect 31299 5956 31303 6012
rect 31303 5956 31359 6012
rect 31359 5956 31363 6012
rect 31299 5952 31363 5956
rect 31379 6012 31443 6016
rect 31379 5956 31383 6012
rect 31383 5956 31439 6012
rect 31439 5956 31443 6012
rect 31379 5952 31443 5956
rect 31459 6012 31523 6016
rect 31459 5956 31463 6012
rect 31463 5956 31519 6012
rect 31519 5956 31523 6012
rect 31459 5952 31523 5956
rect 4252 5468 4316 5472
rect 4252 5412 4256 5468
rect 4256 5412 4312 5468
rect 4312 5412 4316 5468
rect 4252 5408 4316 5412
rect 4332 5468 4396 5472
rect 4332 5412 4336 5468
rect 4336 5412 4392 5468
rect 4392 5412 4396 5468
rect 4332 5408 4396 5412
rect 4412 5468 4476 5472
rect 4412 5412 4416 5468
rect 4416 5412 4472 5468
rect 4472 5412 4476 5468
rect 4412 5408 4476 5412
rect 4492 5468 4556 5472
rect 4492 5412 4496 5468
rect 4496 5412 4552 5468
rect 4552 5412 4556 5468
rect 4492 5408 4556 5412
rect 11957 5468 12021 5472
rect 11957 5412 11961 5468
rect 11961 5412 12017 5468
rect 12017 5412 12021 5468
rect 11957 5408 12021 5412
rect 12037 5468 12101 5472
rect 12037 5412 12041 5468
rect 12041 5412 12097 5468
rect 12097 5412 12101 5468
rect 12037 5408 12101 5412
rect 12117 5468 12181 5472
rect 12117 5412 12121 5468
rect 12121 5412 12177 5468
rect 12177 5412 12181 5468
rect 12117 5408 12181 5412
rect 12197 5468 12261 5472
rect 12197 5412 12201 5468
rect 12201 5412 12257 5468
rect 12257 5412 12261 5468
rect 12197 5408 12261 5412
rect 19662 5468 19726 5472
rect 19662 5412 19666 5468
rect 19666 5412 19722 5468
rect 19722 5412 19726 5468
rect 19662 5408 19726 5412
rect 19742 5468 19806 5472
rect 19742 5412 19746 5468
rect 19746 5412 19802 5468
rect 19802 5412 19806 5468
rect 19742 5408 19806 5412
rect 19822 5468 19886 5472
rect 19822 5412 19826 5468
rect 19826 5412 19882 5468
rect 19882 5412 19886 5468
rect 19822 5408 19886 5412
rect 19902 5468 19966 5472
rect 19902 5412 19906 5468
rect 19906 5412 19962 5468
rect 19962 5412 19966 5468
rect 19902 5408 19966 5412
rect 27367 5468 27431 5472
rect 27367 5412 27371 5468
rect 27371 5412 27427 5468
rect 27427 5412 27431 5468
rect 27367 5408 27431 5412
rect 27447 5468 27511 5472
rect 27447 5412 27451 5468
rect 27451 5412 27507 5468
rect 27507 5412 27511 5468
rect 27447 5408 27511 5412
rect 27527 5468 27591 5472
rect 27527 5412 27531 5468
rect 27531 5412 27587 5468
rect 27587 5412 27591 5468
rect 27527 5408 27591 5412
rect 27607 5468 27671 5472
rect 27607 5412 27611 5468
rect 27611 5412 27667 5468
rect 27667 5412 27671 5468
rect 27607 5408 27671 5412
rect 8104 4924 8168 4928
rect 8104 4868 8108 4924
rect 8108 4868 8164 4924
rect 8164 4868 8168 4924
rect 8104 4864 8168 4868
rect 8184 4924 8248 4928
rect 8184 4868 8188 4924
rect 8188 4868 8244 4924
rect 8244 4868 8248 4924
rect 8184 4864 8248 4868
rect 8264 4924 8328 4928
rect 8264 4868 8268 4924
rect 8268 4868 8324 4924
rect 8324 4868 8328 4924
rect 8264 4864 8328 4868
rect 8344 4924 8408 4928
rect 8344 4868 8348 4924
rect 8348 4868 8404 4924
rect 8404 4868 8408 4924
rect 8344 4864 8408 4868
rect 15809 4924 15873 4928
rect 15809 4868 15813 4924
rect 15813 4868 15869 4924
rect 15869 4868 15873 4924
rect 15809 4864 15873 4868
rect 15889 4924 15953 4928
rect 15889 4868 15893 4924
rect 15893 4868 15949 4924
rect 15949 4868 15953 4924
rect 15889 4864 15953 4868
rect 15969 4924 16033 4928
rect 15969 4868 15973 4924
rect 15973 4868 16029 4924
rect 16029 4868 16033 4924
rect 15969 4864 16033 4868
rect 16049 4924 16113 4928
rect 16049 4868 16053 4924
rect 16053 4868 16109 4924
rect 16109 4868 16113 4924
rect 16049 4864 16113 4868
rect 23514 4924 23578 4928
rect 23514 4868 23518 4924
rect 23518 4868 23574 4924
rect 23574 4868 23578 4924
rect 23514 4864 23578 4868
rect 23594 4924 23658 4928
rect 23594 4868 23598 4924
rect 23598 4868 23654 4924
rect 23654 4868 23658 4924
rect 23594 4864 23658 4868
rect 23674 4924 23738 4928
rect 23674 4868 23678 4924
rect 23678 4868 23734 4924
rect 23734 4868 23738 4924
rect 23674 4864 23738 4868
rect 23754 4924 23818 4928
rect 23754 4868 23758 4924
rect 23758 4868 23814 4924
rect 23814 4868 23818 4924
rect 23754 4864 23818 4868
rect 31219 4924 31283 4928
rect 31219 4868 31223 4924
rect 31223 4868 31279 4924
rect 31279 4868 31283 4924
rect 31219 4864 31283 4868
rect 31299 4924 31363 4928
rect 31299 4868 31303 4924
rect 31303 4868 31359 4924
rect 31359 4868 31363 4924
rect 31299 4864 31363 4868
rect 31379 4924 31443 4928
rect 31379 4868 31383 4924
rect 31383 4868 31439 4924
rect 31439 4868 31443 4924
rect 31379 4864 31443 4868
rect 31459 4924 31523 4928
rect 31459 4868 31463 4924
rect 31463 4868 31519 4924
rect 31519 4868 31523 4924
rect 31459 4864 31523 4868
rect 4252 4380 4316 4384
rect 4252 4324 4256 4380
rect 4256 4324 4312 4380
rect 4312 4324 4316 4380
rect 4252 4320 4316 4324
rect 4332 4380 4396 4384
rect 4332 4324 4336 4380
rect 4336 4324 4392 4380
rect 4392 4324 4396 4380
rect 4332 4320 4396 4324
rect 4412 4380 4476 4384
rect 4412 4324 4416 4380
rect 4416 4324 4472 4380
rect 4472 4324 4476 4380
rect 4412 4320 4476 4324
rect 4492 4380 4556 4384
rect 4492 4324 4496 4380
rect 4496 4324 4552 4380
rect 4552 4324 4556 4380
rect 4492 4320 4556 4324
rect 11957 4380 12021 4384
rect 11957 4324 11961 4380
rect 11961 4324 12017 4380
rect 12017 4324 12021 4380
rect 11957 4320 12021 4324
rect 12037 4380 12101 4384
rect 12037 4324 12041 4380
rect 12041 4324 12097 4380
rect 12097 4324 12101 4380
rect 12037 4320 12101 4324
rect 12117 4380 12181 4384
rect 12117 4324 12121 4380
rect 12121 4324 12177 4380
rect 12177 4324 12181 4380
rect 12117 4320 12181 4324
rect 12197 4380 12261 4384
rect 12197 4324 12201 4380
rect 12201 4324 12257 4380
rect 12257 4324 12261 4380
rect 12197 4320 12261 4324
rect 19662 4380 19726 4384
rect 19662 4324 19666 4380
rect 19666 4324 19722 4380
rect 19722 4324 19726 4380
rect 19662 4320 19726 4324
rect 19742 4380 19806 4384
rect 19742 4324 19746 4380
rect 19746 4324 19802 4380
rect 19802 4324 19806 4380
rect 19742 4320 19806 4324
rect 19822 4380 19886 4384
rect 19822 4324 19826 4380
rect 19826 4324 19882 4380
rect 19882 4324 19886 4380
rect 19822 4320 19886 4324
rect 19902 4380 19966 4384
rect 19902 4324 19906 4380
rect 19906 4324 19962 4380
rect 19962 4324 19966 4380
rect 19902 4320 19966 4324
rect 27367 4380 27431 4384
rect 27367 4324 27371 4380
rect 27371 4324 27427 4380
rect 27427 4324 27431 4380
rect 27367 4320 27431 4324
rect 27447 4380 27511 4384
rect 27447 4324 27451 4380
rect 27451 4324 27507 4380
rect 27507 4324 27511 4380
rect 27447 4320 27511 4324
rect 27527 4380 27591 4384
rect 27527 4324 27531 4380
rect 27531 4324 27587 4380
rect 27587 4324 27591 4380
rect 27527 4320 27591 4324
rect 27607 4380 27671 4384
rect 27607 4324 27611 4380
rect 27611 4324 27667 4380
rect 27667 4324 27671 4380
rect 27607 4320 27671 4324
rect 8104 3836 8168 3840
rect 8104 3780 8108 3836
rect 8108 3780 8164 3836
rect 8164 3780 8168 3836
rect 8104 3776 8168 3780
rect 8184 3836 8248 3840
rect 8184 3780 8188 3836
rect 8188 3780 8244 3836
rect 8244 3780 8248 3836
rect 8184 3776 8248 3780
rect 8264 3836 8328 3840
rect 8264 3780 8268 3836
rect 8268 3780 8324 3836
rect 8324 3780 8328 3836
rect 8264 3776 8328 3780
rect 8344 3836 8408 3840
rect 8344 3780 8348 3836
rect 8348 3780 8404 3836
rect 8404 3780 8408 3836
rect 8344 3776 8408 3780
rect 15809 3836 15873 3840
rect 15809 3780 15813 3836
rect 15813 3780 15869 3836
rect 15869 3780 15873 3836
rect 15809 3776 15873 3780
rect 15889 3836 15953 3840
rect 15889 3780 15893 3836
rect 15893 3780 15949 3836
rect 15949 3780 15953 3836
rect 15889 3776 15953 3780
rect 15969 3836 16033 3840
rect 15969 3780 15973 3836
rect 15973 3780 16029 3836
rect 16029 3780 16033 3836
rect 15969 3776 16033 3780
rect 16049 3836 16113 3840
rect 16049 3780 16053 3836
rect 16053 3780 16109 3836
rect 16109 3780 16113 3836
rect 16049 3776 16113 3780
rect 23514 3836 23578 3840
rect 23514 3780 23518 3836
rect 23518 3780 23574 3836
rect 23574 3780 23578 3836
rect 23514 3776 23578 3780
rect 23594 3836 23658 3840
rect 23594 3780 23598 3836
rect 23598 3780 23654 3836
rect 23654 3780 23658 3836
rect 23594 3776 23658 3780
rect 23674 3836 23738 3840
rect 23674 3780 23678 3836
rect 23678 3780 23734 3836
rect 23734 3780 23738 3836
rect 23674 3776 23738 3780
rect 23754 3836 23818 3840
rect 23754 3780 23758 3836
rect 23758 3780 23814 3836
rect 23814 3780 23818 3836
rect 23754 3776 23818 3780
rect 31219 3836 31283 3840
rect 31219 3780 31223 3836
rect 31223 3780 31279 3836
rect 31279 3780 31283 3836
rect 31219 3776 31283 3780
rect 31299 3836 31363 3840
rect 31299 3780 31303 3836
rect 31303 3780 31359 3836
rect 31359 3780 31363 3836
rect 31299 3776 31363 3780
rect 31379 3836 31443 3840
rect 31379 3780 31383 3836
rect 31383 3780 31439 3836
rect 31439 3780 31443 3836
rect 31379 3776 31443 3780
rect 31459 3836 31523 3840
rect 31459 3780 31463 3836
rect 31463 3780 31519 3836
rect 31519 3780 31523 3836
rect 31459 3776 31523 3780
rect 4252 3292 4316 3296
rect 4252 3236 4256 3292
rect 4256 3236 4312 3292
rect 4312 3236 4316 3292
rect 4252 3232 4316 3236
rect 4332 3292 4396 3296
rect 4332 3236 4336 3292
rect 4336 3236 4392 3292
rect 4392 3236 4396 3292
rect 4332 3232 4396 3236
rect 4412 3292 4476 3296
rect 4412 3236 4416 3292
rect 4416 3236 4472 3292
rect 4472 3236 4476 3292
rect 4412 3232 4476 3236
rect 4492 3292 4556 3296
rect 4492 3236 4496 3292
rect 4496 3236 4552 3292
rect 4552 3236 4556 3292
rect 4492 3232 4556 3236
rect 11957 3292 12021 3296
rect 11957 3236 11961 3292
rect 11961 3236 12017 3292
rect 12017 3236 12021 3292
rect 11957 3232 12021 3236
rect 12037 3292 12101 3296
rect 12037 3236 12041 3292
rect 12041 3236 12097 3292
rect 12097 3236 12101 3292
rect 12037 3232 12101 3236
rect 12117 3292 12181 3296
rect 12117 3236 12121 3292
rect 12121 3236 12177 3292
rect 12177 3236 12181 3292
rect 12117 3232 12181 3236
rect 12197 3292 12261 3296
rect 12197 3236 12201 3292
rect 12201 3236 12257 3292
rect 12257 3236 12261 3292
rect 12197 3232 12261 3236
rect 19662 3292 19726 3296
rect 19662 3236 19666 3292
rect 19666 3236 19722 3292
rect 19722 3236 19726 3292
rect 19662 3232 19726 3236
rect 19742 3292 19806 3296
rect 19742 3236 19746 3292
rect 19746 3236 19802 3292
rect 19802 3236 19806 3292
rect 19742 3232 19806 3236
rect 19822 3292 19886 3296
rect 19822 3236 19826 3292
rect 19826 3236 19882 3292
rect 19882 3236 19886 3292
rect 19822 3232 19886 3236
rect 19902 3292 19966 3296
rect 19902 3236 19906 3292
rect 19906 3236 19962 3292
rect 19962 3236 19966 3292
rect 19902 3232 19966 3236
rect 27367 3292 27431 3296
rect 27367 3236 27371 3292
rect 27371 3236 27427 3292
rect 27427 3236 27431 3292
rect 27367 3232 27431 3236
rect 27447 3292 27511 3296
rect 27447 3236 27451 3292
rect 27451 3236 27507 3292
rect 27507 3236 27511 3292
rect 27447 3232 27511 3236
rect 27527 3292 27591 3296
rect 27527 3236 27531 3292
rect 27531 3236 27587 3292
rect 27587 3236 27591 3292
rect 27527 3232 27591 3236
rect 27607 3292 27671 3296
rect 27607 3236 27611 3292
rect 27611 3236 27667 3292
rect 27667 3236 27671 3292
rect 27607 3232 27671 3236
rect 8104 2748 8168 2752
rect 8104 2692 8108 2748
rect 8108 2692 8164 2748
rect 8164 2692 8168 2748
rect 8104 2688 8168 2692
rect 8184 2748 8248 2752
rect 8184 2692 8188 2748
rect 8188 2692 8244 2748
rect 8244 2692 8248 2748
rect 8184 2688 8248 2692
rect 8264 2748 8328 2752
rect 8264 2692 8268 2748
rect 8268 2692 8324 2748
rect 8324 2692 8328 2748
rect 8264 2688 8328 2692
rect 8344 2748 8408 2752
rect 8344 2692 8348 2748
rect 8348 2692 8404 2748
rect 8404 2692 8408 2748
rect 8344 2688 8408 2692
rect 15809 2748 15873 2752
rect 15809 2692 15813 2748
rect 15813 2692 15869 2748
rect 15869 2692 15873 2748
rect 15809 2688 15873 2692
rect 15889 2748 15953 2752
rect 15889 2692 15893 2748
rect 15893 2692 15949 2748
rect 15949 2692 15953 2748
rect 15889 2688 15953 2692
rect 15969 2748 16033 2752
rect 15969 2692 15973 2748
rect 15973 2692 16029 2748
rect 16029 2692 16033 2748
rect 15969 2688 16033 2692
rect 16049 2748 16113 2752
rect 16049 2692 16053 2748
rect 16053 2692 16109 2748
rect 16109 2692 16113 2748
rect 16049 2688 16113 2692
rect 23514 2748 23578 2752
rect 23514 2692 23518 2748
rect 23518 2692 23574 2748
rect 23574 2692 23578 2748
rect 23514 2688 23578 2692
rect 23594 2748 23658 2752
rect 23594 2692 23598 2748
rect 23598 2692 23654 2748
rect 23654 2692 23658 2748
rect 23594 2688 23658 2692
rect 23674 2748 23738 2752
rect 23674 2692 23678 2748
rect 23678 2692 23734 2748
rect 23734 2692 23738 2748
rect 23674 2688 23738 2692
rect 23754 2748 23818 2752
rect 23754 2692 23758 2748
rect 23758 2692 23814 2748
rect 23814 2692 23818 2748
rect 23754 2688 23818 2692
rect 31219 2748 31283 2752
rect 31219 2692 31223 2748
rect 31223 2692 31279 2748
rect 31279 2692 31283 2748
rect 31219 2688 31283 2692
rect 31299 2748 31363 2752
rect 31299 2692 31303 2748
rect 31303 2692 31359 2748
rect 31359 2692 31363 2748
rect 31299 2688 31363 2692
rect 31379 2748 31443 2752
rect 31379 2692 31383 2748
rect 31383 2692 31439 2748
rect 31439 2692 31443 2748
rect 31379 2688 31443 2692
rect 31459 2748 31523 2752
rect 31459 2692 31463 2748
rect 31463 2692 31519 2748
rect 31519 2692 31523 2748
rect 31459 2688 31523 2692
rect 4252 2204 4316 2208
rect 4252 2148 4256 2204
rect 4256 2148 4312 2204
rect 4312 2148 4316 2204
rect 4252 2144 4316 2148
rect 4332 2204 4396 2208
rect 4332 2148 4336 2204
rect 4336 2148 4392 2204
rect 4392 2148 4396 2204
rect 4332 2144 4396 2148
rect 4412 2204 4476 2208
rect 4412 2148 4416 2204
rect 4416 2148 4472 2204
rect 4472 2148 4476 2204
rect 4412 2144 4476 2148
rect 4492 2204 4556 2208
rect 4492 2148 4496 2204
rect 4496 2148 4552 2204
rect 4552 2148 4556 2204
rect 4492 2144 4556 2148
rect 11957 2204 12021 2208
rect 11957 2148 11961 2204
rect 11961 2148 12017 2204
rect 12017 2148 12021 2204
rect 11957 2144 12021 2148
rect 12037 2204 12101 2208
rect 12037 2148 12041 2204
rect 12041 2148 12097 2204
rect 12097 2148 12101 2204
rect 12037 2144 12101 2148
rect 12117 2204 12181 2208
rect 12117 2148 12121 2204
rect 12121 2148 12177 2204
rect 12177 2148 12181 2204
rect 12117 2144 12181 2148
rect 12197 2204 12261 2208
rect 12197 2148 12201 2204
rect 12201 2148 12257 2204
rect 12257 2148 12261 2204
rect 12197 2144 12261 2148
rect 19662 2204 19726 2208
rect 19662 2148 19666 2204
rect 19666 2148 19722 2204
rect 19722 2148 19726 2204
rect 19662 2144 19726 2148
rect 19742 2204 19806 2208
rect 19742 2148 19746 2204
rect 19746 2148 19802 2204
rect 19802 2148 19806 2204
rect 19742 2144 19806 2148
rect 19822 2204 19886 2208
rect 19822 2148 19826 2204
rect 19826 2148 19882 2204
rect 19882 2148 19886 2204
rect 19822 2144 19886 2148
rect 19902 2204 19966 2208
rect 19902 2148 19906 2204
rect 19906 2148 19962 2204
rect 19962 2148 19966 2204
rect 19902 2144 19966 2148
rect 27367 2204 27431 2208
rect 27367 2148 27371 2204
rect 27371 2148 27427 2204
rect 27427 2148 27431 2204
rect 27367 2144 27431 2148
rect 27447 2204 27511 2208
rect 27447 2148 27451 2204
rect 27451 2148 27507 2204
rect 27507 2148 27511 2204
rect 27447 2144 27511 2148
rect 27527 2204 27591 2208
rect 27527 2148 27531 2204
rect 27531 2148 27587 2204
rect 27587 2148 27591 2204
rect 27527 2144 27591 2148
rect 27607 2204 27671 2208
rect 27607 2148 27611 2204
rect 27611 2148 27667 2204
rect 27667 2148 27671 2204
rect 27607 2144 27671 2148
rect 8104 1660 8168 1664
rect 8104 1604 8108 1660
rect 8108 1604 8164 1660
rect 8164 1604 8168 1660
rect 8104 1600 8168 1604
rect 8184 1660 8248 1664
rect 8184 1604 8188 1660
rect 8188 1604 8244 1660
rect 8244 1604 8248 1660
rect 8184 1600 8248 1604
rect 8264 1660 8328 1664
rect 8264 1604 8268 1660
rect 8268 1604 8324 1660
rect 8324 1604 8328 1660
rect 8264 1600 8328 1604
rect 8344 1660 8408 1664
rect 8344 1604 8348 1660
rect 8348 1604 8404 1660
rect 8404 1604 8408 1660
rect 8344 1600 8408 1604
rect 15809 1660 15873 1664
rect 15809 1604 15813 1660
rect 15813 1604 15869 1660
rect 15869 1604 15873 1660
rect 15809 1600 15873 1604
rect 15889 1660 15953 1664
rect 15889 1604 15893 1660
rect 15893 1604 15949 1660
rect 15949 1604 15953 1660
rect 15889 1600 15953 1604
rect 15969 1660 16033 1664
rect 15969 1604 15973 1660
rect 15973 1604 16029 1660
rect 16029 1604 16033 1660
rect 15969 1600 16033 1604
rect 16049 1660 16113 1664
rect 16049 1604 16053 1660
rect 16053 1604 16109 1660
rect 16109 1604 16113 1660
rect 16049 1600 16113 1604
rect 23514 1660 23578 1664
rect 23514 1604 23518 1660
rect 23518 1604 23574 1660
rect 23574 1604 23578 1660
rect 23514 1600 23578 1604
rect 23594 1660 23658 1664
rect 23594 1604 23598 1660
rect 23598 1604 23654 1660
rect 23654 1604 23658 1660
rect 23594 1600 23658 1604
rect 23674 1660 23738 1664
rect 23674 1604 23678 1660
rect 23678 1604 23734 1660
rect 23734 1604 23738 1660
rect 23674 1600 23738 1604
rect 23754 1660 23818 1664
rect 23754 1604 23758 1660
rect 23758 1604 23814 1660
rect 23814 1604 23818 1660
rect 23754 1600 23818 1604
rect 31219 1660 31283 1664
rect 31219 1604 31223 1660
rect 31223 1604 31279 1660
rect 31279 1604 31283 1660
rect 31219 1600 31283 1604
rect 31299 1660 31363 1664
rect 31299 1604 31303 1660
rect 31303 1604 31359 1660
rect 31359 1604 31363 1660
rect 31299 1600 31363 1604
rect 31379 1660 31443 1664
rect 31379 1604 31383 1660
rect 31383 1604 31439 1660
rect 31439 1604 31443 1660
rect 31379 1600 31443 1604
rect 31459 1660 31523 1664
rect 31459 1604 31463 1660
rect 31463 1604 31519 1660
rect 31519 1604 31523 1660
rect 31459 1600 31523 1604
rect 4252 1116 4316 1120
rect 4252 1060 4256 1116
rect 4256 1060 4312 1116
rect 4312 1060 4316 1116
rect 4252 1056 4316 1060
rect 4332 1116 4396 1120
rect 4332 1060 4336 1116
rect 4336 1060 4392 1116
rect 4392 1060 4396 1116
rect 4332 1056 4396 1060
rect 4412 1116 4476 1120
rect 4412 1060 4416 1116
rect 4416 1060 4472 1116
rect 4472 1060 4476 1116
rect 4412 1056 4476 1060
rect 4492 1116 4556 1120
rect 4492 1060 4496 1116
rect 4496 1060 4552 1116
rect 4552 1060 4556 1116
rect 4492 1056 4556 1060
rect 11957 1116 12021 1120
rect 11957 1060 11961 1116
rect 11961 1060 12017 1116
rect 12017 1060 12021 1116
rect 11957 1056 12021 1060
rect 12037 1116 12101 1120
rect 12037 1060 12041 1116
rect 12041 1060 12097 1116
rect 12097 1060 12101 1116
rect 12037 1056 12101 1060
rect 12117 1116 12181 1120
rect 12117 1060 12121 1116
rect 12121 1060 12177 1116
rect 12177 1060 12181 1116
rect 12117 1056 12181 1060
rect 12197 1116 12261 1120
rect 12197 1060 12201 1116
rect 12201 1060 12257 1116
rect 12257 1060 12261 1116
rect 12197 1056 12261 1060
rect 19662 1116 19726 1120
rect 19662 1060 19666 1116
rect 19666 1060 19722 1116
rect 19722 1060 19726 1116
rect 19662 1056 19726 1060
rect 19742 1116 19806 1120
rect 19742 1060 19746 1116
rect 19746 1060 19802 1116
rect 19802 1060 19806 1116
rect 19742 1056 19806 1060
rect 19822 1116 19886 1120
rect 19822 1060 19826 1116
rect 19826 1060 19882 1116
rect 19882 1060 19886 1116
rect 19822 1056 19886 1060
rect 19902 1116 19966 1120
rect 19902 1060 19906 1116
rect 19906 1060 19962 1116
rect 19962 1060 19966 1116
rect 19902 1056 19966 1060
rect 27367 1116 27431 1120
rect 27367 1060 27371 1116
rect 27371 1060 27427 1116
rect 27427 1060 27431 1116
rect 27367 1056 27431 1060
rect 27447 1116 27511 1120
rect 27447 1060 27451 1116
rect 27451 1060 27507 1116
rect 27507 1060 27511 1116
rect 27447 1056 27511 1060
rect 27527 1116 27591 1120
rect 27527 1060 27531 1116
rect 27531 1060 27587 1116
rect 27587 1060 27591 1116
rect 27527 1056 27591 1060
rect 27607 1116 27671 1120
rect 27607 1060 27611 1116
rect 27611 1060 27667 1116
rect 27667 1060 27671 1116
rect 27607 1056 27671 1060
rect 8104 572 8168 576
rect 8104 516 8108 572
rect 8108 516 8164 572
rect 8164 516 8168 572
rect 8104 512 8168 516
rect 8184 572 8248 576
rect 8184 516 8188 572
rect 8188 516 8244 572
rect 8244 516 8248 572
rect 8184 512 8248 516
rect 8264 572 8328 576
rect 8264 516 8268 572
rect 8268 516 8324 572
rect 8324 516 8328 572
rect 8264 512 8328 516
rect 8344 572 8408 576
rect 8344 516 8348 572
rect 8348 516 8404 572
rect 8404 516 8408 572
rect 8344 512 8408 516
rect 15809 572 15873 576
rect 15809 516 15813 572
rect 15813 516 15869 572
rect 15869 516 15873 572
rect 15809 512 15873 516
rect 15889 572 15953 576
rect 15889 516 15893 572
rect 15893 516 15949 572
rect 15949 516 15953 572
rect 15889 512 15953 516
rect 15969 572 16033 576
rect 15969 516 15973 572
rect 15973 516 16029 572
rect 16029 516 16033 572
rect 15969 512 16033 516
rect 16049 572 16113 576
rect 16049 516 16053 572
rect 16053 516 16109 572
rect 16109 516 16113 572
rect 16049 512 16113 516
rect 23514 572 23578 576
rect 23514 516 23518 572
rect 23518 516 23574 572
rect 23574 516 23578 572
rect 23514 512 23578 516
rect 23594 572 23658 576
rect 23594 516 23598 572
rect 23598 516 23654 572
rect 23654 516 23658 572
rect 23594 512 23658 516
rect 23674 572 23738 576
rect 23674 516 23678 572
rect 23678 516 23734 572
rect 23734 516 23738 572
rect 23674 512 23738 516
rect 23754 572 23818 576
rect 23754 516 23758 572
rect 23758 516 23814 572
rect 23814 516 23818 572
rect 23754 512 23818 516
rect 31219 572 31283 576
rect 31219 516 31223 572
rect 31223 516 31279 572
rect 31279 516 31283 572
rect 31219 512 31283 516
rect 31299 572 31363 576
rect 31299 516 31303 572
rect 31303 516 31359 572
rect 31359 516 31363 572
rect 31299 512 31363 516
rect 31379 572 31443 576
rect 31379 516 31383 572
rect 31383 516 31439 572
rect 31439 516 31443 572
rect 31379 512 31443 516
rect 31459 572 31523 576
rect 31459 516 31463 572
rect 31463 516 31519 572
rect 31519 516 31523 572
rect 31459 512 31523 516
<< metal4 >>
rect 4244 18528 4564 19088
rect 4244 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4564 18528
rect 4244 17440 4564 18464
rect 4244 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4564 17440
rect 4244 16352 4564 17376
rect 4244 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4564 16352
rect 4244 15264 4564 16288
rect 4244 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4564 15264
rect 4244 14176 4564 15200
rect 4244 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4564 14176
rect 4244 13088 4564 14112
rect 4244 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4564 13088
rect 4244 12000 4564 13024
rect 4244 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4564 12000
rect 4244 10912 4564 11936
rect 4244 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4564 10912
rect 4244 9824 4564 10848
rect 4244 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4564 9824
rect 4244 8736 4564 9760
rect 4244 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4564 8736
rect 4244 7648 4564 8672
rect 4244 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4564 7648
rect 4244 6560 4564 7584
rect 4244 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4564 6560
rect 4244 5472 4564 6496
rect 4244 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4564 5472
rect 4244 4384 4564 5408
rect 4244 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4564 4384
rect 4244 3296 4564 4320
rect 4244 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4564 3296
rect 4244 2208 4564 3232
rect 4244 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4564 2208
rect 4244 1120 4564 2144
rect 4244 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4564 1120
rect 4244 496 4564 1056
rect 8096 19072 8416 19088
rect 8096 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8416 19072
rect 8096 17984 8416 19008
rect 8096 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8416 17984
rect 8096 16896 8416 17920
rect 8096 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8416 16896
rect 8096 15808 8416 16832
rect 8096 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8416 15808
rect 8096 14720 8416 15744
rect 8096 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8416 14720
rect 8096 13632 8416 14656
rect 8096 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8416 13632
rect 8096 12544 8416 13568
rect 8096 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8416 12544
rect 8096 11456 8416 12480
rect 8096 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8416 11456
rect 8096 10368 8416 11392
rect 8096 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8416 10368
rect 8096 9280 8416 10304
rect 8096 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8416 9280
rect 8096 8192 8416 9216
rect 8096 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8416 8192
rect 8096 7104 8416 8128
rect 8096 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8416 7104
rect 8096 6016 8416 7040
rect 8096 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8416 6016
rect 8096 4928 8416 5952
rect 8096 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8416 4928
rect 8096 3840 8416 4864
rect 8096 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8416 3840
rect 8096 2752 8416 3776
rect 8096 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8416 2752
rect 8096 1664 8416 2688
rect 8096 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8416 1664
rect 8096 576 8416 1600
rect 8096 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8416 576
rect 8096 496 8416 512
rect 11949 18528 12269 19088
rect 11949 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12269 18528
rect 11949 17440 12269 18464
rect 11949 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12269 17440
rect 11949 16352 12269 17376
rect 11949 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12269 16352
rect 11949 15264 12269 16288
rect 11949 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12269 15264
rect 11949 14176 12269 15200
rect 11949 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12269 14176
rect 11949 13088 12269 14112
rect 11949 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12269 13088
rect 11949 12000 12269 13024
rect 11949 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12269 12000
rect 11949 10912 12269 11936
rect 11949 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12269 10912
rect 11949 9824 12269 10848
rect 11949 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12269 9824
rect 11949 8736 12269 9760
rect 11949 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12269 8736
rect 11949 7648 12269 8672
rect 11949 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12269 7648
rect 11949 6560 12269 7584
rect 11949 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12269 6560
rect 11949 5472 12269 6496
rect 11949 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12269 5472
rect 11949 4384 12269 5408
rect 11949 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12269 4384
rect 11949 3296 12269 4320
rect 11949 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12269 3296
rect 11949 2208 12269 3232
rect 11949 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12269 2208
rect 11949 1120 12269 2144
rect 11949 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12269 1120
rect 11949 496 12269 1056
rect 15801 19072 16121 19088
rect 15801 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16121 19072
rect 15801 17984 16121 19008
rect 15801 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16121 17984
rect 15801 16896 16121 17920
rect 15801 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16121 16896
rect 15801 15808 16121 16832
rect 15801 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16121 15808
rect 15801 14720 16121 15744
rect 15801 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16121 14720
rect 15801 13632 16121 14656
rect 15801 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16121 13632
rect 15801 12544 16121 13568
rect 15801 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16121 12544
rect 15801 11456 16121 12480
rect 15801 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16121 11456
rect 15801 10368 16121 11392
rect 15801 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16121 10368
rect 15801 9280 16121 10304
rect 15801 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16121 9280
rect 15801 8192 16121 9216
rect 15801 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16121 8192
rect 15801 7104 16121 8128
rect 15801 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16121 7104
rect 15801 6016 16121 7040
rect 15801 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16121 6016
rect 15801 4928 16121 5952
rect 15801 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16121 4928
rect 15801 3840 16121 4864
rect 15801 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16121 3840
rect 15801 2752 16121 3776
rect 15801 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16121 2752
rect 15801 1664 16121 2688
rect 15801 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16121 1664
rect 15801 576 16121 1600
rect 15801 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16121 576
rect 15801 496 16121 512
rect 19654 18528 19974 19088
rect 19654 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19974 18528
rect 19654 17440 19974 18464
rect 19654 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19974 17440
rect 19654 16352 19974 17376
rect 19654 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19974 16352
rect 19654 15264 19974 16288
rect 19654 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19974 15264
rect 19654 14176 19974 15200
rect 19654 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19974 14176
rect 19654 13088 19974 14112
rect 19654 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19974 13088
rect 19654 12000 19974 13024
rect 19654 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19974 12000
rect 19654 10912 19974 11936
rect 19654 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19974 10912
rect 19654 9824 19974 10848
rect 19654 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19974 9824
rect 19654 8736 19974 9760
rect 19654 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19974 8736
rect 19654 7648 19974 8672
rect 19654 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19974 7648
rect 19654 6560 19974 7584
rect 19654 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19974 6560
rect 19654 5472 19974 6496
rect 19654 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19974 5472
rect 19654 4384 19974 5408
rect 19654 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19974 4384
rect 19654 3296 19974 4320
rect 19654 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19974 3296
rect 19654 2208 19974 3232
rect 19654 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19974 2208
rect 19654 1120 19974 2144
rect 19654 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19974 1120
rect 19654 496 19974 1056
rect 23506 19072 23826 19088
rect 23506 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23826 19072
rect 23506 17984 23826 19008
rect 23506 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23826 17984
rect 23506 16896 23826 17920
rect 23506 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23826 16896
rect 23506 15808 23826 16832
rect 23506 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23826 15808
rect 23506 14720 23826 15744
rect 23506 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23826 14720
rect 23506 13632 23826 14656
rect 23506 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23826 13632
rect 23506 12544 23826 13568
rect 23506 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23826 12544
rect 23506 11456 23826 12480
rect 23506 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23826 11456
rect 23506 10368 23826 11392
rect 23506 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23826 10368
rect 23506 9280 23826 10304
rect 23506 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23826 9280
rect 23506 8192 23826 9216
rect 23506 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23826 8192
rect 23506 7104 23826 8128
rect 23506 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23826 7104
rect 23506 6016 23826 7040
rect 23506 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23826 6016
rect 23506 4928 23826 5952
rect 23506 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23826 4928
rect 23506 3840 23826 4864
rect 23506 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23826 3840
rect 23506 2752 23826 3776
rect 23506 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23826 2752
rect 23506 1664 23826 2688
rect 23506 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23826 1664
rect 23506 576 23826 1600
rect 23506 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23826 576
rect 23506 496 23826 512
rect 27359 18528 27679 19088
rect 27359 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27679 18528
rect 27359 17440 27679 18464
rect 27359 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27679 17440
rect 27359 16352 27679 17376
rect 27359 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27679 16352
rect 27359 15264 27679 16288
rect 27359 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27679 15264
rect 27359 14176 27679 15200
rect 27359 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27679 14176
rect 27359 13088 27679 14112
rect 27359 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27679 13088
rect 27359 12000 27679 13024
rect 27359 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27679 12000
rect 27359 10912 27679 11936
rect 27359 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27679 10912
rect 27359 9824 27679 10848
rect 27359 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27679 9824
rect 27359 8736 27679 9760
rect 27359 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27679 8736
rect 27359 7648 27679 8672
rect 27359 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27679 7648
rect 27359 6560 27679 7584
rect 27359 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27679 6560
rect 27359 5472 27679 6496
rect 27359 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27679 5472
rect 27359 4384 27679 5408
rect 27359 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27679 4384
rect 27359 3296 27679 4320
rect 27359 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27679 3296
rect 27359 2208 27679 3232
rect 27359 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27679 2208
rect 27359 1120 27679 2144
rect 27359 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27679 1120
rect 27359 496 27679 1056
rect 31211 19072 31531 19088
rect 31211 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31531 19072
rect 31211 17984 31531 19008
rect 31211 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31531 17984
rect 31211 16896 31531 17920
rect 31211 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31531 16896
rect 31211 15808 31531 16832
rect 31211 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31531 15808
rect 31211 14720 31531 15744
rect 31211 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31531 14720
rect 31211 13632 31531 14656
rect 31211 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31531 13632
rect 31211 12544 31531 13568
rect 31211 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31531 12544
rect 31211 11456 31531 12480
rect 31211 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31531 11456
rect 31211 10368 31531 11392
rect 31211 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31531 10368
rect 31211 9280 31531 10304
rect 31211 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31531 9280
rect 31211 8192 31531 9216
rect 31211 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31531 8192
rect 31211 7104 31531 8128
rect 31211 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31531 7104
rect 31211 6016 31531 7040
rect 31211 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31531 6016
rect 31211 4928 31531 5952
rect 31211 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31531 4928
rect 31211 3840 31531 4864
rect 31211 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31531 3840
rect 31211 2752 31531 3776
rect 31211 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31531 2752
rect 31211 1664 31531 2688
rect 31211 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31531 1664
rect 31211 576 31531 1600
rect 31211 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31531 576
rect 31211 496 31531 512
use sky130_fd_sc_hd__dfxtp_2  _00_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13064 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _01_
timestamp 1701704242
transform 1 0 14444 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _02_
timestamp 1701704242
transform -1 0 12880 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _03_
timestamp 1701704242
transform 1 0 14628 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _04_
timestamp 1701704242
transform 1 0 16100 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _05_
timestamp 1701704242
transform -1 0 16100 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _06_
timestamp 1701704242
transform 1 0 13616 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _07_
timestamp 1701704242
transform 1 0 11868 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _08_
timestamp 1701704242
transform 1 0 11040 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _09_
timestamp 1701704242
transform -1 0 10488 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _10_
timestamp 1701704242
transform -1 0 9292 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _11_
timestamp 1701704242
transform -1 0 12512 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _12_
timestamp 1701704242
transform -1 0 8096 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _13_
timestamp 1701704242
transform -1 0 10764 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _14_
timestamp 1701704242
transform -1 0 8188 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _15_
timestamp 1701704242
transform -1 0 10856 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _16_
timestamp 1701704242
transform -1 0 11224 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _17_
timestamp 1701704242
transform -1 0 8556 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _18_
timestamp 1701704242
transform -1 0 9568 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _19_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10488 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _20_
timestamp 1701704242
transform -1 0 12788 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _21_
timestamp 1701704242
transform 1 0 12788 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _22_
timestamp 1701704242
transform 1 0 13984 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _23_
timestamp 1701704242
transform 1 0 12144 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _24_
timestamp 1701704242
transform -1 0 10488 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _25_
timestamp 1701704242
transform -1 0 11500 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _26_
timestamp 1701704242
transform 1 0 13708 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _27_
timestamp 1701704242
transform 1 0 11500 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _28_
timestamp 1701704242
transform 1 0 12880 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _29_
timestamp 1701704242
transform 1 0 14444 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _30_
timestamp 1701704242
transform 1 0 16192 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _31_
timestamp 1701704242
transform 1 0 17572 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _32_
timestamp 1701704242
transform 1 0 16560 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _33_
timestamp 1701704242
transform 1 0 18676 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _34_
timestamp 1701704242
transform 1 0 19596 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _35_
timestamp 1701704242
transform 1 0 22172 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _36_
timestamp 1701704242
transform 1 0 20608 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _37_
timestamp 1701704242
transform 1 0 23368 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _38_
timestamp 1701704242
transform 1 0 17020 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _39_
timestamp 1701704242
transform 1 0 19044 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _40_
timestamp 1701704242
transform 1 0 22172 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _41_
timestamp 1701704242
transform 1 0 22908 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _42_
timestamp 1701704242
transform 1 0 22908 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _43_
timestamp 1701704242
transform 1 0 21988 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _44_
timestamp 1701704242
transform 1 0 17020 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _45_
timestamp 1701704242
transform -1 0 15364 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _46_
timestamp 1701704242
transform 1 0 14536 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _47_
timestamp 1701704242
transform 1 0 16100 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _48_
timestamp 1701704242
transform 1 0 18768 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _49_
timestamp 1701704242
transform 1 0 17020 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _50_
timestamp 1701704242
transform 1 0 20332 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _51_
timestamp 1701704242
transform 1 0 21252 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _52_
timestamp 1701704242
transform 1 0 21988 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _53_
timestamp 1701704242
transform 1 0 21896 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _54_
timestamp 1701704242
transform 1 0 21436 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _55_
timestamp 1701704242
transform 1 0 17756 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _56_
timestamp 1701704242
transform 1 0 19780 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _57_
timestamp 1701704242
transform 1 0 19320 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _58_
timestamp 1701704242
transform 1 0 16192 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _59_
timestamp 1701704242
transform 1 0 18308 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _60_
timestamp 1701704242
transform 1 0 17020 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _61_
timestamp 1701704242
transform 1 0 16100 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _62_
timestamp 1701704242
transform 1 0 14352 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _63_
timestamp 1701704242
transform -1 0 14260 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _64_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16376 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_i_stop pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16100 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_i_stop
timestamp 1701704242
transform -1 0 10856 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_i_stop
timestamp 1701704242
transform -1 0 16008 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_i_stop
timestamp 1701704242
transform 1 0 9844 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_i_stop
timestamp 1701704242
transform -1 0 16560 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_i_stop
timestamp 1701704242
transform -1 0 18584 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_i_stop
timestamp 1701704242
transform 1 0 21344 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_i_stop
timestamp 1701704242
transform 1 0 16928 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_i_stop
timestamp 1701704242
transform 1 0 21528 0 -1 12512
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1701704242
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1701704242
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1701704242
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1701704242
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1701704242
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1701704242
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1701704242
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1701704242
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1701704242
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1701704242
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1701704242
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1701704242
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1701704242
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1701704242
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1701704242
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1701704242
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1701704242
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1701704242
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1701704242
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_237
timestamp 1701704242
transform 1 0 22356 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_250 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 23552 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1701704242
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1701704242
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1701704242
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1701704242
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1701704242
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1701704242
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1701704242
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_321 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 30084 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_329
timestamp 1701704242
transform 1 0 30820 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1701704242
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1701704242
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1701704242
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1701704242
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1701704242
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1701704242
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1701704242
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1701704242
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1701704242
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1701704242
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1701704242
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1701704242
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1701704242
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1701704242
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1701704242
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1701704242
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1701704242
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1701704242
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1701704242
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1701704242
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1701704242
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1701704242
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1701704242
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1701704242
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1701704242
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1701704242
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1701704242
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1701704242
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_329
timestamp 1701704242
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1701704242
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1701704242
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1701704242
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1701704242
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1701704242
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1701704242
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1701704242
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1701704242
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1701704242
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1701704242
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1701704242
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1701704242
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1701704242
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1701704242
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1701704242
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1701704242
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1701704242
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1701704242
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1701704242
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1701704242
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1701704242
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1701704242
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1701704242
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1701704242
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1701704242
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1701704242
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1701704242
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1701704242
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1701704242
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1701704242
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1701704242
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1701704242
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1701704242
transform 1 0 30084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_329
timestamp 1701704242
transform 1 0 30820 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1701704242
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1701704242
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1701704242
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1701704242
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1701704242
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1701704242
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1701704242
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1701704242
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1701704242
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1701704242
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1701704242
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1701704242
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1701704242
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1701704242
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1701704242
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1701704242
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1701704242
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1701704242
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1701704242
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1701704242
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1701704242
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1701704242
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1701704242
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1701704242
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1701704242
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1701704242
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1701704242
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1701704242
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1701704242
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1701704242
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1701704242
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_329
timestamp 1701704242
transform 1 0 30820 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1701704242
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1701704242
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1701704242
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1701704242
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1701704242
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1701704242
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1701704242
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1701704242
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1701704242
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1701704242
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1701704242
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1701704242
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1701704242
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1701704242
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1701704242
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1701704242
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1701704242
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1701704242
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1701704242
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1701704242
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1701704242
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1701704242
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1701704242
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1701704242
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1701704242
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1701704242
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1701704242
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1701704242
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1701704242
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_321
timestamp 1701704242
transform 1 0 30084 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_329
timestamp 1701704242
transform 1 0 30820 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1701704242
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1701704242
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1701704242
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1701704242
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1701704242
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1701704242
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1701704242
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1701704242
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1701704242
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1701704242
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1701704242
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1701704242
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1701704242
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1701704242
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1701704242
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1701704242
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1701704242
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1701704242
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1701704242
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1701704242
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1701704242
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1701704242
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1701704242
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1701704242
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1701704242
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1701704242
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1701704242
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1701704242
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1701704242
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1701704242
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1701704242
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_329
timestamp 1701704242
transform 1 0 30820 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1701704242
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1701704242
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1701704242
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1701704242
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1701704242
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1701704242
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1701704242
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1701704242
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1701704242
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1701704242
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1701704242
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1701704242
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1701704242
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1701704242
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1701704242
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1701704242
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1701704242
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1701704242
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1701704242
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1701704242
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1701704242
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1701704242
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1701704242
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1701704242
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1701704242
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1701704242
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1701704242
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1701704242
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1701704242
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1701704242
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1701704242
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_321
timestamp 1701704242
transform 1 0 30084 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_329
timestamp 1701704242
transform 1 0 30820 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1701704242
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1701704242
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1701704242
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1701704242
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1701704242
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1701704242
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1701704242
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1701704242
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1701704242
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1701704242
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1701704242
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1701704242
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1701704242
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1701704242
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1701704242
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1701704242
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1701704242
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_169
timestamp 1701704242
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_174
timestamp 1701704242
transform 1 0 16560 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_186
timestamp 1701704242
transform 1 0 17664 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_198
timestamp 1701704242
transform 1 0 18768 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_210
timestamp 1701704242
transform 1 0 19872 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1701704242
transform 1 0 20976 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1701704242
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1701704242
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1701704242
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1701704242
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1701704242
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1701704242
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1701704242
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1701704242
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1701704242
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1701704242
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_329
timestamp 1701704242
transform 1 0 30820 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1701704242
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1701704242
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1701704242
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1701704242
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1701704242
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1701704242
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1701704242
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1701704242
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1701704242
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1701704242
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1701704242
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1701704242
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1701704242
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1701704242
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_153
timestamp 1701704242
transform 1 0 14628 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_161
timestamp 1701704242
transform 1 0 15364 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_178
timestamp 1701704242
transform 1 0 16928 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1701704242
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1701704242
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1701704242
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1701704242
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1701704242
transform 1 0 23092 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1701704242
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1701704242
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1701704242
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1701704242
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1701704242
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1701704242
transform 1 0 28244 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1701704242
transform 1 0 28796 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1701704242
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_321
timestamp 1701704242
transform 1 0 30084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_329
timestamp 1701704242
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1701704242
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1701704242
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1701704242
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1701704242
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1701704242
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1701704242
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1701704242
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1701704242
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1701704242
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1701704242
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1701704242
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1701704242
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1701704242
transform 1 0 10948 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_131
timestamp 1701704242
transform 1 0 12604 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_143
timestamp 1701704242
transform 1 0 13708 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1701704242
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1701704242
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_175
timestamp 1701704242
transform 1 0 16652 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_185
timestamp 1701704242
transform 1 0 17572 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_204
timestamp 1701704242
transform 1 0 19320 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_216
timestamp 1701704242
transform 1 0 20424 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1701704242
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1701704242
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1701704242
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1701704242
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1701704242
transform 1 0 25668 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1701704242
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1701704242
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1701704242
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1701704242
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1701704242
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_329
timestamp 1701704242
transform 1 0 30820 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1701704242
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1701704242
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1701704242
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1701704242
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1701704242
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1701704242
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1701704242
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1701704242
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_85
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_111
timestamp 1701704242
transform 1 0 10764 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_115
timestamp 1701704242
transform 1 0 11132 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_141
timestamp 1701704242
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_149
timestamp 1701704242
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1701704242
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_197
timestamp 1701704242
transform 1 0 18676 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_232
timestamp 1701704242
transform 1 0 21896 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_244
timestamp 1701704242
transform 1 0 23000 0 1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1701704242
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1701704242
transform 1 0 24932 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1701704242
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1701704242
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1701704242
transform 1 0 28244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1701704242
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1701704242
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_321
timestamp 1701704242
transform 1 0 30084 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_329
timestamp 1701704242
transform 1 0 30820 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1701704242
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1701704242
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1701704242
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1701704242
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1701704242
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_69
timestamp 1701704242
transform 1 0 6900 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_77
timestamp 1701704242
transform 1 0 7636 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_98
timestamp 1701704242
transform 1 0 9568 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_131
timestamp 1701704242
transform 1 0 12604 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_139
timestamp 1701704242
transform 1 0 13340 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_159
timestamp 1701704242
transform 1 0 15180 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1701704242
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1701704242
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_177
timestamp 1701704242
transform 1 0 16836 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1701704242
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_242
timestamp 1701704242
transform 1 0 22816 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_254
timestamp 1701704242
transform 1 0 23920 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_266
timestamp 1701704242
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 1701704242
transform 1 0 26128 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1701704242
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1701704242
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1701704242
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1701704242
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_329
timestamp 1701704242
transform 1 0 30820 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1701704242
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1701704242
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1701704242
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1701704242
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_65
timestamp 1701704242
transform 1 0 6532 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_73
timestamp 1701704242
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_88
timestamp 1701704242
transform 1 0 8648 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_95
timestamp 1701704242
transform 1 0 9292 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_108
timestamp 1701704242
transform 1 0 10488 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_120
timestamp 1701704242
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1701704242
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_169
timestamp 1701704242
transform 1 0 16100 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_175
timestamp 1701704242
transform 1 0 16652 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_197
timestamp 1701704242
transform 1 0 18676 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_203
timestamp 1701704242
transform 1 0 19228 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_231
timestamp 1701704242
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1701704242
transform 1 0 23552 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1701704242
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1701704242
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1701704242
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1701704242
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1701704242
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1701704242
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1701704242
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_321
timestamp 1701704242
transform 1 0 30084 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_329
timestamp 1701704242
transform 1 0 30820 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1701704242
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1701704242
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1701704242
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1701704242
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1701704242
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1701704242
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1701704242
transform 1 0 5796 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_82
timestamp 1701704242
transform 1 0 8096 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_130
timestamp 1701704242
transform 1 0 12512 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_186
timestamp 1701704242
transform 1 0 17664 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_204
timestamp 1701704242
transform 1 0 19320 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_208
timestamp 1701704242
transform 1 0 19688 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_231
timestamp 1701704242
transform 1 0 21804 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1701704242
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1701704242
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1701704242
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1701704242
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1701704242
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1701704242
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1701704242
transform 1 0 28612 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1701704242
transform 1 0 29716 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_329
timestamp 1701704242
transform 1 0 30820 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1701704242
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1701704242
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1701704242
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1701704242
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1701704242
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_77
timestamp 1701704242
transform 1 0 7636 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1701704242
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_93
timestamp 1701704242
transform 1 0 9108 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_111
timestamp 1701704242
transform 1 0 10764 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_134
timestamp 1701704242
transform 1 0 12880 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_170
timestamp 1701704242
transform 1 0 16192 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_182
timestamp 1701704242
transform 1 0 17296 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1701704242
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp 1701704242
transform 1 0 18676 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_249
timestamp 1701704242
transform 1 0 23460 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1701704242
transform 1 0 23828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1701704242
transform 1 0 24932 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1701704242
transform 1 0 26036 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1701704242
transform 1 0 27140 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1701704242
transform 1 0 28244 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1701704242
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1701704242
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_321
timestamp 1701704242
transform 1 0 30084 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_329
timestamp 1701704242
transform 1 0 30820 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1701704242
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1701704242
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1701704242
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1701704242
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1701704242
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1701704242
transform 1 0 5796 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_65
timestamp 1701704242
transform 1 0 6532 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1701704242
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_125
timestamp 1701704242
transform 1 0 12052 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_137
timestamp 1701704242
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_169
timestamp 1701704242
transform 1 0 16100 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_187
timestamp 1701704242
transform 1 0 17756 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1701704242
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_225
timestamp 1701704242
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_246
timestamp 1701704242
transform 1 0 23184 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_258
timestamp 1701704242
transform 1 0 24288 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_270
timestamp 1701704242
transform 1 0 25392 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 1701704242
transform 1 0 26128 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1701704242
transform 1 0 26404 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1701704242
transform 1 0 27508 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1701704242
transform 1 0 28612 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1701704242
transform 1 0 29716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_329
timestamp 1701704242
transform 1 0 30820 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1701704242
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1701704242
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1701704242
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1701704242
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1701704242
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_77
timestamp 1701704242
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_88
timestamp 1701704242
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_98
timestamp 1701704242
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_116
timestamp 1701704242
transform 1 0 11224 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1701704242
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_144
timestamp 1701704242
transform 1 0 13800 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_160
timestamp 1701704242
transform 1 0 15272 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_183
timestamp 1701704242
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1701704242
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_203
timestamp 1701704242
transform 1 0 19228 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1701704242
transform 1 0 20884 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1701704242
transform 1 0 23552 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1701704242
transform 1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1701704242
transform 1 0 24932 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1701704242
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1701704242
transform 1 0 27140 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1701704242
transform 1 0 28244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1701704242
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1701704242
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_321
timestamp 1701704242
transform 1 0 30084 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_329
timestamp 1701704242
transform 1 0 30820 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1701704242
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1701704242
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1701704242
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1701704242
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1701704242
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1701704242
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_69
timestamp 1701704242
transform 1 0 6900 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_87
timestamp 1701704242
transform 1 0 8556 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_94
timestamp 1701704242
transform 1 0 9200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_106
timestamp 1701704242
transform 1 0 10304 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_125
timestamp 1701704242
transform 1 0 12052 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_129
timestamp 1701704242
transform 1 0 12420 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_149
timestamp 1701704242
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_192
timestamp 1701704242
transform 1 0 18216 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_210
timestamp 1701704242
transform 1 0 19872 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_222
timestamp 1701704242
transform 1 0 20976 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_260
timestamp 1701704242
transform 1 0 24472 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_272
timestamp 1701704242
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1701704242
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1701704242
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1701704242
transform 1 0 28612 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1701704242
transform 1 0 29716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_329
timestamp 1701704242
transform 1 0 30820 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1701704242
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1701704242
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1701704242
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1701704242
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1701704242
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1701704242
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1701704242
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1701704242
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1701704242
transform 1 0 8372 0 1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_127
timestamp 1701704242
transform 1 0 12236 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1701704242
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_141
timestamp 1701704242
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_152
timestamp 1701704242
transform 1 0 14536 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_158
timestamp 1701704242
transform 1 0 15088 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_162
timestamp 1701704242
transform 1 0 15456 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_169
timestamp 1701704242
transform 1 0 16100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_177
timestamp 1701704242
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1701704242
transform 1 0 18676 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1701704242
transform 1 0 19780 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_221
timestamp 1701704242
transform 1 0 20884 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_244
timestamp 1701704242
transform 1 0 23000 0 1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1701704242
transform 1 0 23828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1701704242
transform 1 0 24932 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1701704242
transform 1 0 26036 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1701704242
transform 1 0 27140 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1701704242
transform 1 0 28244 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1701704242
transform 1 0 28796 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1701704242
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_321
timestamp 1701704242
transform 1 0 30084 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_329
timestamp 1701704242
transform 1 0 30820 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1701704242
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1701704242
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1701704242
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1701704242
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1701704242
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1701704242
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_98
timestamp 1701704242
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1701704242
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1701704242
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_186
timestamp 1701704242
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_198
timestamp 1701704242
transform 1 0 18768 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1701704242
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_260
timestamp 1701704242
transform 1 0 24472 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_272
timestamp 1701704242
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1701704242
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1701704242
transform 1 0 27508 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1701704242
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1701704242
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_329
timestamp 1701704242
transform 1 0 30820 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1701704242
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1701704242
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1701704242
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1701704242
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1701704242
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1701704242
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1701704242
transform 1 0 6532 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1701704242
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1701704242
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 1701704242
transform 1 0 8372 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_91
timestamp 1701704242
transform 1 0 8924 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_121
timestamp 1701704242
transform 1 0 11684 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_134
timestamp 1701704242
transform 1 0 12880 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_141
timestamp 1701704242
transform 1 0 13524 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_145
timestamp 1701704242
transform 1 0 13892 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_163
timestamp 1701704242
transform 1 0 15548 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_175
timestamp 1701704242
transform 1 0 16652 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_197
timestamp 1701704242
transform 1 0 18676 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_205
timestamp 1701704242
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_234
timestamp 1701704242
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1701704242
transform 1 0 23828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1701704242
transform 1 0 24932 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1701704242
transform 1 0 26036 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1701704242
transform 1 0 27140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1701704242
transform 1 0 28244 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1701704242
transform 1 0 28796 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1701704242
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_321
timestamp 1701704242
transform 1 0 30084 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_329
timestamp 1701704242
transform 1 0 30820 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1701704242
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1701704242
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1701704242
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1701704242
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1701704242
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1701704242
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1701704242
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1701704242
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_81
timestamp 1701704242
transform 1 0 8004 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_89
timestamp 1701704242
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_108
timestamp 1701704242
transform 1 0 10488 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_122
timestamp 1701704242
transform 1 0 11776 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_160
timestamp 1701704242
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1701704242
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 1701704242
transform 1 0 16100 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_173
timestamp 1701704242
transform 1 0 16468 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_177
timestamp 1701704242
transform 1 0 16836 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_198
timestamp 1701704242
transform 1 0 18768 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_205
timestamp 1701704242
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1701704242
transform 1 0 20976 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_225
timestamp 1701704242
transform 1 0 21252 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_265
timestamp 1701704242
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_277
timestamp 1701704242
transform 1 0 26036 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1701704242
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1701704242
transform 1 0 27508 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1701704242
transform 1 0 28612 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1701704242
transform 1 0 29716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_329
timestamp 1701704242
transform 1 0 30820 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1701704242
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1701704242
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1701704242
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1701704242
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1701704242
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1701704242
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1701704242
transform 1 0 6532 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1701704242
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1701704242
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1701704242
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_97
timestamp 1701704242
transform 1 0 9476 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_101
timestamp 1701704242
transform 1 0 9844 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_122
timestamp 1701704242
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_136
timestamp 1701704242
transform 1 0 13064 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1701704242
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_153
timestamp 1701704242
transform 1 0 14628 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1701704242
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1701704242
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1701704242
transform 1 0 24932 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1701704242
transform 1 0 26036 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1701704242
transform 1 0 27140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1701704242
transform 1 0 28244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1701704242
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1701704242
transform 1 0 28980 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_321
timestamp 1701704242
transform 1 0 30084 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_329
timestamp 1701704242
transform 1 0 30820 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1701704242
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1701704242
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1701704242
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1701704242
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1701704242
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1701704242
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1701704242
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1701704242
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1701704242
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1701704242
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_105
timestamp 1701704242
transform 1 0 10212 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_116
timestamp 1701704242
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_124
timestamp 1701704242
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_138
timestamp 1701704242
transform 1 0 13248 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_148
timestamp 1701704242
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_172
timestamp 1701704242
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_177
timestamp 1701704242
transform 1 0 16836 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_184
timestamp 1701704242
transform 1 0 17480 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_202
timestamp 1701704242
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1701704242
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1701704242
transform 1 0 22356 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1701704242
transform 1 0 23460 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1701704242
transform 1 0 24564 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1701704242
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1701704242
transform 1 0 26220 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1701704242
transform 1 0 26404 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1701704242
transform 1 0 27508 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1701704242
transform 1 0 28612 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1701704242
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_329
timestamp 1701704242
transform 1 0 30820 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1701704242
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1701704242
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1701704242
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1701704242
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1701704242
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1701704242
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1701704242
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1701704242
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1701704242
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1701704242
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1701704242
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_109
timestamp 1701704242
transform 1 0 10580 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_136
timestamp 1701704242
transform 1 0 13064 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_141
timestamp 1701704242
transform 1 0 13524 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_148
timestamp 1701704242
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_153
timestamp 1701704242
transform 1 0 14628 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_157
timestamp 1701704242
transform 1 0 14996 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_161
timestamp 1701704242
transform 1 0 15364 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_169
timestamp 1701704242
transform 1 0 16100 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_214
timestamp 1701704242
transform 1 0 20240 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1701704242
transform 1 0 20884 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1701704242
transform 1 0 21988 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1701704242
transform 1 0 23092 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1701704242
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1701704242
transform 1 0 23828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1701704242
transform 1 0 24932 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1701704242
transform 1 0 26036 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1701704242
transform 1 0 27140 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1701704242
transform 1 0 28244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1701704242
transform 1 0 28796 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1701704242
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_321
timestamp 1701704242
transform 1 0 30084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_329
timestamp 1701704242
transform 1 0 30820 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1701704242
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1701704242
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1701704242
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1701704242
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1701704242
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1701704242
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1701704242
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1701704242
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1701704242
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1701704242
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1701704242
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1701704242
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1701704242
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_125
timestamp 1701704242
transform 1 0 12052 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_133
timestamp 1701704242
transform 1 0 12788 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1701704242
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1701704242
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_196
timestamp 1701704242
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_208
timestamp 1701704242
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_220
timestamp 1701704242
transform 1 0 20792 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1701704242
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1701704242
transform 1 0 22356 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1701704242
transform 1 0 23460 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1701704242
transform 1 0 24564 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1701704242
transform 1 0 25668 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1701704242
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1701704242
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1701704242
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1701704242
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1701704242
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_329
timestamp 1701704242
transform 1 0 30820 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1701704242
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1701704242
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1701704242
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1701704242
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1701704242
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1701704242
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1701704242
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1701704242
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1701704242
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1701704242
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1701704242
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1701704242
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1701704242
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1701704242
transform 1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1701704242
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1701704242
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1701704242
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1701704242
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1701704242
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1701704242
transform 1 0 17940 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1701704242
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1701704242
transform 1 0 18676 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1701704242
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1701704242
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1701704242
transform 1 0 21988 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1701704242
transform 1 0 23092 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1701704242
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1701704242
transform 1 0 23828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1701704242
transform 1 0 24932 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1701704242
transform 1 0 26036 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1701704242
transform 1 0 27140 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1701704242
transform 1 0 28244 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1701704242
transform 1 0 28796 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1701704242
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1701704242
transform 1 0 30084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_329
timestamp 1701704242
transform 1 0 30820 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1701704242
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1701704242
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1701704242
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1701704242
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1701704242
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1701704242
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1701704242
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1701704242
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1701704242
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1701704242
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1701704242
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1701704242
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1701704242
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1701704242
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1701704242
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1701704242
transform 1 0 14260 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1701704242
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1701704242
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1701704242
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1701704242
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1701704242
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1701704242
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1701704242
transform 1 0 20516 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1701704242
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1701704242
transform 1 0 21252 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1701704242
transform 1 0 22356 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1701704242
transform 1 0 23460 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1701704242
transform 1 0 24564 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1701704242
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1701704242
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1701704242
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1701704242
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1701704242
transform 1 0 28612 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1701704242
transform 1 0 29716 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_329
timestamp 1701704242
transform 1 0 30820 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1701704242
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1701704242
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1701704242
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1701704242
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1701704242
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1701704242
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1701704242
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1701704242
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1701704242
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1701704242
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1701704242
transform 1 0 9476 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1701704242
transform 1 0 10580 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1701704242
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1701704242
transform 1 0 12788 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1701704242
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1701704242
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1701704242
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1701704242
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1701704242
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1701704242
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1701704242
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1701704242
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1701704242
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1701704242
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1701704242
transform 1 0 21988 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1701704242
transform 1 0 23092 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1701704242
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1701704242
transform 1 0 23828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1701704242
transform 1 0 24932 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1701704242
transform 1 0 26036 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1701704242
transform 1 0 27140 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1701704242
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1701704242
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1701704242
transform 1 0 28980 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_321
timestamp 1701704242
transform 1 0 30084 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_329
timestamp 1701704242
transform 1 0 30820 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1701704242
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1701704242
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1701704242
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1701704242
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1701704242
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1701704242
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1701704242
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1701704242
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1701704242
transform 1 0 8004 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1701704242
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1701704242
transform 1 0 10212 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1701704242
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1701704242
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1701704242
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1701704242
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1701704242
transform 1 0 14260 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1701704242
transform 1 0 15364 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1701704242
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1701704242
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1701704242
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1701704242
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1701704242
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1701704242
transform 1 0 20516 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1701704242
transform 1 0 21068 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1701704242
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1701704242
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1701704242
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1701704242
transform 1 0 24564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1701704242
transform 1 0 25668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1701704242
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1701704242
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1701704242
transform 1 0 27508 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1701704242
transform 1 0 28612 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1701704242
transform 1 0 29716 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_329
timestamp 1701704242
transform 1 0 30820 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1701704242
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1701704242
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1701704242
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1701704242
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1701704242
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1701704242
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1701704242
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1701704242
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1701704242
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1701704242
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1701704242
transform 1 0 10580 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1701704242
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1701704242
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1701704242
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1701704242
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1701704242
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1701704242
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1701704242
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1701704242
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1701704242
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1701704242
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1701704242
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1701704242
transform 1 0 20884 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1701704242
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1701704242
transform 1 0 23092 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1701704242
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1701704242
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1701704242
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1701704242
transform 1 0 26036 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1701704242
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1701704242
transform 1 0 28244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1701704242
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1701704242
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_321
timestamp 1701704242
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_329
timestamp 1701704242
transform 1 0 30820 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1701704242
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1701704242
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1701704242
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1701704242
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1701704242
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1701704242
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1701704242
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1701704242
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1701704242
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1701704242
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1701704242
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1701704242
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1701704242
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1701704242
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1701704242
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1701704242
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1701704242
transform 1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1701704242
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1701704242
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1701704242
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1701704242
transform 1 0 18308 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1701704242
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1701704242
transform 1 0 20516 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1701704242
transform 1 0 21068 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1701704242
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1701704242
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1701704242
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1701704242
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1701704242
transform 1 0 25668 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1701704242
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1701704242
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1701704242
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1701704242
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1701704242
transform 1 0 29716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_329
timestamp 1701704242
transform 1 0 30820 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1701704242
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1701704242
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1701704242
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1701704242
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1701704242
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1701704242
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1701704242
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1701704242
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1701704242
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1701704242
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1701704242
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1701704242
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1701704242
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1701704242
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1701704242
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1701704242
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1701704242
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1701704242
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1701704242
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1701704242
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1701704242
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1701704242
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1701704242
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1701704242
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1701704242
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1701704242
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1701704242
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1701704242
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1701704242
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1701704242
transform 1 0 26036 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1701704242
transform 1 0 27140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1701704242
transform 1 0 28244 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1701704242
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1701704242
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1701704242
transform 1 0 30084 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_329
timestamp 1701704242
transform 1 0 30820 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1701704242
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1701704242
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_27
timestamp 1701704242
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1701704242
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1701704242
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1701704242
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1701704242
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1701704242
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1701704242
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_85
timestamp 1701704242
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1701704242
transform 1 0 9476 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1701704242
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1701704242
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1701704242
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_137
timestamp 1701704242
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_141
timestamp 1701704242
transform 1 0 13524 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_153
timestamp 1701704242
transform 1 0 14628 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1701704242
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1701704242
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1701704242
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_193
timestamp 1701704242
transform 1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_197
timestamp 1701704242
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_209
timestamp 1701704242
transform 1 0 19780 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1701704242
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1701704242
transform 1 0 21252 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1701704242
transform 1 0 22356 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_249
timestamp 1701704242
transform 1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1701704242
transform 1 0 23828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_265
timestamp 1701704242
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1701704242
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1701704242
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1701704242
transform 1 0 27508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_305
timestamp 1701704242
transform 1 0 28612 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_309
timestamp 1701704242
transform 1 0 28980 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_321
timestamp 1701704242
transform 1 0 30084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_329
timestamp 1701704242
transform 1 0 30820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[0\].dly_stg1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15732 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[0\].dly_stg2
timestamp 1701704242
transform 1 0 16652 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[1\].dly_stg1
timestamp 1701704242
transform -1 0 16652 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[1\].dly_stg2
timestamp 1701704242
transform 1 0 16376 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[2\].dly_stg1
timestamp 1701704242
transform -1 0 17572 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[2\].dly_stg2
timestamp 1701704242
transform -1 0 17296 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[3\].dly_stg1
timestamp 1701704242
transform 1 0 18216 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[3\].dly_stg2
timestamp 1701704242
transform -1 0 17940 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[4\].dly_stg1
timestamp 1701704242
transform 1 0 17940 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[4\].dly_stg2
timestamp 1701704242
transform 1 0 18216 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[5\].dly_stg1
timestamp 1701704242
transform -1 0 19320 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[5\].dly_stg2
timestamp 1701704242
transform -1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[6\].dly_stg1
timestamp 1701704242
transform 1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[6\].dly_stg2
timestamp 1701704242
transform -1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[7\].dly_stg1
timestamp 1701704242
transform -1 0 19872 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[7\].dly_stg2
timestamp 1701704242
transform 1 0 19872 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[8\].dly_stg1
timestamp 1701704242
transform -1 0 21252 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[8\].dly_stg2
timestamp 1701704242
transform 1 0 20700 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[9\].dly_stg1
timestamp 1701704242
transform 1 0 23184 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[9\].dly_stg2
timestamp 1701704242
transform -1 0 21804 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[10\].dly_stg1
timestamp 1701704242
transform 1 0 20332 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[10\].dly_stg2
timestamp 1701704242
transform 1 0 21252 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[11\].dly_stg1
timestamp 1701704242
transform -1 0 21160 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[11\].dly_stg2
timestamp 1701704242
transform -1 0 20608 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[12\].dly_stg1
timestamp 1701704242
transform -1 0 20056 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[12\].dly_stg2
timestamp 1701704242
transform 1 0 20056 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[13\].dly_stg1
timestamp 1701704242
transform -1 0 19780 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[13\].dly_stg2
timestamp 1701704242
transform -1 0 19504 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[14\].dly_stg1
timestamp 1701704242
transform -1 0 19228 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[14\].dly_stg2
timestamp 1701704242
transform -1 0 18952 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[15\].dly_stg1
timestamp 1701704242
transform -1 0 18400 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[15\].dly_stg2
timestamp 1701704242
transform -1 0 18124 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[16\].dly_stg1
timestamp 1701704242
transform -1 0 18216 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[16\].dly_stg2
timestamp 1701704242
transform -1 0 16836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[17\].dly_stg1
timestamp 1701704242
transform -1 0 16284 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[17\].dly_stg2
timestamp 1701704242
transform -1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[18\].dly_stg1
timestamp 1701704242
transform 1 0 15180 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[18\].dly_stg2
timestamp 1701704242
transform 1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[19\].dly_stg1
timestamp 1701704242
transform 1 0 14628 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[19\].dly_stg2
timestamp 1701704242
transform -1 0 14628 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[20\].dly_stg1
timestamp 1701704242
transform -1 0 14536 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[20\].dly_stg2
timestamp 1701704242
transform -1 0 14444 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[21\].dly_stg1
timestamp 1701704242
transform -1 0 13156 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[21\].dly_stg2
timestamp 1701704242
transform 1 0 13524 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[22\].dly_stg1
timestamp 1701704242
transform -1 0 14168 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[22\].dly_stg2
timestamp 1701704242
transform -1 0 13616 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[23\].dly_stg1
timestamp 1701704242
transform 1 0 13524 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[23\].dly_stg2
timestamp 1701704242
transform -1 0 14352 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[24\].dly_stg1
timestamp 1701704242
transform -1 0 13616 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[24\].dly_stg2
timestamp 1701704242
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[25\].dly_stg1
timestamp 1701704242
transform 1 0 13064 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[25\].dly_stg2
timestamp 1701704242
transform -1 0 13984 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[26\].dly_stg1
timestamp 1701704242
transform 1 0 12604 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[26\].dly_stg2
timestamp 1701704242
transform -1 0 13156 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[27\].dly_stg1
timestamp 1701704242
transform -1 0 12328 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[27\].dly_stg2
timestamp 1701704242
transform -1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[28\].dly_stg1
timestamp 1701704242
transform -1 0 12052 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[28\].dly_stg2
timestamp 1701704242
transform -1 0 11776 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[29\].dly_stg1
timestamp 1701704242
transform -1 0 10856 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[29\].dly_stg2
timestamp 1701704242
transform -1 0 11132 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[30\].dly_stg1
timestamp 1701704242
transform 1 0 9752 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[30\].dly_stg2
timestamp 1701704242
transform 1 0 10028 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[31\].dly_stg1
timestamp 1701704242
transform -1 0 9936 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[31\].dly_stg2
timestamp 1701704242
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[32\].dly_stg1
timestamp 1701704242
transform -1 0 9016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[32\].dly_stg2
timestamp 1701704242
transform 1 0 9936 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[33\].dly_stg1
timestamp 1701704242
transform 1 0 8004 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[33\].dly_stg2
timestamp 1701704242
transform -1 0 8464 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[34\].dly_stg1
timestamp 1701704242
transform -1 0 8280 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[34\].dly_stg2
timestamp 1701704242
transform -1 0 8004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[35\].dly_stg1
timestamp 1701704242
transform 1 0 8464 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[35\].dly_stg2
timestamp 1701704242
transform 1 0 9016 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[36\].dly_stg1
timestamp 1701704242
transform -1 0 8280 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[36\].dly_stg2
timestamp 1701704242
transform 1 0 9292 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[37\].dly_stg1
timestamp 1701704242
transform -1 0 9016 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[37\].dly_stg2
timestamp 1701704242
transform -1 0 9200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[38\].dly_stg1
timestamp 1701704242
transform 1 0 9752 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[38\].dly_stg2
timestamp 1701704242
transform -1 0 9752 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[39\].dly_stg1
timestamp 1701704242
transform -1 0 9660 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[39\].dly_stg2
timestamp 1701704242
transform -1 0 10212 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[40\].dly_stg1
timestamp 1701704242
transform -1 0 10212 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[40\].dly_stg2
timestamp 1701704242
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[41\].dly_stg1
timestamp 1701704242
transform -1 0 11224 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[41\].dly_stg2
timestamp 1701704242
transform -1 0 10488 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[42\].dly_stg1
timestamp 1701704242
transform -1 0 12328 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[42\].dly_stg2
timestamp 1701704242
transform -1 0 12604 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[43\].dly_stg1
timestamp 1701704242
transform -1 0 11776 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[43\].dly_stg2
timestamp 1701704242
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[44\].dly_stg1
timestamp 1701704242
transform -1 0 11776 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[44\].dly_stg2
timestamp 1701704242
transform -1 0 9568 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[45\].dly_stg1
timestamp 1701704242
transform 1 0 11684 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[45\].dly_stg2
timestamp 1701704242
transform 1 0 11960 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[46\].dly_stg1
timestamp 1701704242
transform 1 0 12788 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[46\].dly_stg2
timestamp 1701704242
transform -1 0 12788 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[47\].dly_stg1
timestamp 1701704242
transform -1 0 12972 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[47\].dly_stg2
timestamp 1701704242
transform -1 0 12696 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[48\].dly_stg1
timestamp 1701704242
transform 1 0 13892 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[48\].dly_stg2
timestamp 1701704242
transform -1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[49\].dly_stg1
timestamp 1701704242
transform -1 0 14628 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[49\].dly_stg2
timestamp 1701704242
transform 1 0 14720 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[50\].dly_stg1
timestamp 1701704242
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[50\].dly_stg2
timestamp 1701704242
transform 1 0 15548 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[51\].dly_stg1
timestamp 1701704242
transform 1 0 15732 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[51\].dly_stg2
timestamp 1701704242
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[52\].dly_stg1
timestamp 1701704242
transform -1 0 17480 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[52\].dly_stg2
timestamp 1701704242
transform -1 0 17204 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[53\].dly_stg1
timestamp 1701704242
transform 1 0 18676 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[53\].dly_stg2
timestamp 1701704242
transform -1 0 18584 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[54\].dly_stg1
timestamp 1701704242
transform -1 0 19228 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[54\].dly_stg2
timestamp 1701704242
transform -1 0 19504 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[55\].dly_stg1
timestamp 1701704242
transform 1 0 19136 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[55\].dly_stg2
timestamp 1701704242
transform 1 0 20056 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[56\].dly_stg1
timestamp 1701704242
transform -1 0 19596 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[56\].dly_stg2
timestamp 1701704242
transform -1 0 20608 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[57\].dly_stg1
timestamp 1701704242
transform 1 0 19872 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[57\].dly_stg2
timestamp 1701704242
transform 1 0 20148 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[58\].dly_stg1
timestamp 1701704242
transform -1 0 20700 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[58\].dly_stg2
timestamp 1701704242
transform -1 0 20148 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[59\].dly_stg1
timestamp 1701704242
transform 1 0 21528 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[59\].dly_stg2
timestamp 1701704242
transform -1 0 21528 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[60\].dly_stg1
timestamp 1701704242
transform 1 0 21804 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[60\].dly_stg2
timestamp 1701704242
transform -1 0 21068 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[61\].dly_stg1
timestamp 1701704242
transform -1 0 22632 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[61\].dly_stg2
timestamp 1701704242
transform -1 0 22356 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[62\].dly_stg1
timestamp 1701704242
transform -1 0 22448 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[62\].dly_stg2
timestamp 1701704242
transform -1 0 22724 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[63\].dly_stg1
timestamp 1701704242
transform -1 0 22080 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[63\].dly_stg2
timestamp 1701704242
transform -1 0 21528 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[64\].dly_stg1
timestamp 1701704242
transform 1 0 22724 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_even\[64\].dly_stg2
timestamp 1701704242
transform -1 0 21804 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg1
timestamp 1701704242
transform 1 0 15732 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg2
timestamp 1701704242
transform -1 0 16560 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg1
timestamp 1701704242
transform 1 0 18492 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg2
timestamp 1701704242
transform -1 0 16376 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg1
timestamp 1701704242
transform 1 0 17940 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg2
timestamp 1701704242
transform -1 0 17020 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg1
timestamp 1701704242
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg2
timestamp 1701704242
transform 1 0 18768 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg1
timestamp 1701704242
transform 1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg2
timestamp 1701704242
transform 1 0 18584 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg1
timestamp 1701704242
transform 1 0 19964 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg2
timestamp 1701704242
transform 1 0 19688 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg1
timestamp 1701704242
transform 1 0 19320 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg2
timestamp 1701704242
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg1
timestamp 1701704242
transform 1 0 20792 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg2
timestamp 1701704242
transform 1 0 20424 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg1
timestamp 1701704242
transform 1 0 21252 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg2
timestamp 1701704242
transform -1 0 20332 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg1
timestamp 1701704242
transform -1 0 20424 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg2
timestamp 1701704242
transform -1 0 21804 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg1
timestamp 1701704242
transform -1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg2
timestamp 1701704242
transform -1 0 19504 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg1
timestamp 1701704242
transform -1 0 19780 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg2
timestamp 1701704242
transform -1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg1
timestamp 1701704242
transform -1 0 18124 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg2
timestamp 1701704242
transform -1 0 20056 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg1
timestamp 1701704242
transform -1 0 18676 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg2
timestamp 1701704242
transform -1 0 18400 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[14\].dly_stg1
timestamp 1701704242
transform -1 0 18952 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[14\].dly_stg2
timestamp 1701704242
transform 1 0 18952 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[15\].dly_stg1
timestamp 1701704242
transform -1 0 17388 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[15\].dly_stg2
timestamp 1701704242
transform -1 0 17848 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[16\].dly_stg1
timestamp 1701704242
transform -1 0 16560 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[16\].dly_stg2
timestamp 1701704242
transform -1 0 17112 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[17\].dly_stg1
timestamp 1701704242
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[17\].dly_stg2
timestamp 1701704242
transform -1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[18\].dly_stg1
timestamp 1701704242
transform -1 0 15180 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[18\].dly_stg2
timestamp 1701704242
transform -1 0 15456 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[19\].dly_stg1
timestamp 1701704242
transform -1 0 14720 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[19\].dly_stg2
timestamp 1701704242
transform -1 0 14996 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[20\].dly_stg1
timestamp 1701704242
transform -1 0 13340 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[20\].dly_stg2
timestamp 1701704242
transform 1 0 14996 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[21\].dly_stg1
timestamp 1701704242
transform -1 0 13892 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[21\].dly_stg2
timestamp 1701704242
transform -1 0 12880 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[22\].dly_stg1
timestamp 1701704242
transform -1 0 14444 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[22\].dly_stg2
timestamp 1701704242
transform -1 0 14076 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[23\].dly_stg1
timestamp 1701704242
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[23\].dly_stg2
timestamp 1701704242
transform 1 0 14352 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[24\].dly_stg1
timestamp 1701704242
transform -1 0 13892 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[24\].dly_stg2
timestamp 1701704242
transform -1 0 14168 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[25\].dly_stg1
timestamp 1701704242
transform -1 0 13064 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[25\].dly_stg2
timestamp 1701704242
transform 1 0 13984 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[26\].dly_stg1
timestamp 1701704242
transform -1 0 12604 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[26\].dly_stg2
timestamp 1701704242
transform 1 0 13156 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[27\].dly_stg1
timestamp 1701704242
transform -1 0 12328 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[27\].dly_stg2
timestamp 1701704242
transform 1 0 12328 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[28\].dly_stg1
timestamp 1701704242
transform -1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[28\].dly_stg2
timestamp 1701704242
transform -1 0 11500 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[29\].dly_stg1
timestamp 1701704242
transform -1 0 10580 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[29\].dly_stg2
timestamp 1701704242
transform -1 0 10764 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[30\].dly_stg1
timestamp 1701704242
transform -1 0 9568 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[30\].dly_stg2
timestamp 1701704242
transform -1 0 10488 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[31\].dly_stg1
timestamp 1701704242
transform -1 0 7728 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[31\].dly_stg2
timestamp 1701704242
transform -1 0 8004 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[32\].dly_stg1
timestamp 1701704242
transform -1 0 9016 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[32\].dly_stg2
timestamp 1701704242
transform -1 0 8740 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[33\].dly_stg1
timestamp 1701704242
transform -1 0 9660 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[33\].dly_stg2
timestamp 1701704242
transform -1 0 8648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[34\].dly_stg1
timestamp 1701704242
transform -1 0 8832 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[34\].dly_stg2
timestamp 1701704242
transform -1 0 9108 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[35\].dly_stg1
timestamp 1701704242
transform -1 0 8464 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[35\].dly_stg2
timestamp 1701704242
transform -1 0 9016 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[36\].dly_stg1
timestamp 1701704242
transform -1 0 9292 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[36\].dly_stg2
timestamp 1701704242
transform -1 0 8648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[37\].dly_stg1
timestamp 1701704242
transform -1 0 10304 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[37\].dly_stg2
timestamp 1701704242
transform -1 0 8924 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[38\].dly_stg1
timestamp 1701704242
transform 1 0 9108 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[38\].dly_stg2
timestamp 1701704242
transform 1 0 9660 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[39\].dly_stg1
timestamp 1701704242
transform 1 0 9016 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[39\].dly_stg2
timestamp 1701704242
transform 1 0 10212 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[40\].dly_stg1
timestamp 1701704242
transform -1 0 10764 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[40\].dly_stg2
timestamp 1701704242
transform 1 0 9568 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[41\].dly_stg1
timestamp 1701704242
transform 1 0 11776 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[41\].dly_stg2
timestamp 1701704242
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[42\].dly_stg1
timestamp 1701704242
transform -1 0 11500 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[42\].dly_stg2
timestamp 1701704242
transform 1 0 12604 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[43\].dly_stg1
timestamp 1701704242
transform -1 0 10856 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[43\].dly_stg2
timestamp 1701704242
transform -1 0 10856 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[44\].dly_stg1
timestamp 1701704242
transform -1 0 12144 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[44\].dly_stg2
timestamp 1701704242
transform 1 0 10948 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[45\].dly_stg1
timestamp 1701704242
transform -1 0 11684 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[45\].dly_stg2
timestamp 1701704242
transform 1 0 12236 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[46\].dly_stg1
timestamp 1701704242
transform 1 0 12144 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[46\].dly_stg2
timestamp 1701704242
transform -1 0 11500 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[47\].dly_stg1
timestamp 1701704242
transform 1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[47\].dly_stg2
timestamp 1701704242
transform 1 0 12972 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[48\].dly_stg1
timestamp 1701704242
transform 1 0 13340 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[48\].dly_stg2
timestamp 1701704242
transform 1 0 14352 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[49\].dly_stg1
timestamp 1701704242
transform 1 0 14628 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[49\].dly_stg2
timestamp 1701704242
transform 1 0 15088 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[50\].dly_stg1
timestamp 1701704242
transform 1 0 15180 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[50\].dly_stg2
timestamp 1701704242
transform 1 0 15456 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[51\].dly_stg1
timestamp 1701704242
transform 1 0 16560 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[51\].dly_stg2
timestamp 1701704242
transform 1 0 16192 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[52\].dly_stg1
timestamp 1701704242
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[52\].dly_stg2
timestamp 1701704242
transform 1 0 17756 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[53\].dly_stg1
timestamp 1701704242
transform 1 0 18124 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[53\].dly_stg2
timestamp 1701704242
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[54\].dly_stg1
timestamp 1701704242
transform 1 0 19780 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[54\].dly_stg2
timestamp 1701704242
transform 1 0 19504 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[55\].dly_stg1
timestamp 1701704242
transform 1 0 20608 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[55\].dly_stg2
timestamp 1701704242
transform 1 0 20332 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[56\].dly_stg1
timestamp 1701704242
transform -1 0 20700 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[56\].dly_stg2
timestamp 1701704242
transform 1 0 20700 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[57\].dly_stg1
timestamp 1701704242
transform -1 0 19872 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[57\].dly_stg2
timestamp 1701704242
transform -1 0 20424 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[58\].dly_stg1
timestamp 1701704242
transform 1 0 20700 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[58\].dly_stg2
timestamp 1701704242
transform -1 0 19872 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[59\].dly_stg1
timestamp 1701704242
transform -1 0 21252 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[59\].dly_stg2
timestamp 1701704242
transform 1 0 21804 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[60\].dly_stg1
timestamp 1701704242
transform 1 0 21528 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[60\].dly_stg2
timestamp 1701704242
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[61\].dly_stg1
timestamp 1701704242
transform 1 0 22632 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[61\].dly_stg2
timestamp 1701704242
transform 1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[62\].dly_stg1
timestamp 1701704242
transform -1 0 22172 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[62\].dly_stg2
timestamp 1701704242
transform -1 0 22356 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[63\].dly_stg1
timestamp 1701704242
transform -1 0 22908 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[63\].dly_stg2
timestamp 1701704242
transform 1 0 22356 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 22632 0 1 544
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 31372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 31372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 31372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 31372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 31372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 31372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 31372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 31372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 31372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 31372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 31372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 31372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 31372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 31372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 31372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 31372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 31372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 31372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1701704242
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 31372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1701704242
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 31372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1701704242
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 31372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1701704242
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 31372 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1701704242
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 31372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1701704242
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 31372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1701704242
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 31372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1701704242
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 31372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1701704242
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 31372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1701704242
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 31372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1701704242
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 31372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1701704242
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 31372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1701704242
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 31372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1701704242
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1701704242
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1701704242
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1701704242
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1701704242
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1701704242
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1701704242
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1701704242
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1701704242
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_82
timestamp 1701704242
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp 1701704242
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 1701704242
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 1701704242
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 1701704242
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 1701704242
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 1701704242
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp 1701704242
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 1701704242
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_97
timestamp 1701704242
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 1701704242
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 1701704242
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 1701704242
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_101
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_103
timestamp 1701704242
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_104
timestamp 1701704242
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_105
timestamp 1701704242
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_108
timestamp 1701704242
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_109
timestamp 1701704242
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_110
timestamp 1701704242
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_111
timestamp 1701704242
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_112
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_113
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_114
timestamp 1701704242
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_115
timestamp 1701704242
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1701704242
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_117
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_118
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_119
timestamp 1701704242
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1701704242
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1701704242
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1701704242
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_123
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1701704242
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1701704242
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1701704242
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1701704242
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1701704242
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_132
timestamp 1701704242
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_133
timestamp 1701704242
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp 1701704242
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp 1701704242
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp 1701704242
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_140
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_141
timestamp 1701704242
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_142
timestamp 1701704242
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_143
timestamp 1701704242
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_144
timestamp 1701704242
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_145
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_146
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_147
timestamp 1701704242
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_148
timestamp 1701704242
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_149
timestamp 1701704242
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_150
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_152
timestamp 1701704242
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_153
timestamp 1701704242
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_154
timestamp 1701704242
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_155
timestamp 1701704242
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_156
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_157
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_158
timestamp 1701704242
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_159
timestamp 1701704242
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 1701704242
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_162
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_163
timestamp 1701704242
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 1701704242
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 1701704242
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 1701704242
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_167
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_168
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 1701704242
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_170
timestamp 1701704242
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 1701704242
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_172
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 1701704242
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 1701704242
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 1701704242
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 1701704242
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 1701704242
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 1701704242
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 1701704242
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_183
timestamp 1701704242
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_184
timestamp 1701704242
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_185
timestamp 1701704242
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 1701704242
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 1701704242
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 1701704242
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 1701704242
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_190
timestamp 1701704242
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_191
timestamp 1701704242
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_192
timestamp 1701704242
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 1701704242
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_194
timestamp 1701704242
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1701704242
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 1701704242
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 1701704242
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 1701704242
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 1701704242
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_200
timestamp 1701704242
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_201
timestamp 1701704242
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 1701704242
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 1701704242
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 1701704242
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_205
timestamp 1701704242
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 1701704242
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 1701704242
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 1701704242
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_209
timestamp 1701704242
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_210
timestamp 1701704242
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 1701704242
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 1701704242
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_213
timestamp 1701704242
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_214
timestamp 1701704242
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_215
timestamp 1701704242
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 1701704242
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 1701704242
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_218
timestamp 1701704242
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_219
timestamp 1701704242
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_220
timestamp 1701704242
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_221
timestamp 1701704242
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_222
timestamp 1701704242
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_223
timestamp 1701704242
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_224
timestamp 1701704242
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_225
timestamp 1701704242
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_226
timestamp 1701704242
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_227
timestamp 1701704242
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_228
timestamp 1701704242
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_229
timestamp 1701704242
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_230
timestamp 1701704242
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_231
timestamp 1701704242
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_232
timestamp 1701704242
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_233
timestamp 1701704242
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_234
timestamp 1701704242
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_235
timestamp 1701704242
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_236
timestamp 1701704242
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_237
timestamp 1701704242
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_238
timestamp 1701704242
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_239
timestamp 1701704242
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_240
timestamp 1701704242
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_241
timestamp 1701704242
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_242
timestamp 1701704242
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_243
timestamp 1701704242
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_244
timestamp 1701704242
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_245
timestamp 1701704242
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_246
timestamp 1701704242
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_247
timestamp 1701704242
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_248
timestamp 1701704242
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_249
timestamp 1701704242
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_250
timestamp 1701704242
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_251
timestamp 1701704242
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_252
timestamp 1701704242
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_253
timestamp 1701704242
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_254
timestamp 1701704242
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_255
timestamp 1701704242
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_256
timestamp 1701704242
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_257
timestamp 1701704242
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_258
timestamp 1701704242
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_259
timestamp 1701704242
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_260
timestamp 1701704242
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_261
timestamp 1701704242
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_262
timestamp 1701704242
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_263
timestamp 1701704242
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp 1701704242
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1701704242
transform 1 0 28888 0 -1 19040
box -38 -48 130 592
<< labels >>
flabel metal4 s 8096 496 8416 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15801 496 16121 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23506 496 23826 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 31211 496 31531 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4244 496 4564 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11949 496 12269 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19654 496 19974 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 27359 496 27679 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 22558 0 22614 400 0 FreeSans 224 90 0 0 i_start
port 2 nsew signal input
flabel metal2 s 7102 0 7158 400 0 FreeSans 224 90 0 0 i_stop
port 3 nsew signal input
flabel metal2 s 21270 0 21326 400 0 FreeSans 224 90 0 0 o_result[0]
port 4 nsew signal tristate
flabel metal3 s 31600 5448 32000 5568 0 FreeSans 480 0 0 0 o_result[10]
port 5 nsew signal tristate
flabel metal2 s 19982 0 20038 400 0 FreeSans 224 90 0 0 o_result[11]
port 6 nsew signal tristate
flabel metal3 s 31600 8848 32000 8968 0 FreeSans 480 0 0 0 o_result[12]
port 7 nsew signal tristate
flabel metal3 s 31600 9528 32000 9648 0 FreeSans 480 0 0 0 o_result[13]
port 8 nsew signal tristate
flabel metal2 s 18694 0 18750 400 0 FreeSans 224 90 0 0 o_result[14]
port 9 nsew signal tristate
flabel metal3 s 31600 10208 32000 10328 0 FreeSans 480 0 0 0 o_result[15]
port 10 nsew signal tristate
flabel metal2 s 21270 19600 21326 20000 0 FreeSans 224 90 0 0 o_result[16]
port 11 nsew signal tristate
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 224 90 0 0 o_result[17]
port 12 nsew signal tristate
flabel metal2 s 16118 19600 16174 20000 0 FreeSans 224 90 0 0 o_result[18]
port 13 nsew signal tristate
flabel metal2 s 9034 0 9090 400 0 FreeSans 224 90 0 0 o_result[19]
port 14 nsew signal tristate
flabel metal2 s 14186 0 14242 400 0 FreeSans 224 90 0 0 o_result[1]
port 15 nsew signal tristate
flabel metal2 s 10322 0 10378 400 0 FreeSans 224 90 0 0 o_result[20]
port 16 nsew signal tristate
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 o_result[21]
port 17 nsew signal tristate
flabel metal2 s 11610 0 11666 400 0 FreeSans 224 90 0 0 o_result[22]
port 18 nsew signal tristate
flabel metal2 s 16118 0 16174 400 0 FreeSans 224 90 0 0 o_result[23]
port 19 nsew signal tristate
flabel metal2 s 17406 0 17462 400 0 FreeSans 224 90 0 0 o_result[24]
port 20 nsew signal tristate
flabel metal2 s 12898 0 12954 400 0 FreeSans 224 90 0 0 o_result[25]
port 21 nsew signal tristate
flabel metal2 s 14830 0 14886 400 0 FreeSans 224 90 0 0 o_result[26]
port 22 nsew signal tristate
flabel metal2 s 13542 0 13598 400 0 FreeSans 224 90 0 0 o_result[27]
port 23 nsew signal tristate
flabel metal2 s 12254 0 12310 400 0 FreeSans 224 90 0 0 o_result[28]
port 24 nsew signal tristate
flabel metal2 s 9678 0 9734 400 0 FreeSans 224 90 0 0 o_result[29]
port 25 nsew signal tristate
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 o_result[2]
port 26 nsew signal tristate
flabel metal3 s 0 6128 400 6248 0 FreeSans 480 0 0 0 o_result[30]
port 27 nsew signal tristate
flabel metal2 s 10966 0 11022 400 0 FreeSans 224 90 0 0 o_result[31]
port 28 nsew signal tristate
flabel metal3 s 0 6808 400 6928 0 FreeSans 480 0 0 0 o_result[32]
port 29 nsew signal tristate
flabel metal3 s 0 7488 400 7608 0 FreeSans 480 0 0 0 o_result[33]
port 30 nsew signal tristate
flabel metal3 s 0 8848 400 8968 0 FreeSans 480 0 0 0 o_result[34]
port 31 nsew signal tristate
flabel metal3 s 0 8168 400 8288 0 FreeSans 480 0 0 0 o_result[35]
port 32 nsew signal tristate
flabel metal3 s 0 9528 400 9648 0 FreeSans 480 0 0 0 o_result[36]
port 33 nsew signal tristate
flabel metal3 s 0 10208 400 10328 0 FreeSans 480 0 0 0 o_result[37]
port 34 nsew signal tristate
flabel metal3 s 0 11568 400 11688 0 FreeSans 480 0 0 0 o_result[38]
port 35 nsew signal tristate
flabel metal3 s 0 10888 400 11008 0 FreeSans 480 0 0 0 o_result[39]
port 36 nsew signal tristate
flabel metal2 s 18050 0 18106 400 0 FreeSans 224 90 0 0 o_result[3]
port 37 nsew signal tristate
flabel metal2 s 11610 19600 11666 20000 0 FreeSans 224 90 0 0 o_result[40]
port 38 nsew signal tristate
flabel metal2 s 13542 19600 13598 20000 0 FreeSans 224 90 0 0 o_result[41]
port 39 nsew signal tristate
flabel metal2 s 15474 19600 15530 20000 0 FreeSans 224 90 0 0 o_result[42]
port 40 nsew signal tristate
flabel metal2 s 12898 19600 12954 20000 0 FreeSans 224 90 0 0 o_result[43]
port 41 nsew signal tristate
flabel metal3 s 0 12248 400 12368 0 FreeSans 480 0 0 0 o_result[44]
port 42 nsew signal tristate
flabel metal2 s 10966 19600 11022 20000 0 FreeSans 224 90 0 0 o_result[45]
port 43 nsew signal tristate
flabel metal2 s 14830 19600 14886 20000 0 FreeSans 224 90 0 0 o_result[46]
port 44 nsew signal tristate
flabel metal2 s 12254 19600 12310 20000 0 FreeSans 224 90 0 0 o_result[47]
port 45 nsew signal tristate
flabel metal2 s 14186 19600 14242 20000 0 FreeSans 224 90 0 0 o_result[48]
port 46 nsew signal tristate
flabel metal2 s 16762 19600 16818 20000 0 FreeSans 224 90 0 0 o_result[49]
port 47 nsew signal tristate
flabel metal2 s 20626 0 20682 400 0 FreeSans 224 90 0 0 o_result[4]
port 48 nsew signal tristate
flabel metal2 s 18050 19600 18106 20000 0 FreeSans 224 90 0 0 o_result[50]
port 49 nsew signal tristate
flabel metal2 s 19982 19600 20038 20000 0 FreeSans 224 90 0 0 o_result[51]
port 50 nsew signal tristate
flabel metal2 s 18694 19600 18750 20000 0 FreeSans 224 90 0 0 o_result[52]
port 51 nsew signal tristate
flabel metal2 s 20626 19600 20682 20000 0 FreeSans 224 90 0 0 o_result[53]
port 52 nsew signal tristate
flabel metal2 s 21914 19600 21970 20000 0 FreeSans 224 90 0 0 o_result[54]
port 53 nsew signal tristate
flabel metal3 s 31600 14968 32000 15088 0 FreeSans 480 0 0 0 o_result[55]
port 54 nsew signal tristate
flabel metal3 s 31600 12928 32000 13048 0 FreeSans 480 0 0 0 o_result[56]
port 55 nsew signal tristate
flabel metal3 s 31600 14288 32000 14408 0 FreeSans 480 0 0 0 o_result[57]
port 56 nsew signal tristate
flabel metal2 s 19338 19600 19394 20000 0 FreeSans 224 90 0 0 o_result[58]
port 57 nsew signal tristate
flabel metal3 s 31600 12248 32000 12368 0 FreeSans 480 0 0 0 o_result[59]
port 58 nsew signal tristate
flabel metal2 s 19338 0 19394 400 0 FreeSans 224 90 0 0 o_result[5]
port 59 nsew signal tristate
flabel metal3 s 31600 13608 32000 13728 0 FreeSans 480 0 0 0 o_result[60]
port 60 nsew signal tristate
flabel metal3 s 31600 11568 32000 11688 0 FreeSans 480 0 0 0 o_result[61]
port 61 nsew signal tristate
flabel metal3 s 31600 10888 32000 11008 0 FreeSans 480 0 0 0 o_result[62]
port 62 nsew signal tristate
flabel metal3 s 31600 8168 32000 8288 0 FreeSans 480 0 0 0 o_result[63]
port 63 nsew signal tristate
flabel metal2 s 21914 0 21970 400 0 FreeSans 224 90 0 0 o_result[6]
port 64 nsew signal tristate
flabel metal3 s 31600 6128 32000 6248 0 FreeSans 480 0 0 0 o_result[7]
port 65 nsew signal tristate
flabel metal3 s 31600 6808 32000 6928 0 FreeSans 480 0 0 0 o_result[8]
port 66 nsew signal tristate
flabel metal3 s 31600 7488 32000 7608 0 FreeSans 480 0 0 0 o_result[9]
port 67 nsew signal tristate
rlabel via1 16041 19040 16041 19040 0 VGND
rlabel metal1 15962 18496 15962 18496 0 VPWR
rlabel metal1 17296 12274 17296 12274 0 clknet_0_i_stop
rlabel metal1 10488 6222 10488 6222 0 clknet_3_0__leaf_i_stop
rlabel metal1 14628 6222 14628 6222 0 clknet_3_1__leaf_i_stop
rlabel metal1 11408 12750 11408 12750 0 clknet_3_2__leaf_i_stop
rlabel metal1 14490 14484 14490 14484 0 clknet_3_3__leaf_i_stop
rlabel metal1 17066 6732 17066 6732 0 clknet_3_4__leaf_i_stop
rlabel metal1 21206 8942 21206 8942 0 clknet_3_5__leaf_i_stop
rlabel metal1 17618 13396 17618 13396 0 clknet_3_6__leaf_i_stop
rlabel metal1 20332 12818 20332 12818 0 clknet_3_7__leaf_i_stop
rlabel metal2 22586 415 22586 415 0 i_start
rlabel metal1 14306 10132 14306 10132 0 i_stop
rlabel metal1 16284 5134 16284 5134 0 net1
rlabel metal2 21298 2676 21298 2676 0 o_result[0]
rlabel metal2 28474 7157 28474 7157 0 o_result[10]
rlabel metal1 19596 7718 19596 7718 0 o_result[11]
rlabel metal2 28290 8721 28290 8721 0 o_result[12]
rlabel metal1 22218 9418 22218 9418 0 o_result[13]
rlabel metal1 18170 8806 18170 8806 0 o_result[14]
rlabel metal2 20930 9792 20930 9792 0 o_result[15]
rlabel metal1 19872 10778 19872 10778 0 o_result[16]
rlabel metal1 17480 11322 17480 11322 0 o_result[17]
rlabel metal2 16192 19244 16192 19244 0 o_result[18]
rlabel metal2 12650 6664 12650 6664 0 o_result[19]
rlabel metal1 14076 5542 14076 5542 0 o_result[1]
rlabel metal1 10810 4114 10810 4114 0 o_result[20]
rlabel metal1 15686 8806 15686 8806 0 o_result[21]
rlabel metal2 11638 1557 11638 1557 0 o_result[22]
rlabel metal1 16192 8262 16192 8262 0 o_result[23]
rlabel metal2 17434 1571 17434 1571 0 o_result[24]
rlabel metal1 13708 6970 13708 6970 0 o_result[25]
rlabel metal2 14858 1557 14858 1557 0 o_result[26]
rlabel metal1 13432 6086 13432 6086 0 o_result[27]
rlabel metal2 12282 619 12282 619 0 o_result[28]
rlabel metal1 9384 6086 9384 6086 0 o_result[29]
rlabel metal1 16376 6086 16376 6086 0 o_result[2]
rlabel metal2 7866 6409 7866 6409 0 o_result[30]
rlabel metal1 11040 7718 11040 7718 0 o_result[31]
rlabel metal2 6670 7293 6670 7293 0 o_result[32]
rlabel metal3 1533 7548 1533 7548 0 o_result[33]
rlabel via2 6762 8891 6762 8891 0 o_result[34]
rlabel metal3 1533 8228 1533 8228 0 o_result[35]
rlabel via2 9798 9605 9798 9605 0 o_result[36]
rlabel via2 7130 10251 7130 10251 0 o_result[37]
rlabel metal1 7544 11322 7544 11322 0 o_result[38]
rlabel metal3 1533 10948 1533 10948 0 o_result[39]
rlabel metal2 17986 6460 17986 6460 0 o_result[3]
rlabel metal1 11500 11322 11500 11322 0 o_result[40]
rlabel metal1 13892 11322 13892 11322 0 o_result[41]
rlabel metal1 15456 11866 15456 11866 0 o_result[42]
rlabel metal1 13248 12410 13248 12410 0 o_result[43]
rlabel metal2 6946 12359 6946 12359 0 o_result[44]
rlabel metal2 10994 18099 10994 18099 0 o_result[45]
rlabel metal1 14996 12410 14996 12410 0 o_result[46]
rlabel metal2 12328 18700 12328 18700 0 o_result[47]
rlabel metal1 14260 14586 14260 14586 0 o_result[48]
rlabel metal1 16330 14586 16330 14586 0 o_result[49]
rlabel metal1 20332 6086 20332 6086 0 o_result[4]
rlabel metal1 17848 14042 17848 14042 0 o_result[50]
rlabel metal1 19504 13498 19504 13498 0 o_result[51]
rlabel metal1 18262 12954 18262 12954 0 o_result[52]
rlabel metal1 20378 14042 20378 14042 0 o_result[53]
rlabel metal1 21482 13498 21482 13498 0 o_result[54]
rlabel metal2 28014 13957 28014 13957 0 o_result[55]
rlabel via2 28290 12971 28290 12971 0 o_result[56]
rlabel metal2 28474 13379 28474 13379 0 o_result[57]
rlabel metal1 18906 11866 18906 11866 0 o_result[58]
rlabel metal1 20884 11254 20884 11254 0 o_result[59]
rlabel metal2 19228 6732 19228 6732 0 o_result[5]
rlabel metal1 26082 11866 26082 11866 0 o_result[60]
rlabel metal2 28290 11475 28290 11475 0 o_result[61]
rlabel metal2 28290 10591 28290 10591 0 o_result[62]
rlabel metal2 23414 8925 23414 8925 0 o_result[63]
rlabel metal2 21758 5803 21758 5803 0 o_result[6]
rlabel metal2 28290 6409 28290 6409 0 o_result[7]
rlabel metal2 28290 7021 28290 7021 0 o_result[8]
rlabel metal2 28290 7633 28290 7633 0 o_result[9]
rlabel metal1 22116 7922 22116 7922 0 w_dly_sig\[10\]
rlabel metal1 21114 7956 21114 7956 0 w_dly_sig\[11\]
rlabel metal1 19412 8262 19412 8262 0 w_dly_sig\[12\]
rlabel via1 20097 8330 20097 8330 0 w_dly_sig\[13\]
rlabel metal1 19258 9418 19258 9418 0 w_dly_sig\[14\]
rlabel metal2 17342 9282 17342 9282 0 w_dly_sig\[15\]
rlabel metal1 17250 9418 17250 9418 0 w_dly_sig\[16\]
rlabel metal1 16652 9690 16652 9690 0 w_dly_sig\[17\]
rlabel metal2 15870 9622 15870 9622 0 w_dly_sig\[18\]
rlabel metal2 14674 10336 14674 10336 0 w_dly_sig\[19\]
rlabel metal1 17935 5134 17935 5134 0 w_dly_sig\[1\]
rlabel metal1 13892 10030 13892 10030 0 w_dly_sig\[20\]
rlabel metal1 14582 9350 14582 9350 0 w_dly_sig\[21\]
rlabel metal1 14122 9078 14122 9078 0 w_dly_sig\[22\]
rlabel metal1 13110 8874 13110 8874 0 w_dly_sig\[23\]
rlabel metal1 14566 8330 14566 8330 0 w_dly_sig\[24\]
rlabel metal1 14628 8262 14628 8262 0 w_dly_sig\[25\]
rlabel via1 14122 7378 14122 7378 0 w_dly_sig\[26\]
rlabel metal1 14025 6902 14025 6902 0 w_dly_sig\[27\]
rlabel metal1 12236 7446 12236 7446 0 w_dly_sig\[28\]
rlabel metal1 10810 6800 10810 6800 0 w_dly_sig\[29\]
rlabel metal1 16330 5610 16330 5610 0 w_dly_sig\[2\]
rlabel metal1 11178 6426 11178 6426 0 w_dly_sig\[30\]
rlabel viali 8974 6834 8974 6834 0 w_dly_sig\[31\]
rlabel metal2 10350 7718 10350 7718 0 w_dly_sig\[32\]
rlabel metal1 9867 7378 9867 7378 0 w_dly_sig\[33\]
rlabel metal1 8786 8364 8786 8364 0 w_dly_sig\[34\]
rlabel metal1 8280 8330 8280 8330 0 w_dly_sig\[35\]
rlabel metal1 9246 9554 9246 9554 0 w_dly_sig\[36\]
rlabel metal1 8924 9486 8924 9486 0 w_dly_sig\[37\]
rlabel metal1 8336 10098 8336 10098 0 w_dly_sig\[38\]
rlabel metal1 9158 11254 9158 11254 0 w_dly_sig\[39\]
rlabel metal2 16238 6018 16238 6018 0 w_dly_sig\[3\]
rlabel metal1 9936 10778 9936 10778 0 w_dly_sig\[40\]
rlabel metal1 11822 11594 11822 11594 0 w_dly_sig\[41\]
rlabel metal1 12926 11628 12926 11628 0 w_dly_sig\[42\]
rlabel metal1 12742 11798 12742 11798 0 w_dly_sig\[43\]
rlabel metal1 11730 12784 11730 12784 0 w_dly_sig\[44\]
rlabel metal1 10442 13158 10442 13158 0 w_dly_sig\[45\]
rlabel via1 11182 12750 11182 12750 0 w_dly_sig\[46\]
rlabel metal1 13984 13362 13984 13362 0 w_dly_sig\[47\]
rlabel metal1 11674 13838 11674 13838 0 w_dly_sig\[48\]
rlabel metal1 13156 13430 13156 13430 0 w_dly_sig\[49\]
rlabel metal1 17986 6290 17986 6290 0 w_dly_sig\[4\]
rlabel metal1 14812 14042 14812 14042 0 w_dly_sig\[50\]
rlabel metal1 15732 13362 15732 13362 0 w_dly_sig\[51\]
rlabel metal1 15916 13498 15916 13498 0 w_dly_sig\[52\]
rlabel metal1 16928 13158 16928 13158 0 w_dly_sig\[53\]
rlabel metal1 18170 13906 18170 13906 0 w_dly_sig\[54\]
rlabel metal1 19412 12954 19412 12954 0 w_dly_sig\[55\]
rlabel metal1 20424 12614 20424 12614 0 w_dly_sig\[56\]
rlabel metal2 20470 13328 20470 13328 0 w_dly_sig\[57\]
rlabel metal1 20562 12070 20562 12070 0 w_dly_sig\[58\]
rlabel metal1 18671 11594 18671 11594 0 w_dly_sig\[59\]
rlabel metal1 19591 6222 19591 6222 0 w_dly_sig\[5\]
rlabel metal1 19550 11526 19550 11526 0 w_dly_sig\[60\]
rlabel metal1 21436 11866 21436 11866 0 w_dly_sig\[61\]
rlabel metal1 21942 11016 21942 11016 0 w_dly_sig\[62\]
rlabel metal1 22172 10506 22172 10506 0 w_dly_sig\[63\]
rlabel metal2 21942 9860 21942 9860 0 w_dly_sig\[64\]
rlabel metal1 22080 9962 22080 9962 0 w_dly_sig\[65\]
rlabel metal1 18400 6766 18400 6766 0 w_dly_sig\[6\]
rlabel metal2 19826 7140 19826 7140 0 w_dly_sig\[7\]
rlabel metal2 20654 7208 20654 7208 0 w_dly_sig\[8\]
rlabel metal1 20700 7242 20700 7242 0 w_dly_sig\[9\]
rlabel metal1 16698 5100 16698 5100 0 w_dly_sig_n\[0\]
rlabel metal1 20056 7990 20056 7990 0 w_dly_sig_n\[10\]
rlabel metal1 20654 9010 20654 9010 0 w_dly_sig_n\[11\]
rlabel metal1 19780 8262 19780 8262 0 w_dly_sig_n\[12\]
rlabel metal1 19458 8976 19458 8976 0 w_dly_sig_n\[13\]
rlabel metal1 19044 9146 19044 9146 0 w_dly_sig_n\[14\]
rlabel metal1 18538 9418 18538 9418 0 w_dly_sig_n\[15\]
rlabel metal1 17664 9622 17664 9622 0 w_dly_sig_n\[16\]
rlabel metal1 15824 10098 15824 10098 0 w_dly_sig_n\[17\]
rlabel metal1 15502 10438 15502 10438 0 w_dly_sig_n\[18\]
rlabel metal1 14904 9894 14904 9894 0 w_dly_sig_n\[19\]
rlabel metal1 16330 5712 16330 5712 0 w_dly_sig_n\[1\]
rlabel metal1 14490 9690 14490 9690 0 w_dly_sig_n\[20\]
rlabel metal1 13386 9418 13386 9418 0 w_dly_sig_n\[21\]
rlabel metal1 13892 8806 13892 8806 0 w_dly_sig_n\[22\]
rlabel metal2 14306 8602 14306 8602 0 w_dly_sig_n\[23\]
rlabel metal1 13386 8058 13386 8058 0 w_dly_sig_n\[24\]
rlabel metal1 13478 7786 13478 7786 0 w_dly_sig_n\[25\]
rlabel metal1 12834 7514 12834 7514 0 w_dly_sig_n\[26\]
rlabel metal1 12098 7310 12098 7310 0 w_dly_sig_n\[27\]
rlabel metal1 12052 6698 12052 6698 0 w_dly_sig_n\[28\]
rlabel metal1 10902 6630 10902 6630 0 w_dly_sig_n\[29\]
rlabel metal1 18032 5542 18032 5542 0 w_dly_sig_n\[2\]
rlabel metal2 10442 7140 10442 7140 0 w_dly_sig_n\[30\]
rlabel metal1 8694 6970 8694 6970 0 w_dly_sig_n\[31\]
rlabel metal1 9982 7242 9982 7242 0 w_dly_sig_n\[32\]
rlabel metal1 8464 7922 8464 7922 0 w_dly_sig_n\[33\]
rlabel metal1 9292 8398 9292 8398 0 w_dly_sig_n\[34\]
rlabel metal1 8648 8806 8648 8806 0 w_dly_sig_n\[35\]
rlabel metal1 8602 9452 8602 9452 0 w_dly_sig_n\[36\]
rlabel metal1 9016 10098 9016 10098 0 w_dly_sig_n\[37\]
rlabel metal1 9844 10234 9844 10234 0 w_dly_sig_n\[38\]
rlabel metal1 9384 10506 9384 10506 0 w_dly_sig_n\[39\]
rlabel metal1 18170 5610 18170 5610 0 w_dly_sig_n\[3\]
rlabel metal1 9890 11186 9890 11186 0 w_dly_sig_n\[40\]
rlabel metal1 11040 11322 11040 11322 0 w_dly_sig_n\[41\]
rlabel metal1 12558 11628 12558 11628 0 w_dly_sig_n\[42\]
rlabel metal1 11132 13362 11132 13362 0 w_dly_sig_n\[43\]
rlabel metal1 11178 12614 11178 12614 0 w_dly_sig_n\[44\]
rlabel metal1 12006 12784 12006 12784 0 w_dly_sig_n\[45\]
rlabel metal1 11500 13498 11500 13498 0 w_dly_sig_n\[46\]
rlabel metal1 12742 13362 12742 13362 0 w_dly_sig_n\[47\]
rlabel metal2 14030 13600 14030 13600 0 w_dly_sig_n\[48\]
rlabel metal1 14444 13702 14444 13702 0 w_dly_sig_n\[49\]
rlabel metal1 18124 6222 18124 6222 0 w_dly_sig_n\[4\]
rlabel metal1 15502 13328 15502 13328 0 w_dly_sig_n\[50\]
rlabel metal1 16238 13362 16238 13362 0 w_dly_sig_n\[51\]
rlabel metal1 17572 13498 17572 13498 0 w_dly_sig_n\[52\]
rlabel metal1 18584 13838 18584 13838 0 w_dly_sig_n\[53\]
rlabel metal1 18676 12682 18676 12682 0 w_dly_sig_n\[54\]
rlabel metal1 20010 12750 20010 12750 0 w_dly_sig_n\[55\]
rlabel metal1 20700 13702 20700 13702 0 w_dly_sig_n\[56\]
rlabel metal1 20286 12138 20286 12138 0 w_dly_sig_n\[57\]
rlabel metal1 19688 11662 19688 11662 0 w_dly_sig_n\[58\]
rlabel metal1 21252 11798 21252 11798 0 w_dly_sig_n\[59\]
rlabel metal1 19090 6630 19090 6630 0 w_dly_sig_n\[5\]
rlabel metal1 21068 11186 21068 11186 0 w_dly_sig_n\[60\]
rlabel metal2 21666 10914 21666 10914 0 w_dly_sig_n\[61\]
rlabel metal1 22678 10608 22678 10608 0 w_dly_sig_n\[62\]
rlabel metal1 21620 9894 21620 9894 0 w_dly_sig_n\[63\]
rlabel metal1 21758 10166 21758 10166 0 w_dly_sig_n\[64\]
rlabel metal1 20010 6698 20010 6698 0 w_dly_sig_n\[6\]
rlabel metal1 19596 7242 19596 7242 0 w_dly_sig_n\[7\]
rlabel metal1 20700 7174 20700 7174 0 w_dly_sig_n\[8\]
rlabel metal1 21758 7412 21758 7412 0 w_dly_sig_n\[9\]
<< properties >>
string FIXED_BBOX 0 0 32000 20000
<< end >>
