* PEX produced on Fri Mar 15 07:13:16 PM CET 2024 using /foss/tools/osic-multitool/iic-pex.sh with m=1 and s=1
* NGSPICE file created from tdc.ext - technology: sky130A

.subckt tdc i_start i_stop o_result[0] o_result[14] o_result[16] o_result[19] o_result[20]
+ o_result[21] o_result[22] o_result[23] o_result[24] o_result[25] o_result[26] o_result[27]
+ o_result[28] o_result[2] o_result[32] o_result[35] o_result[37] o_result[38] o_result[3]
+ o_result[40] o_result[41] o_result[42] o_result[43] o_result[44] o_result[45] o_result[49]
+ o_result[50] o_result[51] o_result[53] o_result[54] o_result[56] o_result[57] o_result[59]
+ o_result[5] o_result[60] o_result[61] o_result[62] o_result[6] o_result[7] o_result[8]
+ o_result[46] o_result[11] o_result[48] o_result[29] o_result[34] o_result[31] o_result[13]
+ o_result[18] o_result[10] o_result[58] o_result[63] o_result[55] o_result[47] o_result[52]
+ o_result[39] o_result[36] o_result[33] o_result[30] o_result[15] o_result[12] o_result[17]
+ o_result[4] o_result[9] VPWR o_result[1] VGND
X0 VPWR a_15319_10901# o_result[55] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR clknet_3_0__leaf_i_stop a_8767_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2 a_18298_11989# a_18130_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8 o_result[32] a_11639_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_21023_11739# o_result[60] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR w_dly_sig[40] a_13262_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0672 ps=0.74 w=0.42 l=0.15
X12 a_18130_12015# a_17857_12021# a_18045_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X13 VGND a_14894_10901# a_14852_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14 VGND a_20138_7637# a_20096_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X16 VGND a_13295_11989# a_13253_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X17 VGND a_14599_9839# a_14767_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 w_dly_sig_n[11] w_dly_sig[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_21633_7663# w_dly_sig[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X26 VGND a_17159_8725# o_result[42] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 w_dly_sig_n[0] net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 VPWR a_9389_11445# clknet_3_2__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X31 VGND a_18539_10901# a_18497_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X32 VGND w_dly_sig_n[41] w_dly_sig[42] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 clknet_0_i_stop a_16197_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X34 a_11694_9661# a_11447_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X35 w_dly_sig_n[37] w_dly_sig[37] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X36 clknet_3_5__leaf_i_stop a_21822_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X37 a_19329_6581# a_19163_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X39 a_20295_10927# a_19513_10933# a_20211_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X40 VGND w_dly_sig[40] w_dly_sig_n[40] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X44 VGND w_dly_sig[54] w_dly_sig_n[54] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X45 a_15649_6397# a_15115_6031# a_15554_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X46 a_15036_9129# a_14637_8757# a_14910_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X48 a_8946_8207# a_8559_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X51 VPWR a_14691_12015# a_14859_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X54 VGND a_21822_8207# clknet_3_5__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X57 VPWR a_9111_13335# o_result[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X59 clknet_3_3__leaf_i_stop a_14449_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X61 a_14174_6575# a_13901_6581# a_14089_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X62 VGND clknet_3_4__leaf_i_stop a_17967_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X64 a_17359_10749# a_16495_10383# a_17102_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X65 a_14637_8757# a_14471_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X67 VPWR clknet_3_7__leaf_i_stop a_19991_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X68 a_12023_10927# a_11159_10933# a_11766_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X70 VGND a_14817_7093# clknet_3_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X73 VGND a_16197_9813# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X74 clknet_3_4__leaf_i_stop a_16854_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X75 VPWR a_12835_6549# o_result[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X77 VPWR a_9665_7093# clknet_3_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X78 o_result[45] a_20566_10636# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X81 VGND w_dly_sig_n[28] w_dly_sig[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X82 a_12889_10933# a_12723_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X83 a_11693_10927# a_11159_10933# a_11598_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X86 VPWR clknet_3_1__leaf_i_stop a_13735_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X88 o_result[24] a_8559_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X89 VGND a_17010_7637# a_16968_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X90 VPWR w_dly_sig_n[5] w_dly_sig[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X91 VPWR w_dly_sig[29] w_dly_sig_n[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X92 VGND a_16854_8207# clknet_3_4__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X96 VGND a_11639_12827# o_result[32] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X98 a_16941_6575# w_dly_sig[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X100 a_19421_12021# a_19255_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X101 VGND clknet_0_i_stop a_16749_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X102 a_8743_6005# a_8911_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X103 w_dly_sig[53] w_dly_sig_n[52] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X104 a_11411_7895# a_11579_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X105 clknet_0_i_stop a_16197_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X110 w_dly_sig[4] w_dly_sig_n[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X113 VGND clknet_3_7__leaf_i_stop a_19623_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X115 a_20855_11837# a_20157_11471# a_20598_11583# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X116 a_16661_10383# a_16495_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X120 a_15036_8041# a_14637_7669# a_14910_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X122 VGND w_dly_sig_n[36] w_dly_sig[37] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X124 clknet_3_0__leaf_i_stop a_9665_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X125 w_dly_sig_n[55] w_dly_sig[55] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X127 a_10117_13481# a_9570_13225# a_9770_13380# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X128 a_17102_10495# a_16934_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X129 a_12157_6575# w_dly_sig[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X130 o_result[61] a_20655_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X131 a_17861_10927# w_dly_sig[54] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X132 a_13254_8751# a_12981_8757# a_13169_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X135 clknet_3_7__leaf_i_stop a_21822_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X136 VPWR a_11766_10901# a_11693_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X137 VPWR a_22679_10651# o_result[50] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X138 VPWR w_dly_sig_n[61] w_dly_sig[62] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X143 w_dly_sig[30] w_dly_sig_n[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X145 VGND a_12191_10901# a_12149_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X148 a_11447_9295# a_11318_9569# a_11027_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X152 w_dly_sig_n[44] w_dly_sig[44] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X154 a_9647_10357# a_9938_10657# a_9889_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X155 a_11865_9295# a_11318_9569# a_11518_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X156 a_16293_8757# a_16127_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X158 VGND a_10859_9269# o_result[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X160 a_22580_10217# a_22181_9845# a_22454_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X161 a_20571_13103# a_19789_13109# a_20487_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X164 w_dly_sig[52] w_dly_sig_n[51] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X165 w_dly_sig_n[51] w_dly_sig[51] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X166 VGND a_14767_9813# o_result[40] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X168 w_dly_sig[14] w_dly_sig_n[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X170 VPWR w_dly_sig[62] w_dly_sig_n[62] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X171 VPWR clknet_3_0__leaf_i_stop a_11251_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X178 o_result[14] a_17619_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X179 w_dly_sig_n[21] w_dly_sig[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X180 a_18406_7663# a_18133_7669# a_18321_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X181 VPWR a_19735_8475# o_result[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X184 VGND w_dly_sig_n[20] w_dly_sig[21] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X185 VPWR a_16975_12827# a_16891_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X186 VPWR clknet_3_6__leaf_i_stop a_19255_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X187 o_result[28] a_8927_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X188 VPWR a_14342_6549# a_14269_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X189 a_12797_12015# a_12263_12021# a_12702_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X192 VPWR w_dly_sig[47] w_dly_sig_n[47] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X195 VPWR w_dly_sig_n[34] w_dly_sig[35] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X200 o_result[20] a_11363_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X204 o_result[39] a_12050_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.185 ps=1.87 w=0.65 l=0.15
X205 VPWR w_dly_sig[11] w_dly_sig_n[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X208 a_9195_6005# clknet_3_0__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X209 VGND a_13330_10901# a_13288_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X211 VPWR w_dly_sig[23] w_dly_sig_n[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X214 clknet_3_2__leaf_i_stop a_9389_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X215 a_22086_10749# a_21647_10383# a_22001_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X216 VPWR a_12050_9813# o_result[39] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X217 clknet_3_6__leaf_i_stop a_16749_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X219 a_20153_6953# a_19163_6581# a_20027_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X222 VPWR a_9931_10357# a_9938_10657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X223 VPWR a_22311_8725# o_result[47] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X224 o_result[52] a_20379_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X226 VGND clknet_3_4__leaf_i_stop a_16403_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X227 w_dly_sig[15] w_dly_sig_n[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X229 VGND a_15319_10901# o_result[55] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X233 VPWR a_20211_10927# a_20379_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X234 o_result[26] a_9203_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X235 VPWR a_13422_8725# a_13349_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X238 VGND a_14817_7093# clknet_3_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X239 a_9379_11145# clknet_3_2__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X240 VGND w_dly_sig[27] w_dly_sig_n[27] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X241 a_22089_6031# a_21923_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X242 VPWR a_11471_12925# a_11639_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X243 o_result[60] a_21023_11739# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X245 w_dly_sig_n[19] w_dly_sig[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X246 VPWR w_dly_sig_n[9] w_dly_sig[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X247 a_13671_10927# a_12889_10933# a_13587_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X249 VPWR w_dly_sig[36] w_dly_sig_n[36] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X251 w_dly_sig[23] w_dly_sig_n[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X252 w_dly_sig[26] w_dly_sig_n[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X254 a_9758_7663# a_9485_7669# a_9673_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X257 VGND a_14817_7093# clknet_3_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X258 VPWR a_14817_7093# clknet_3_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X261 w_dly_sig_n[59] w_dly_sig[59] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X262 VGND w_dly_sig[39] w_dly_sig_n[39] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X263 VGND w_dly_sig[45] w_dly_sig_n[45] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X266 VGND clknet_0_i_stop a_9665_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X268 a_22270_13103# a_21831_13109# a_22185_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X269 a_10209_10217# a_9655_10057# a_9862_10116# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X270 VPWR w_dly_sig[8] w_dly_sig_n[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X271 a_16749_11445# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X272 a_18681_9129# a_17691_8757# a_18555_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X275 VPWR a_13295_11989# o_result[36] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X276 clknet_3_7__leaf_i_stop a_21822_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X278 a_18045_12015# w_dly_sig[59] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X279 a_11724_11471# a_11325_11471# a_11598_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X281 VGND w_dly_sig_n[63] w_dly_sig[64] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X282 VGND a_13295_11989# o_result[36] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X283 a_20525_11837# a_19991_11471# a_20430_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X286 VPWR a_14875_12925# a_15043_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X287 a_14434_11989# a_14266_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X290 clknet_3_3__leaf_i_stop a_14449_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X293 VPWR a_18574_7637# a_18501_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X294 clknet_3_3__leaf_i_stop a_14449_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X298 a_12107_11837# a_11325_11471# a_12023_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X301 VGND a_22587_10901# a_22545_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X302 w_dly_sig[13] w_dly_sig_n[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X303 a_22913_7119# a_21923_7119# a_22787_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X305 a_21633_8751# w_dly_sig[48] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X306 w_dly_sig[29] w_dly_sig_n[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X307 VGND w_dly_sig[52] w_dly_sig_n[52] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X309 VGND a_16854_8207# clknet_3_4__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X310 VPWR w_dly_sig[30] w_dly_sig_n[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X311 VGND a_16749_11445# clknet_3_6__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X312 a_20521_8041# a_19531_7669# a_20395_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X313 VPWR clknet_3_7__leaf_i_stop a_22199_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X315 VGND clknet_0_i_stop a_9389_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X321 w_dly_sig_n[13] w_dly_sig[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X324 VGND clknet_3_0__leaf_i_stop a_11251_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X328 VPWR clknet_0_i_stop a_14817_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X329 a_13427_7881# clknet_3_1__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X332 VPWR a_18723_11989# a_18639_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X333 VPWR a_20598_11583# a_20525_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X334 a_22365_9295# a_22199_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 a_8969_8573# a_8559_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X336 a_18501_7663# a_17967_7669# a_18406_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X338 VGND w_dly_sig[17] w_dly_sig_n[17] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X339 clknet_3_0__leaf_i_stop a_9665_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X341 VGND clknet_3_6__leaf_i_stop a_16495_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X346 VPWR a_15503_7637# o_result[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X348 w_dly_sig[37] w_dly_sig_n[36] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X349 w_dly_sig_n[18] w_dly_sig[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X350 a_22806_11989# a_22638_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X351 VPWR a_20487_13103# a_20655_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X352 a_14775_12015# a_13993_12021# a_14691_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X353 a_18072_11305# a_17673_10933# a_17946_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X355 VGND a_20487_13103# a_20655_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X356 VPWR w_dly_sig_n[31] w_dly_sig[32] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X359 clknet_0_i_stop a_16197_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X362 a_22913_6031# a_21923_6031# a_22787_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X364 a_9203_10071# a_9371_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X367 VPWR a_9926_7637# a_9853_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X368 VPWR w_dly_sig[34] w_dly_sig_n[34] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X370 a_17393_8041# a_16403_7669# a_17267_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X371 a_22530_7231# a_22362_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X374 a_9590_10205# a_9203_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X377 a_20487_13103# a_19623_13109# a_20230_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X379 a_14825_7663# w_dly_sig[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X381 VPWR a_11639_12827# o_result[32] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X382 VGND a_9126_9269# a_9055_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X387 o_result[1] a_12283_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X389 a_20157_13103# a_19623_13109# a_20062_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X390 VGND a_12191_10901# o_result[38] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X393 a_9665_7093# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X397 w_dly_sig[55] w_dly_sig_n[54] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X398 w_dly_sig_n[28] w_dly_sig[28] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X399 a_19885_10383# w_dly_sig[46] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X400 VPWR a_18723_8725# o_result[43] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X403 a_12828_12393# a_12429_12021# a_12702_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X404 clknet_3_5__leaf_i_stop a_21822_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X405 w_dly_sig_n[15] w_dly_sig[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X407 o_result[38] a_12191_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X408 a_19786_10927# a_19513_10933# a_19701_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X409 a_15001_12559# a_14011_12559# a_14875_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X412 VPWR a_12667_6575# a_12835_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X413 VPWR w_dly_sig[44] w_dly_sig_n[44] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X415 a_22001_10383# w_dly_sig[51] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X418 VPWR w_dly_sig_n[14] w_dly_sig[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X420 a_14817_7093# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X422 VPWR w_dly_sig[27] w_dly_sig_n[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X423 a_9853_7663# a_9319_7669# a_9758_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X426 VPWR a_16854_8207# clknet_3_4__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X428 VPWR a_22695_13103# a_22863_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X429 VGND a_22695_13103# a_22863_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X434 a_19697_10383# a_19531_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X435 a_19310_8319# a_19142_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X437 o_result[21] a_8743_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X440 a_20345_11471# w_dly_sig[61] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X442 clknet_3_4__leaf_i_stop a_16854_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X446 w_dly_sig[63] w_dly_sig_n[62] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X447 clknet_3_2__leaf_i_stop a_9389_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X448 w_dly_sig_n[38] w_dly_sig[38] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X449 VGND w_dly_sig[6] w_dly_sig_n[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X450 VPWR w_dly_sig_n[22] w_dly_sig[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X452 a_22530_6143# a_22362_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X453 a_12107_10927# a_11325_10933# a_12023_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X454 VPWR a_13587_10927# a_13755_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X455 a_21813_10383# a_21647_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X456 VPWR a_9862_10116# a_9791_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X457 VGND w_dly_sig[53] w_dly_sig_n[53] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X458 VPWR a_16197_9813# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X460 w_dly_sig_n[58] w_dly_sig[58] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X461 a_14449_11445# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X462 a_18045_8751# w_dly_sig[44] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X464 a_14959_12925# a_14177_12559# a_14875_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X466 VGND a_12835_6549# o_result[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X468 VGND clknet_3_4__leaf_i_stop a_16587_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X469 a_12751_6575# a_11969_6581# a_12667_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X470 VGND w_dly_sig_n[8] w_dly_sig[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X473 a_10770_6397# a_10331_6031# a_10685_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X475 a_16481_9295# w_dly_sig[42] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X476 VGND a_9665_7093# clknet_3_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X478 VGND w_dly_sig_n[52] w_dly_sig[53] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X479 VPWR w_dly_sig[2] w_dly_sig_n[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X480 o_result[18] a_11411_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X482 VPWR a_14449_11445# clknet_3_3__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X484 a_13783_8029# a_13563_8041# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X486 a_8727_8181# a_9018_8481# a_8969_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X488 VGND clknet_3_1__leaf_i_stop a_15115_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X489 VPWR w_dly_sig_n[62] w_dly_sig[63] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X491 a_11046_12925# a_10607_12559# a_10961_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X493 VPWR w_dly_sig[1] a_11865_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X494 a_22269_9129# a_21279_8757# a_22143_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X497 a_13587_10927# a_12723_10933# a_13330_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X498 w_dly_sig_n[41] w_dly_sig[41] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X499 VGND a_9218_8181# a_9147_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X501 a_13257_10927# a_12723_10933# a_13162_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X502 a_11863_7881# clknet_3_1__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X504 VPWR a_23047_9813# a_22963_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X505 w_dly_sig_n[43] w_dly_sig[43] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X508 VPWR a_20655_13077# o_result[61] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X510 VGND a_20655_13077# o_result[61] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X514 a_21718_7663# a_21445_7669# a_21633_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X515 VGND a_22311_7637# o_result[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X516 a_12610_13103# a_12337_13109# a_12525_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X517 a_18681_12393# a_17691_12021# a_18555_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X520 VPWR a_17159_9563# o_result[41] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X521 o_result[36] a_13295_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X522 a_11195_6397# a_10331_6031# a_10938_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X523 a_9371_10071# a_9655_10057# a_9590_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X524 VPWR a_9665_7093# clknet_3_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X525 a_9011_8181# clknet_3_0__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X530 VGND a_14342_6549# a_14300_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X531 VGND w_dly_sig[32] w_dly_sig_n[32] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X532 a_10896_6031# a_10497_6031# a_10770_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X534 VPWR a_17159_11989# a_17075_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X535 VPWR a_20566_10636# a_20479_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X537 VGND clknet_0_i_stop a_16854_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X539 a_19694_12015# a_19255_12021# a_19609_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X540 w_dly_sig[51] w_dly_sig_n[50] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X544 a_9643_12381# a_9423_12393# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X547 clknet_0_i_stop a_16197_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X548 VGND a_22622_9813# a_22580_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X549 a_21886_8725# a_21718_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X551 a_22269_8041# a_21279_7669# a_22143_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X554 w_dly_sig[49] w_dly_sig_n[48] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X556 a_17673_10933# a_17507_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X557 w_dly_sig_n[46] w_dly_sig[46] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X558 clknet_3_0__leaf_i_stop a_9665_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X564 VGND a_12070_7940# a_11999_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X568 VGND w_dly_sig_n[11] w_dly_sig[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X569 a_11325_11471# a_11159_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X571 VGND a_22162_10901# a_22120_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X572 o_result[51] a_22587_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X577 a_22277_7119# w_dly_sig[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X579 a_11046_12925# a_10773_12559# a_10961_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X581 VGND a_10938_6143# a_10896_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X583 clknet_3_1__leaf_i_stop a_14817_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X584 a_10309_8041# a_9319_7669# a_10183_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X585 o_result[15] a_16147_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X587 a_16297_12559# w_dly_sig[58] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X589 a_8919_9269# clknet_3_0__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X590 VPWR a_21822_11471# clknet_3_7__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X592 w_dly_sig[48] w_dly_sig_n[47] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X593 a_12975_7895# a_13143_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X596 w_dly_sig[32] w_dly_sig_n[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X597 VPWR a_13755_10901# o_result[37] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X598 VGND a_17159_9563# o_result[41] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X599 VGND clknet_3_0__leaf_i_stop a_8767_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X602 VPWR a_22143_8751# a_22311_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X607 a_22511_10749# a_21813_10383# a_22254_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X610 a_22503_10927# a_21721_10933# a_22419_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X616 a_16481_8751# w_dly_sig[43] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X618 VPWR a_21886_7637# a_21813_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X619 a_12337_6575# a_11803_6581# a_12242_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X622 a_8559_8181# a_8727_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X624 a_20188_13481# a_19789_13109# a_20062_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X625 VGND a_15043_12827# o_result[34] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X626 VPWR w_dly_sig[22] w_dly_sig_n[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X627 VPWR a_11363_6299# a_11279_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X629 a_16749_11445# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X630 a_9389_11445# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X631 clknet_3_7__leaf_i_stop a_21822_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X632 o_result[55] a_15319_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X634 a_10938_6143# a_10770_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X636 o_result[38] a_12191_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X637 VGND a_14449_11445# clknet_3_3__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X638 VPWR clknet_3_4__leaf_i_stop a_17691_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X640 a_17857_12021# a_17691_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X641 VPWR a_17619_6549# a_17535_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X643 VPWR w_dly_sig[13] w_dly_sig_n[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X645 a_14089_6575# w_dly_sig[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X649 VGND net1 a_10975_8759# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X650 clknet_3_5__leaf_i_stop a_21822_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X651 clknet_3_5__leaf_i_stop a_21822_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X654 w_dly_sig[44] w_dly_sig_n[43] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X659 VPWR w_dly_sig[5] w_dly_sig_n[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X660 VGND clknet_3_5__leaf_i_stop a_19531_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X661 a_19786_10927# a_19347_10933# a_19701_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X662 clknet_3_4__leaf_i_stop a_16854_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X663 VGND clknet_3_1__leaf_i_stop a_13735_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X664 a_21813_7663# a_21279_7669# a_21718_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X665 a_16933_12559# a_15943_12559# a_16807_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X666 a_15235_10927# a_14453_10933# a_15151_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X667 o_result[12] a_20195_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X668 VPWR a_13634_7940# a_13563_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X673 a_15722_6143# a_15554_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X674 a_11999_8041# a_11863_7881# a_11579_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X675 VGND a_13587_10927# a_13755_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X678 VPWR a_16197_9813# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X679 a_9011_8181# clknet_3_0__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X681 o_result[31] a_9111_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X682 clknet_3_3__leaf_i_stop a_14449_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X684 VPWR w_dly_sig[57] w_dly_sig_n[57] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X685 VPWR clknet_3_7__leaf_i_stop a_21647_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X687 a_10961_12559# w_dly_sig[33] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X689 VGND w_dly_sig_n[57] w_dly_sig[58] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X691 VGND a_18114_10901# a_18072_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X693 VPWR a_14859_11989# o_result[35] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X696 a_16991_12015# a_16293_12021# a_16734_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X697 VGND a_14859_11989# o_result[35] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X698 a_17117_12393# a_16127_12021# a_16991_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X699 a_16734_11989# a_16566_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X700 a_10685_6031# w_dly_sig[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X702 VPWR a_14817_7093# clknet_3_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X705 a_12736_13481# a_12337_13109# a_12610_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X709 a_16566_12015# a_16293_12021# a_16481_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X711 a_18574_7637# a_18406_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X712 w_dly_sig_n[54] w_dly_sig[54] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X716 a_13901_9845# a_13735_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X721 VGND a_15503_7637# o_result[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X723 a_14599_6575# a_13735_6581# a_14342_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X725 clknet_3_2__leaf_i_stop a_9389_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X728 VPWR clknet_3_5__leaf_i_stop a_21279_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X731 VPWR w_dly_sig_n[4] w_dly_sig[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X734 a_20076_10383# a_19697_10383# a_19979_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X735 VPWR clknet_3_0__leaf_i_stop a_10331_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X737 a_15078_8725# a_14910_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X738 VPWR w_dly_sig[12] w_dly_sig_n[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X740 a_19954_9407# a_19786_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X742 a_20111_6575# a_19329_6581# a_20027_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X744 a_11411_7895# a_11579_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X745 w_dly_sig[62] w_dly_sig_n[61] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X747 w_dly_sig[38] w_dly_sig_n[37] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X748 clknet_0_i_stop a_16197_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X749 a_13679_8751# a_12981_8757# a_13422_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X754 VPWR a_9665_7093# clknet_3_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X756 VPWR a_23231_11989# o_result[63] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X758 a_9121_6575# w_dly_sig[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X760 VPWR clknet_0_i_stop a_21822_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X761 w_dly_sig_n[46] w_dly_sig[46] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X763 VGND a_9926_7637# a_9884_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X765 o_result[44] a_19091_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X769 a_15078_8725# a_14910_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X770 a_22511_10749# a_21647_10383# a_22254_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X771 w_dly_sig[41] w_dly_sig_n[40] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X772 VGND w_dly_sig_n[38] w_dly_sig[39] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X774 a_20395_10749# a_19697_10383# a_20138_10519# VGND sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X776 a_14089_9839# w_dly_sig[41] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X778 a_22181_10749# a_21647_10383# a_22086_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X779 VGND a_22955_7387# o_result[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X780 w_dly_sig_n[26] w_dly_sig[26] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X782 VGND a_20563_7637# a_20521_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X784 VGND a_9389_11445# clknet_3_2__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X785 VGND clknet_3_6__leaf_i_stop a_17507_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X786 a_12821_10217# a_12688_10057# a_12400_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X787 a_9055_9295# a_8919_9269# a_8635_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X788 a_13679_8751# a_12815_8757# a_13422_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X789 a_17117_9129# a_16127_8757# a_16991_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X790 VGND w_dly_sig_n[16] w_dly_sig[17] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X791 o_result[51] a_22587_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X792 a_9245_12015# a_8835_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X794 VGND a_12667_6575# a_12835_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X797 VPWR clknet_3_5__leaf_i_stop a_21279_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X798 clknet_0_i_stop a_16197_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X799 VPWR a_22419_10927# a_22587_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X800 a_16566_9661# a_16293_9295# a_16481_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X801 a_22362_6397# a_22089_6031# a_22277_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X802 a_18321_7663# w_dly_sig[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X805 a_12337_13109# a_12171_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X806 VPWR a_16749_11445# clknet_3_6__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X807 o_result[8] a_22311_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X809 VGND a_13755_10901# o_result[37] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X811 a_14894_10901# a_14726_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X812 w_dly_sig[7] w_dly_sig_n[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X814 o_result[37] a_13755_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X815 VPWR a_15335_8751# a_15503_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X817 w_dly_sig_n[60] w_dly_sig[60] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X818 w_dly_sig_n[24] w_dly_sig[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X820 a_20524_10383# a_19531_10383# a_20395_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X823 VPWR a_22254_10495# a_22181_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X825 VGND a_9402_6005# a_9331_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X826 VPWR a_17010_7637# a_16937_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X827 a_22419_10927# a_21555_10933# a_22162_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X829 VGND w_dly_sig[31] w_dly_sig_n[31] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X830 VGND a_22955_6299# o_result[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X831 VPWR a_14767_6549# a_14683_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X832 VGND a_17159_11989# a_17117_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X833 o_result[23] a_10351_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X834 a_22089_10927# a_21555_10933# a_21994_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X835 VPWR a_16991_9661# a_17159_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X836 w_dly_sig_n[1] w_dly_sig[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X837 clknet_3_6__leaf_i_stop a_16749_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X839 a_21822_11471# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X840 VGND a_17435_7637# a_17393_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X841 o_result[55] a_15319_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X842 a_19701_10927# w_dly_sig[53] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X844 a_9389_11445# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X846 w_dly_sig_n[17] w_dly_sig[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X847 a_22227_7663# a_21445_7669# a_22143_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X848 o_result[34] a_15043_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X849 VGND a_14449_11445# clknet_3_3__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X850 VGND w_dly_sig[19] a_12417_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X851 VGND a_14449_11445# clknet_3_3__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X852 VPWR a_15151_10927# a_15319_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X854 a_9153_6397# a_8743_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X855 clknet_3_0__leaf_i_stop a_9665_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X856 w_dly_sig_n[27] w_dly_sig[27] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X857 VPWR a_9379_11145# a_9386_11049# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X860 a_18831_7663# a_17967_7669# a_18574_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X862 VPWR a_20379_10901# o_result[52] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X864 VPWR w_dly_sig[18] a_13981_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X868 a_16382_12925# a_15943_12559# a_16297_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X869 VPWR a_11639_12827# a_11555_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X870 w_dly_sig[31] w_dly_sig_n[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X871 VPWR a_23231_11989# a_23147_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X873 w_dly_sig[3] w_dly_sig_n[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X874 a_15005_7663# a_14471_7669# a_14910_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X875 VPWR w_dly_sig_n[43] w_dly_sig[44] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X878 a_9314_11293# a_8927_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X879 VPWR a_16197_9813# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X881 a_16569_7669# a_16403_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X882 a_9699_13481# a_9563_13321# a_9279_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X883 VPWR w_dly_sig[29] a_9933_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X884 a_9673_7663# w_dly_sig[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X885 a_19602_6575# a_19329_6581# a_19517_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X886 w_dly_sig_n[25] w_dly_sig[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X887 VGND w_dly_sig[9] w_dly_sig_n[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X893 VPWR clknet_3_6__leaf_i_stop a_18059_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X894 VPWR a_13847_8725# a_13763_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X895 clknet_3_3__leaf_i_stop a_14449_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X897 VPWR a_12050_9813# o_result[39] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X901 VGND clknet_0_i_stop a_14817_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X902 VGND a_9665_7093# clknet_3_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X904 a_20345_11471# w_dly_sig[61] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X905 a_22871_7485# a_22089_7119# a_22787_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X906 w_dly_sig[8] w_dly_sig_n[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X907 VPWR clknet_3_7__leaf_i_stop a_21831_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X908 a_9287_12233# clknet_3_2__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X909 w_dly_sig[58] w_dly_sig_n[57] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X910 VPWR a_16734_9407# a_16661_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X911 VPWR a_22530_6143# a_22457_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X914 VPWR a_15043_12827# a_14959_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X917 VPWR a_15043_12827# o_result[34] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X920 VGND a_9111_13335# o_result[31] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X921 VPWR w_dly_sig_n[26] w_dly_sig[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X923 a_16197_9813# i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X928 a_20157_11471# a_19991_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X931 w_dly_sig[10] w_dly_sig_n[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X933 VPWR a_12892_10116# a_12821_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X935 a_16566_8751# a_16293_8757# a_16481_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X936 VPWR a_18999_7637# a_18915_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X938 VGND a_12283_8475# a_12241_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X940 a_22695_13103# a_21831_13109# a_22438_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X941 a_18371_10927# a_17507_10933# a_18114_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X942 a_16661_9661# a_16127_9295# a_16566_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X943 VPWR clknet_3_1__leaf_i_stop a_14471_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X946 a_19142_8573# a_18869_8207# a_19057_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X948 a_22365_13103# a_21831_13109# a_22270_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X951 a_18041_10927# a_17507_10933# a_17946_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X953 a_8743_6005# a_8911_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X954 a_9933_11305# a_9386_11049# a_9586_11204# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X955 VPWR a_14767_9813# o_result[40] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X957 a_19789_13109# a_19623_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X959 a_18225_9845# a_18059_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X960 a_9331_6031# a_9195_6005# a_8911_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X961 VPWR w_dly_sig[35] w_dly_sig_n[35] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X962 VPWR a_9586_11204# a_9515_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X963 w_dly_sig[18] w_dly_sig_n[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X964 w_dly_sig_n[52] w_dly_sig[52] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X965 a_12219_8029# a_11999_8041# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X968 VPWR w_dly_sig[55] w_dly_sig_n[55] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X972 a_19609_12015# w_dly_sig[60] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X974 w_dly_sig_n[7] w_dly_sig[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X975 VGND w_dly_sig[4] w_dly_sig_n[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X979 w_dly_sig_n[39] w_dly_sig[39] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X980 VPWR a_20395_10749# a_20566_10636# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X981 clknet_3_6__leaf_i_stop a_16749_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X982 a_18666_9813# a_18498_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X983 VPWR a_20379_9563# a_20295_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X985 VPWR a_21822_8207# clknet_3_5__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X987 VPWR a_19770_6549# a_19697_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X989 a_14725_10217# a_13735_9845# a_14599_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X990 VPWR w_dly_sig_n[40] w_dly_sig[41] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X991 VGND a_18723_8725# o_result[43] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X994 VGND a_16854_8207# clknet_3_4__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X996 a_14875_12925# a_14177_12559# a_14618_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X997 VGND a_9389_11445# clknet_3_2__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1000 VPWR a_22438_13077# a_22365_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1001 VPWR a_18114_10901# a_18041_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1003 a_9563_13321# clknet_3_2__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1005 VPWR w_dly_sig_n[0] w_dly_sig[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1007 VGND a_22419_10927# a_22587_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1008 a_14089_9839# w_dly_sig[41] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1009 a_15554_6397# a_15281_6031# a_15469_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1010 w_dly_sig[46] w_dly_sig_n[45] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1011 VPWR a_12023_10927# a_12191_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1012 o_result[5] a_17435_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1013 VPWR a_16749_11445# clknet_3_6__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1014 VGND clknet_3_7__leaf_i_stop a_19531_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1015 a_19513_9295# a_19347_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1017 clknet_3_1__leaf_i_stop a_14817_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1019 VGND w_dly_sig[3] w_dly_sig_n[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1022 a_12793_6953# a_11803_6581# a_12667_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1023 VPWR a_9389_11445# clknet_3_2__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1024 VGND w_dly_sig_n[51] w_dly_sig[52] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1025 VPWR w_dly_sig[51] w_dly_sig_n[51] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1027 VPWR w_dly_sig_n[35] w_dly_sig[36] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1030 clknet_3_3__leaf_i_stop a_14449_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1031 w_dly_sig_n[48] w_dly_sig[48] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1032 a_12115_8573# a_11251_8207# a_11858_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1034 VGND w_dly_sig[61] w_dly_sig_n[61] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1038 VGND clknet_3_7__leaf_i_stop a_21555_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1039 VGND w_dly_sig[38] w_dly_sig_n[38] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1040 clknet_3_1__leaf_i_stop a_14817_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1046 VGND w_dly_sig_n[58] w_dly_sig[59] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1047 a_10287_10383# a_10067_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1048 a_12050_9813# a_12400_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.162 ps=1.33 w=1 l=0.15
X1050 VPWR w_dly_sig_n[1] w_dly_sig[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1051 VPWR a_16734_8725# a_16661_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1053 VPWR a_22863_13077# o_result[62] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1054 VGND a_22863_13077# o_result[62] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1056 VGND a_16147_6299# o_result[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1057 a_22457_7485# a_21923_7119# a_22362_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1059 w_dly_sig[25] w_dly_sig_n[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1060 w_dly_sig_n[10] w_dly_sig[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1064 clknet_3_6__leaf_i_stop a_16749_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1066 a_12975_7895# a_13143_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1067 a_21822_11471# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1068 w_dly_sig[47] w_dly_sig_n[46] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1069 VPWR a_19310_8319# a_19237_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1071 clknet_3_2__leaf_i_stop a_9389_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1072 VGND a_12050_9813# o_result[39] VGND sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X1073 a_15419_7663# a_14637_7669# a_15335_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1077 VPWR a_17194_6549# a_17121_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1078 VGND a_14449_11445# clknet_3_3__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1080 VGND a_14449_11445# clknet_3_3__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1081 a_12688_10057# clknet_3_3__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1083 w_dly_sig[12] w_dly_sig_n[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1086 w_dly_sig[22] w_dly_sig_n[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1087 clknet_3_5__leaf_i_stop a_21822_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1089 a_11214_12671# a_11046_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1090 VPWR w_dly_sig_n[27] w_dly_sig[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1093 a_9931_10357# clknet_3_2__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1094 a_9206_6575# a_8933_6581# a_9121_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1095 VGND a_20379_10901# o_result[52] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1098 VPWR a_23047_9813# o_result[49] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1099 a_22637_10383# a_21647_10383# a_22511_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1102 a_9841_12393# a_9294_12137# a_9494_12292# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1104 a_14450_12925# a_14177_12559# a_14365_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1105 a_18555_12015# a_17857_12021# a_18298_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1106 clknet_3_0__leaf_i_stop a_9665_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1108 a_16661_8751# a_16127_8757# a_16566_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1114 VPWR a_9494_12292# a_9423_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1115 a_21822_8207# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1117 VGND w_dly_sig[40] a_13262_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1119 VGND a_22787_7485# a_22955_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1123 clknet_3_4__leaf_i_stop a_16854_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1127 a_17121_6575# a_16587_6581# a_17026_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1128 VPWR a_13127_12015# a_13295_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1129 a_20072_10749# a_19531_10383# a_19979_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X1130 VGND a_13127_12015# a_13295_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1131 a_22212_10383# a_21813_10383# a_22086_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1133 VPWR a_20287_11989# a_20203_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1135 VPWR a_15722_6143# a_15649_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1138 VPWR a_14817_7093# clknet_3_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1139 VGND a_18371_10927# a_18539_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1140 VPWR clknet_3_4__leaf_i_stop a_16127_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1141 a_16854_8207# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1142 VGND a_14767_9813# a_14725_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1143 VGND a_21886_8725# a_21844_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1145 a_22369_9839# w_dly_sig[50] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1147 a_16481_12015# w_dly_sig[57] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1148 clknet_0_i_stop a_16197_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1149 a_17075_9661# a_16293_9295# a_16991_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1151 VPWR a_12283_8475# a_12199_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1153 w_dly_sig[34] w_dly_sig_n[33] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1154 o_result[34] a_15043_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1156 a_18923_9839# a_18059_9845# a_18666_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1157 a_16197_9813# i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1161 w_dly_sig[43] w_dly_sig_n[42] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1163 VPWR w_dly_sig[63] w_dly_sig_n[63] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1165 o_result[20] a_11363_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1168 o_result[48] a_23231_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1171 VGND a_22787_6397# a_22955_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1173 VGND clknet_3_2__leaf_i_stop a_11159_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1176 a_22396_13481# a_21997_13109# a_22270_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1178 a_22365_12021# a_22199_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1179 w_dly_sig[50] w_dly_sig_n[49] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1180 a_20230_13077# a_20062_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1182 o_result[8] a_22311_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1183 VGND a_11766_11583# a_11724_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1189 VGND a_22143_8751# a_22311_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1191 VPWR a_14449_11445# clknet_3_3__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1194 a_20430_11837# a_19991_11471# a_20345_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1195 VPWR a_9374_6549# a_9301_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1197 VGND w_dly_sig[64] w_dly_sig_n[64] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1200 VPWR a_21822_11471# clknet_3_7__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1204 clknet_3_6__leaf_i_stop a_16749_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1205 clknet_3_6__leaf_i_stop a_16749_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1207 o_result[61] a_20655_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1210 o_result[23] a_10351_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1211 VPWR w_dly_sig_n[41] w_dly_sig[42] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1212 VPWR w_dly_sig_n[10] w_dly_sig[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1215 a_19770_6549# a_19602_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1217 VGND a_9389_11445# clknet_3_2__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1227 VGND w_dly_sig_n[55] w_dly_sig[56] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1228 VPWR a_9563_13321# a_9570_13225# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1229 VGND a_12023_10927# a_12191_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1231 a_14817_7093# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1233 VPWR a_12191_11739# a_12107_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1234 clknet_3_7__leaf_i_stop a_21822_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1236 a_9301_6575# a_8767_6581# a_9206_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1237 o_result[48] a_23231_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1238 w_dly_sig[6] w_dly_sig_n[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1240 a_14181_12015# w_dly_sig[36] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1241 VPWR a_9389_11445# clknet_3_2__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1245 clknet_3_3__leaf_i_stop a_14449_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1246 a_21718_6575# a_21279_6581# a_21633_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1247 w_dly_sig[20] w_dly_sig_n[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1249 w_dly_sig[33] w_dly_sig_n[32] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1252 VPWR a_19862_11989# a_19789_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1253 a_21633_8751# w_dly_sig[48] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1260 a_12778_13077# a_12610_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1261 w_dly_sig_n[61] w_dly_sig[61] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1262 VPWR a_12191_10901# o_result[38] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1263 a_19513_10933# a_19347_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1264 a_10685_6031# w_dly_sig[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1265 a_11027_9269# a_11318_9569# a_11269_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1266 a_21886_6549# a_21718_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1269 w_dly_sig[59] w_dly_sig_n[58] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1270 VGND a_18298_8725# a_18256_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1271 VPWR clknet_3_4__leaf_i_stop a_19163_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1272 o_result[62] a_22863_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1273 w_dly_sig_n[57] w_dly_sig[57] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1274 o_result[62] a_22863_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1275 o_result[39] a_12050_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X1278 a_17075_8751# a_16293_8757# a_16991_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1280 o_result[21] a_8743_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1282 VPWR a_10975_8759# _64_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1286 clknet_3_5__leaf_i_stop a_21822_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1287 a_9613_9839# a_9203_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1288 w_dly_sig[2] w_dly_sig_n[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1292 a_20395_7663# a_19531_7669# a_20138_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1295 a_19697_7669# a_19531_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1296 VPWR w_dly_sig[58] w_dly_sig_n[58] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1297 w_dly_sig[28] w_dly_sig_n[27] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1298 a_10314_10749# a_10067_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1299 o_result[49] a_23047_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1301 a_21844_6953# a_21445_6581# a_21718_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1302 a_16734_9407# a_16566_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1304 a_22553_12015# w_dly_sig[64] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1307 a_16734_9407# a_16566_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1308 clknet_3_0__leaf_i_stop a_9665_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1313 VGND a_16197_9813# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1314 VGND a_17102_10495# a_17060_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1315 VGND a_19770_6549# a_19728_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1317 clknet_3_4__leaf_i_stop a_16854_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1320 VGND a_9665_7093# clknet_3_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1321 a_9866_10383# a_9479_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1322 VPWR w_dly_sig_n[59] w_dly_sig[60] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1323 a_9770_13380# a_9570_13225# a_9919_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1324 VPWR a_11311_9269# a_11318_9569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1327 a_14825_7663# w_dly_sig[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1328 VPWR w_dly_sig_n[49] w_dly_sig[50] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1331 a_16293_12021# a_16127_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1332 a_14683_9839# a_13901_9845# a_14599_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1335 VPWR clknet_0_i_stop a_14449_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1338 a_10138_10357# a_9931_10357# a_10314_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1339 VPWR w_dly_sig[56] w_dly_sig_n[56] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1340 w_dly_sig[4] w_dly_sig_n[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1341 VGND clknet_3_5__leaf_i_stop a_21279_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1342 o_result[46] a_20379_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1343 a_16063_6397# a_15281_6031# a_15979_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1344 clknet_0_i_stop a_16197_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1346 a_17267_7663# a_16403_7669# a_17010_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1348 a_10067_10383# a_9931_10357# a_9647_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1350 a_16293_9295# a_16127_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1352 w_dly_sig[54] w_dly_sig_n[53] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1353 w_dly_sig_n[23] w_dly_sig[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1358 VGND a_13847_8725# a_13805_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1361 a_11172_12559# a_10773_12559# a_11046_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1362 VPWR w_dly_sig_n[42] w_dly_sig[43] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1364 VGND clknet_3_6__leaf_i_stop a_17691_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1366 VGND a_15979_6397# a_16147_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1368 VGND a_16749_11445# clknet_3_6__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1369 VPWR a_12191_10901# a_12107_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1373 a_18498_9839# a_18059_9845# a_18413_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1376 a_18225_12015# a_17691_12021# a_18130_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1377 a_18045_8751# w_dly_sig[44] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1379 a_16297_12559# w_dly_sig[58] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1381 a_14726_10927# a_14453_10933# a_14641_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1382 VGND a_15335_8751# a_15503_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1384 a_22185_13103# w_dly_sig[63] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1385 a_9791_10217# a_9655_10057# a_9371_10071# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1387 a_19770_6549# a_19602_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1388 a_16842_7663# a_16403_7669# a_16757_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1391 VPWR a_20563_7637# a_20479_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1392 VGND a_9770_13380# a_9699_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1393 a_12981_8757# a_12815_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1394 VGND clknet_3_4__leaf_i_stop a_17691_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1395 VGND w_dly_sig[16] w_dly_sig_n[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1396 VPWR w_dly_sig[20] w_dly_sig_n[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1397 VGND a_9862_10116# a_9791_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1398 VPWR a_22879_9839# a_23047_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1400 VPWR a_21822_11471# clknet_3_7__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1401 VPWR a_22587_10901# o_result[51] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1402 VPWR a_21822_8207# clknet_3_5__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1406 a_22143_6575# a_21279_6581# a_21886_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1407 a_19820_12393# a_19421_12021# a_19694_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1410 VGND a_16734_8725# a_16692_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1412 VPWR w_dly_sig_n[19] w_dly_sig[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1415 VPWR a_9665_7093# clknet_3_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1416 o_result[46] a_20379_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1417 VGND a_17194_6549# a_17152_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1418 w_dly_sig_n[31] w_dly_sig[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1419 a_22787_6397# a_21923_6031# a_22530_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1424 VPWR a_18298_11989# a_18225_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1425 a_11766_11583# a_11598_11837# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1426 a_19517_6575# w_dly_sig[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1429 VPWR a_16854_8207# clknet_3_4__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1433 w_dly_sig[64] w_dly_sig_n[63] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1435 o_result[16] a_14767_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1436 clknet_3_7__leaf_i_stop a_21822_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1437 w_dly_sig[56] w_dly_sig_n[55] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1439 a_16968_8041# a_16569_7669# a_16842_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1440 VGND w_dly_sig[11] w_dly_sig_n[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1441 VPWR a_9389_11445# clknet_3_2__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1443 VGND clknet_0_i_stop a_14449_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1444 a_22963_9839# a_22181_9845# a_22879_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1445 VPWR a_11863_7881# a_11870_7785# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1446 a_16550_12671# a_16382_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1447 VPWR net1 w_dly_sig_n[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1449 a_22089_7119# a_21923_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1451 clknet_3_1__leaf_i_stop a_14817_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1453 VPWR clknet_0_i_stop a_16854_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1454 VPWR a_17435_7637# a_17351_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1459 a_19567_8573# a_18869_8207# a_19310_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1464 w_dly_sig_n[20] w_dly_sig[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1465 a_13330_10901# a_13162_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1466 VGND a_16991_8751# a_17159_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1467 a_17194_6549# a_17026_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1468 VPWR a_13295_11989# a_13211_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1470 a_9279_13335# a_9570_13225# a_9521_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1476 VGND clknet_3_7__leaf_i_stop a_19347_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1477 a_14342_6549# a_14174_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1478 a_10961_12559# w_dly_sig[33] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1481 a_14269_9839# a_13735_9845# a_14174_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1483 a_22530_7231# a_22362_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1485 a_9578_6397# a_9331_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1487 a_22638_9661# a_22199_9295# a_22553_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1492 VGND w_dly_sig_n[9] w_dly_sig[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1496 VPWR a_16749_11445# clknet_3_6__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1497 a_10038_9839# a_9791_10217# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1498 a_13385_7663# a_12975_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1500 VGND a_9287_12233# a_9294_12137# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1503 w_dly_sig_n[14] w_dly_sig[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1504 VGND clknet_3_5__leaf_i_stop a_21279_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1505 VGND a_12191_11739# a_12149_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1506 VGND w_dly_sig_n[54] w_dly_sig[55] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1507 VGND clknet_3_7__leaf_i_stop a_19991_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1508 o_result[2] a_13847_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1509 VGND a_14817_7093# clknet_3_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1511 w_dly_sig[24] w_dly_sig_n[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1514 o_result[31] a_9111_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1515 VPWR clknet_3_6__leaf_i_stop a_15943_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1516 w_dly_sig_n[29] w_dly_sig[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1517 clknet_3_0__leaf_i_stop a_9665_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1520 VGND w_dly_sig[8] w_dly_sig_n[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1521 a_20027_6575# a_19163_6581# a_19770_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1522 a_21822_8207# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1524 VGND a_22879_9839# a_23047_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1526 VPWR a_22311_6549# a_22227_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1529 a_15151_10927# a_14453_10933# a_14894_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1530 VGND a_16197_9813# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1533 a_18045_12015# w_dly_sig[59] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1535 VGND clknet_3_3__leaf_i_stop a_12171_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1540 VPWR a_22955_6299# a_22871_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1541 VPWR w_dly_sig[19] w_dly_sig_n[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1542 a_19912_11305# a_19513_10933# a_19786_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1543 VGND w_dly_sig[48] w_dly_sig_n[48] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1544 a_16481_8751# w_dly_sig[43] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1548 a_22530_6143# a_22362_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1549 VGND a_20566_10636# o_result[45] VGND sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X1550 a_22764_9295# a_22365_9295# a_22638_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1553 w_dly_sig[60] w_dly_sig_n[59] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1555 VPWR a_17451_6575# a_17619_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1556 VPWR w_dly_sig[54] w_dly_sig_n[54] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1558 VGND a_9374_6549# a_9332_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1559 o_result[13] a_18999_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1561 VPWR a_9655_10057# a_9662_9961# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1562 VPWR a_15503_8725# o_result[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1564 VGND clknet_3_6__leaf_i_stop a_18059_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1565 w_dly_sig_n[3] w_dly_sig[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1566 w_dly_sig_n[35] w_dly_sig[35] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1567 VGND clknet_3_6__leaf_i_stop a_16127_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1570 a_19862_11989# a_19694_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1572 a_12242_6575# a_11969_6581# a_12157_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1574 VPWR clknet_3_0__leaf_i_stop a_9319_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1576 a_9655_10057# clknet_3_2__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1578 a_17117_9295# a_16127_9295# a_16991_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1580 VGND clknet_0_i_stop a_14817_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1583 VGND a_18666_9813# a_18624_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1584 w_dly_sig_n[56] w_dly_sig[56] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1585 a_14599_9839# a_13901_9845# a_14342_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1586 a_14174_9839# a_13735_9845# a_14089_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1587 a_15281_6031# a_15115_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1588 VPWR clknet_3_7__leaf_i_stop a_19347_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1591 VPWR clknet_3_0__leaf_i_stop a_11803_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1592 clknet_3_3__leaf_i_stop a_14449_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1593 VGND a_15078_7637# a_15036_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1598 a_13993_12021# a_13827_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1599 VPWR w_dly_sig_n[28] w_dly_sig[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1601 w_dly_sig_n[18] w_dly_sig[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1603 a_19567_8573# a_18703_8207# a_19310_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1604 VPWR w_dly_sig_n[13] w_dly_sig[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1605 VPWR w_dly_sig_n[37] w_dly_sig[38] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1606 a_9749_6031# a_9195_6005# a_9402_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1608 VGND w_dly_sig[21] w_dly_sig_n[21] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1610 w_dly_sig_n[47] w_dly_sig[47] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1611 a_9749_6031# a_9202_6305# a_9402_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1612 a_9374_6549# a_9206_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1613 w_dly_sig[53] w_dly_sig_n[52] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1615 VGND a_22806_9407# a_22764_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1616 a_14825_8751# w_dly_sig[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1619 w_dly_sig_n[53] w_dly_sig[53] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1620 a_22595_10749# a_21813_10383# a_22511_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1621 a_10209_10217# a_9662_9961# a_9862_10116# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1622 a_22549_9839# a_22015_9845# a_22454_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1625 VGND a_16749_11445# clknet_3_6__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1626 a_13563_8041# a_13427_7881# a_13143_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1628 VGND clknet_0_i_stop a_21822_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1632 w_dly_sig[35] w_dly_sig_n[34] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1633 VGND a_9389_11445# clknet_3_2__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1635 a_22089_7119# a_21923_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1637 a_13713_11305# a_12723_10933# a_13587_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1638 w_dly_sig[16] w_dly_sig_n[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1639 w_dly_sig[36] w_dly_sig_n[35] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1641 a_18574_7637# a_18406_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1642 VGND a_11639_12827# a_11597_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1644 a_23063_12015# a_22365_12021# a_22806_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1646 VPWR a_21822_11471# clknet_3_7__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1647 VGND a_22587_10901# o_result[51] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1652 VPWR clknet_0_i_stop a_9389_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1653 VPWR a_21822_11471# clknet_3_7__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1655 a_12821_10217# a_12698_9961# a_12400_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0657 ps=0.725 w=0.36 l=0.15
X1656 a_13901_9845# a_13735_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1658 a_17451_6575# a_16587_6581# a_17194_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1661 a_13143_7895# a_13427_7881# a_13362_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1666 o_result[22] a_9799_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1668 a_19954_10901# a_19786_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1669 a_9195_6005# clknet_3_0__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1671 VPWR a_9665_7093# clknet_3_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1675 a_15979_6397# a_15115_6031# a_15722_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1678 a_16569_7669# a_16403_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1680 VGND a_9931_10357# a_9938_10657# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1681 VGND w_dly_sig_n[14] w_dly_sig[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1682 VPWR clknet_3_5__leaf_i_stop a_21923_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1683 a_12702_12015# a_12429_12021# a_12617_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1684 w_dly_sig_n[42] w_dly_sig[42] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1685 a_14817_7093# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1686 a_11821_7663# a_11411_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1687 VGND w_dly_sig[60] w_dly_sig_n[60] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1688 VPWR a_16854_8207# clknet_3_4__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1689 VGND a_16854_8207# clknet_3_4__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1691 a_11195_6397# a_10497_6031# a_10938_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1693 w_dly_sig[45] w_dly_sig_n[44] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1694 VPWR a_16550_12671# a_16477_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1695 a_8727_8181# a_9011_8181# a_8946_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1696 VGND clknet_3_6__leaf_i_stop a_15943_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1697 w_dly_sig[52] w_dly_sig_n[51] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1699 VGND w_dly_sig[33] w_dly_sig_n[33] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1700 a_14342_6549# a_14174_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1701 a_11325_10933# a_11159_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1703 VPWR a_12410_6549# a_12337_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1704 clknet_3_6__leaf_i_stop a_16749_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1705 w_dly_sig_n[36] w_dly_sig[36] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1706 VGND a_14449_11445# clknet_3_3__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1707 a_22089_6031# a_21923_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1708 w_dly_sig_n[32] w_dly_sig[32] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1710 VGND w_dly_sig_n[22] w_dly_sig[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1715 a_9735_11293# a_9515_11305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1716 clknet_3_5__leaf_i_stop a_21822_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1724 VPWR a_10938_6143# a_10865_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1728 w_dly_sig_n[16] w_dly_sig[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1729 VPWR a_19735_8475# a_19651_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1730 clknet_3_1__leaf_i_stop a_14817_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1732 a_21718_8751# a_21445_8757# a_21633_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1735 VPWR clknet_3_3__leaf_i_stop a_12723_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1739 VGND a_18723_11989# a_18681_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1740 VPWR a_16749_11445# clknet_3_6__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1741 VPWR w_dly_sig_n[30] w_dly_sig[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1742 VPWR a_16749_11445# clknet_3_6__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1744 VPWR a_22955_7387# o_result[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1745 VGND clknet_3_1__leaf_i_stop a_14471_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1747 a_22438_13077# a_22270_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1748 VPWR w_dly_sig[49] w_dly_sig_n[49] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1749 a_19142_8573# a_18703_8207# a_19057_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1750 VGND w_dly_sig_n[12] w_dly_sig[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1751 a_9337_10927# a_8927_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1752 VGND a_17159_9563# a_17117_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1753 a_22553_9295# w_dly_sig[49] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1754 a_20855_11837# a_19991_11471# a_20598_11583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1756 w_dly_sig_n[43] w_dly_sig[43] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1758 a_13422_8725# a_13254_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1759 clknet_3_2__leaf_i_stop a_9389_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1760 clknet_3_0__leaf_i_stop a_9665_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1763 w_dly_sig_n[30] w_dly_sig[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1764 a_17102_10495# a_16934_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1768 a_10865_6397# a_10331_6031# a_10770_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1772 a_19954_10901# a_19786_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1773 a_21997_13109# a_21831_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1775 clknet_3_4__leaf_i_stop a_16854_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1776 VPWR a_14599_6575# a_14767_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1777 a_14599_6575# a_13901_6581# a_14342_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1778 w_dly_sig_n[63] w_dly_sig[63] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1779 VPWR a_11518_9269# a_11447_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1780 VGND a_9665_7093# clknet_3_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1783 a_13422_8725# a_13254_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1786 o_result[53] a_18539_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1787 a_18923_9839# a_18225_9845# a_18666_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1789 a_9631_6575# a_8767_6581# a_9374_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1791 a_9111_13335# a_9279_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1792 a_16508_12559# a_16109_12559# a_16382_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1796 a_19049_10217# a_18059_9845# a_18923_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1797 a_16566_12015# a_16127_12021# a_16481_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1799 w_dly_sig[26] w_dly_sig_n[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1800 a_15722_6143# a_15554_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1803 VGND clknet_0_i_stop a_16749_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1804 a_16854_8207# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1805 VPWR a_13203_13077# a_13119_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1806 a_11605_8207# w_dly_sig[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1810 a_12429_12021# a_12263_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1811 o_result[45] a_20566_10636# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X1812 VGND clknet_3_6__leaf_i_stop a_19255_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1813 a_19268_8207# a_18869_8207# a_19142_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1815 VPWR a_22955_6299# o_result[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1818 a_14365_12559# w_dly_sig[35] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1819 a_20598_11583# a_20430_11837# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1822 a_23063_9661# a_22199_9295# a_22806_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1823 VGND a_21822_11471# clknet_3_7__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1825 a_22779_13103# a_21997_13109# a_22695_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1827 VGND a_19862_11989# a_19820_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1828 VGND a_18999_7637# a_18957_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1832 a_18455_10927# a_17673_10933# a_18371_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1833 VGND a_9655_10057# a_9662_9961# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1834 a_11579_7895# a_11863_7881# a_11798_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1835 w_dly_sig_n[34] w_dly_sig[34] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1837 w_dly_sig_n[40] w_dly_sig[40] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1839 VGND w_dly_sig[18] a_13981_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1841 VGND w_dly_sig[26] w_dly_sig_n[26] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1843 VGND w_dly_sig_n[60] w_dly_sig[61] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1844 a_15461_9129# a_14471_8757# a_15335_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1849 VPWR clknet_3_3__leaf_i_stop a_13827_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1850 w_dly_sig[29] w_dly_sig_n[28] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1851 VPWR w_dly_sig[52] w_dly_sig_n[52] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1852 o_result[27] a_9479_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1853 a_20211_9661# a_19513_9295# a_19954_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1856 VPWR clknet_3_4__leaf_i_stop a_18703_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1859 a_19970_7663# a_19531_7669# a_19885_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1860 VPWR a_21886_8725# a_21813_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1861 w_dly_sig_n[2] w_dly_sig[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1862 o_result[16] a_14767_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1863 VGND w_dly_sig[15] w_dly_sig_n[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1865 a_14910_7663# a_14637_7669# a_14825_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1866 a_18133_7669# a_17967_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1869 VGND w_dly_sig_n[24] w_dly_sig[25] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1870 o_result[19] a_12835_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1871 a_21721_10933# a_21555_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1872 VGND clknet_3_4__leaf_i_stop a_19163_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1873 VPWR a_9799_6549# a_9715_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1874 VGND a_19310_8319# a_19268_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1875 VPWR a_21822_8207# clknet_3_5__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1877 VGND w_dly_sig[24] w_dly_sig_n[24] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1880 VPWR clknet_0_i_stop a_21822_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1881 VGND a_21023_11739# a_20981_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1882 a_9130_6031# a_8743_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1883 a_9919_13469# a_9699_13481# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1884 VGND a_8743_6005# o_result[21] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1887 VGND w_dly_sig_n[56] w_dly_sig[57] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1890 VPWR a_17527_10651# a_17443_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1891 a_19697_10383# a_19531_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1892 VGND clknet_3_3__leaf_i_stop a_13735_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1894 a_20230_13077# a_20062_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1897 a_21813_8751# a_21279_8757# a_21718_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1898 a_15461_8041# a_14471_7669# a_15335_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1900 a_20062_13103# a_19789_13109# a_19977_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1901 VGND a_19954_10901# a_19912_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1902 a_21813_10383# a_21647_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1908 VGND a_13203_13077# a_13161_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1909 a_16109_12559# a_15943_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1910 clknet_3_5__leaf_i_stop a_21822_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1912 a_18130_8751# a_17857_8757# a_18045_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1914 w_dly_sig_n[62] w_dly_sig[62] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1915 a_14453_10933# a_14287_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1916 a_12241_8207# a_11251_8207# a_12115_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1919 VGND w_dly_sig[5] w_dly_sig_n[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1920 a_9147_8207# a_9011_8181# a_8727_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1921 w_dly_sig_n[21] w_dly_sig[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1923 clknet_3_6__leaf_i_stop a_16749_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1924 VPWR a_23231_9563# a_23147_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1927 w_dly_sig_n[64] w_dly_sig[64] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1930 VPWR w_dly_sig_n[20] w_dly_sig[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1933 VGND a_19091_9813# a_19049_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1934 VPWR w_dly_sig[41] w_dly_sig_n[41] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1935 VGND clknet_3_4__leaf_i_stop a_16127_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1937 o_result[0] a_10859_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1941 a_12617_12015# w_dly_sig[37] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1942 VGND a_16991_12015# a_17159_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1943 VGND clknet_3_7__leaf_i_stop a_22199_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1945 VGND w_dly_sig_n[48] w_dly_sig[49] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1948 clknet_3_1__leaf_i_stop a_14817_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1951 w_dly_sig[39] w_dly_sig_n[38] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1952 VGND a_22311_8725# o_result[47] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1955 a_12870_11989# a_12702_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1956 a_11279_6397# a_10497_6031# a_11195_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1957 o_result[13] a_18999_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1959 o_result[6] a_19735_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1962 a_10138_10357# a_9938_10657# a_10287_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1963 w_dly_sig[21] w_dly_sig_n[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1965 VGND w_dly_sig[59] w_dly_sig_n[59] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1966 VGND a_14817_7093# clknet_3_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1967 a_18114_10901# a_17946_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1968 VPWR clknet_3_5__leaf_i_stop a_21279_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1971 a_13161_13481# a_12171_13109# a_13035_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1972 a_12778_13077# a_12610_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1976 VPWR w_dly_sig_n[50] w_dly_sig[51] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1978 VGND a_16734_11989# a_16692_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1981 a_13330_10901# a_13162_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1982 a_19057_8207# w_dly_sig[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1984 VGND a_22311_6549# a_22269_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1985 VGND a_20195_6549# a_20153_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1990 a_13162_10927# a_12889_10933# a_13077_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1991 VPWR a_18298_8725# a_18225_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1998 a_11858_8319# a_11690_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1999 VPWR a_9195_6005# a_9202_6305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2000 clknet_3_7__leaf_i_stop a_21822_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2001 a_8911_6005# a_9195_6005# a_9130_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2003 VPWR w_dly_sig_n[52] w_dly_sig[53] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2004 VGND w_dly_sig_n[4] w_dly_sig[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2007 VGND clknet_3_4__leaf_i_stop a_18703_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2010 o_result[53] a_18539_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2012 VGND w_dly_sig[12] w_dly_sig_n[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2013 a_10773_12559# a_10607_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2014 VGND a_12283_8475# o_result[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2017 a_20211_9661# a_19347_9295# a_19954_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2018 VPWR a_18371_10927# a_18539_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2020 VPWR w_dly_sig_n[33] w_dly_sig[34] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2024 VGND a_9665_7093# clknet_3_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2026 VGND clknet_0_i_stop a_21822_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2027 VPWR a_20563_7637# o_result[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2028 o_result[54] a_17527_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2030 VPWR a_16147_6299# o_result[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2034 VGND a_22254_10495# a_22212_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2035 VGND w_dly_sig_n[47] w_dly_sig[48] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2036 a_22362_7485# a_22089_7119# a_22277_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2038 VGND a_12410_6549# a_12368_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2040 VGND a_21822_11471# clknet_3_7__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2041 a_18225_8751# a_17691_8757# a_18130_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2043 a_12525_13103# w_dly_sig[34] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2044 VPWR clknet_3_5__leaf_i_stop a_22199_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2046 VGND a_18723_8725# a_18681_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2047 o_result[47] a_22311_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2051 VGND a_16975_12827# a_16933_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2052 clknet_3_2__leaf_i_stop a_9389_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2054 VGND w_dly_sig_n[49] w_dly_sig[50] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2055 w_dly_sig[13] w_dly_sig_n[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2056 o_result[22] a_9799_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2057 a_15277_11305# a_14287_10933# a_15151_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2058 VGND a_16991_9661# a_17159_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2059 w_dly_sig_n[45] w_dly_sig[45] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2060 w_dly_sig_n[49] w_dly_sig[49] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2064 a_11513_10927# w_dly_sig[39] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2067 w_dly_sig_n[8] w_dly_sig[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2071 a_19977_13103# w_dly_sig[62] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2075 w_dly_sig[61] w_dly_sig_n[60] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2076 a_16105_6031# a_15115_6031# a_15979_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2077 a_16109_12559# a_15943_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2078 VGND w_dly_sig_n[64] g_dly_chain_even[64].dly_stg2.Y VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2079 a_16934_10749# a_16661_10383# a_16849_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2082 VPWR w_dly_sig_n[18] w_dly_sig[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2083 w_dly_sig_n[13] w_dly_sig[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2084 a_14691_12015# a_13993_12021# a_14434_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2085 VGND w_dly_sig[26] a_9473_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2086 VPWR a_22787_7485# a_22955_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2087 w_dly_sig[7] w_dly_sig_n[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2088 a_17857_8757# a_17691_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2091 o_result[24] a_8559_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2093 a_14434_11989# a_14266_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2095 a_9379_11145# clknet_3_2__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2096 VPWR a_20379_10901# a_20295_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2097 a_22227_8751# a_21445_8757# a_22143_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2098 w_dly_sig_n[6] w_dly_sig[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2099 a_20138_7637# a_19970_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2100 VPWR a_17435_7637# o_result[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2101 VPWR w_dly_sig[40] w_dly_sig_n[40] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2102 a_14266_12015# a_13993_12021# a_14181_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2105 VGND w_dly_sig[28] w_dly_sig_n[28] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2107 a_14450_12925# a_14011_12559# a_14365_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2108 a_19697_7669# a_19531_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2111 VPWR a_9665_7093# clknet_3_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2113 w_dly_sig[9] w_dly_sig_n[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2115 a_20556_11471# a_20157_11471# a_20430_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2116 VPWR a_22311_6549# o_result[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2117 w_dly_sig[57] w_dly_sig_n[56] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2119 a_15005_8751# a_14471_8757# a_14910_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2121 w_dly_sig_n[17] w_dly_sig[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2124 VPWR a_16854_8207# clknet_3_4__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2127 VGND w_dly_sig[37] w_dly_sig_n[37] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2128 o_result[6] a_19735_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2129 clknet_3_0__leaf_i_stop a_9665_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2130 o_result[4] a_15503_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2131 a_8927_11159# a_9095_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2133 VGND w_dly_sig_n[32] w_dly_sig[33] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2134 o_result[2] a_13847_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2137 VGND clknet_3_7__leaf_i_stop a_21647_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2139 clknet_0_i_stop a_16197_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2140 a_18831_7663# a_18133_7669# a_18574_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2143 a_13254_8751# a_12815_8757# a_13169_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2145 a_16757_7663# w_dly_sig[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2146 VPWR a_22787_6397# a_22955_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2147 VGND a_22311_7637# a_22269_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2148 VPWR clknet_0_i_stop a_16749_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2149 VPWR a_22530_7231# a_22457_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2150 a_23189_12393# a_22199_12021# a_23063_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2151 VPWR clknet_3_3__leaf_i_stop a_14287_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2152 clknet_3_5__leaf_i_stop a_21822_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2153 a_22806_11989# a_22638_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2154 a_14449_11445# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2155 VPWR a_9203_10071# o_result[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2156 a_14342_9813# a_14174_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2158 w_dly_sig_n[15] w_dly_sig[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2159 a_17010_7637# a_16842_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2160 VGND a_12050_9813# o_result[39] VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2161 VGND a_14599_6575# a_14767_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2163 a_22638_12015# a_22365_12021# a_22553_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2164 a_12157_6575# w_dly_sig[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2167 VGND a_20566_10636# o_result[45] VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X2168 a_10773_12559# a_10607_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2169 VPWR w_dly_sig_n[36] w_dly_sig[37] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2172 VGND w_dly_sig[25] a_9565_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2174 a_19979_10749# a_19531_10383# a_19885_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2179 a_19881_10927# a_19347_10933# a_19786_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2182 VGND a_10351_7637# a_10309_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2183 VGND a_15503_8725# o_result[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2184 o_result[12] a_20195_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2185 VGND clknet_3_0__leaf_i_stop a_11803_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2188 VGND a_23047_9813# o_result[49] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2189 a_21445_7669# a_21279_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2192 a_17485_10383# a_16495_10383# a_17359_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2193 o_result[43] a_18723_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2194 a_10497_6031# a_10331_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2196 w_dly_sig[63] w_dly_sig_n[62] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2197 VGND w_dly_sig[22] w_dly_sig_n[22] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2198 VPWR clknet_3_1__leaf_i_stop a_14471_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2200 VGND clknet_3_0__leaf_i_stop a_10331_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2202 w_dly_sig_n[44] w_dly_sig[44] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2203 a_13380_9129# a_12981_8757# a_13254_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2205 a_18130_12015# a_17691_12021# a_18045_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2206 a_21633_6575# w_dly_sig[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2208 a_9275_9295# a_9055_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2212 w_dly_sig[10] w_dly_sig_n[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2213 VPWR a_20655_13077# a_20571_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2214 a_19786_9661# a_19347_9295# a_19701_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2216 VGND a_17619_6549# a_17577_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2218 VGND w_dly_sig[27] a_10209_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2219 VPWR a_19091_9813# o_result[44] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2220 a_21886_6549# a_21718_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2223 a_12981_8757# a_12815_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2225 VGND w_dly_sig_n[29] w_dly_sig[30] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2226 clknet_3_7__leaf_i_stop a_21822_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2227 a_8635_9269# a_8926_9569# a_8877_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2228 VGND w_dly_sig_n[44] w_dly_sig[45] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2230 clknet_3_7__leaf_i_stop a_21822_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2231 VPWR w_dly_sig_n[7] w_dly_sig[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2234 VPWR a_19954_10901# a_19881_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2236 VGND a_16147_6299# a_16105_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2244 VPWR clknet_3_2__leaf_i_stop a_10607_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2245 w_dly_sig[18] w_dly_sig_n[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2246 w_dly_sig_n[27] w_dly_sig[27] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2248 a_13587_10927# a_12889_10933# a_13330_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2250 a_21445_6581# a_21279_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2252 a_12667_6575# a_11803_6581# a_12410_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2253 VGND w_dly_sig_n[53] w_dly_sig[54] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2254 VPWR a_11858_8319# a_11785_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2258 VGND a_12191_11739# o_result[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2259 a_9126_9269# a_8926_9569# a_9275_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2260 a_17857_12021# a_17691_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2261 VGND a_17359_10749# a_17527_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2262 VGND a_21822_8207# clknet_3_5__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2263 VGND a_21822_11471# clknet_3_7__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2264 a_19912_9295# a_19513_9295# a_19786_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2265 VPWR w_dly_sig_n[6] w_dly_sig[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2267 VPWR a_18831_7663# a_18999_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2268 VGND a_10138_10357# a_10067_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2270 clknet_3_2__leaf_i_stop a_9389_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2271 VPWR clknet_3_3__leaf_i_stop a_14011_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2273 VPWR a_8835_12247# o_result[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2274 VGND a_16197_9813# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2276 VGND a_11863_7881# a_11870_7785# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2277 a_14641_10927# w_dly_sig[56] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2280 VPWR a_21822_8207# clknet_3_5__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2283 a_20138_7637# a_19970_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2285 VGND a_16197_9813# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2286 VPWR a_10351_7637# o_result[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2288 VGND a_23231_11989# a_23189_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2289 VPWR a_8919_9269# a_8926_9569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2290 VGND w_dly_sig[1] w_dly_sig_n[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2292 a_11785_8573# a_11251_8207# a_11690_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2293 a_9367_8207# a_9147_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2294 a_13981_8041# a_13434_7785# a_13634_7940# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2298 VPWR a_14817_7093# clknet_3_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2300 VGND a_11214_12671# a_11172_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2301 g_dly_chain_even[64].dly_stg2.Y w_dly_sig_n[64] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2302 VPWR a_13755_10901# a_13671_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2304 VPWR w_dly_sig[7] w_dly_sig_n[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2305 VPWR a_12070_7940# a_11999_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2306 a_22254_10495# a_22086_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2309 clknet_3_2__leaf_i_stop a_9389_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2311 a_9946_13103# a_9699_13481# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2312 a_19789_12015# a_19255_12021# a_19694_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2313 w_dly_sig[40] w_dly_sig_n[39] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2316 w_dly_sig_n[33] w_dly_sig[33] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2317 a_18624_10217# a_18225_9845# a_18498_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2318 a_15419_8751# a_14637_8757# a_15335_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2321 a_9473_9295# a_8919_9269# a_9126_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2322 clknet_3_1__leaf_i_stop a_14817_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2323 VPWR a_15078_7637# a_15005_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2324 VPWR clknet_3_2__leaf_i_stop a_11159_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2327 VPWR w_dly_sig[39] w_dly_sig_n[39] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2328 VGND a_19954_9407# a_19912_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2329 VGND a_20655_13077# a_20613_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2330 a_22181_9845# a_22015_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2333 VPWR w_dly_sig[45] w_dly_sig_n[45] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2335 VGND w_dly_sig[14] w_dly_sig_n[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2338 o_result[54] a_17527_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2340 a_16749_11445# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2341 clknet_3_7__leaf_i_stop a_21822_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2342 VGND w_dly_sig_n[2] w_dly_sig[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2343 a_11471_12925# a_10607_12559# a_11214_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2346 VPWR w_dly_sig_n[63] w_dly_sig[64] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2347 VGND a_11518_9269# a_11447_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2348 a_22162_10901# a_21994_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2350 VPWR a_17619_6549# o_result[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2351 VGND a_9799_6549# a_9757_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2352 a_9521_13103# a_9111_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2354 VGND w_dly_sig[25] w_dly_sig_n[25] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2355 a_11141_12925# a_10607_12559# a_11046_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2356 a_18666_9813# a_18498_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2360 VGND a_12115_8573# a_12283_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2364 o_result[42] a_17159_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2365 w_dly_sig[12] w_dly_sig_n[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2366 VGND a_9389_11445# clknet_3_2__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2367 a_9218_8181# a_9018_8481# a_9367_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2368 clknet_3_5__leaf_i_stop a_21822_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2369 a_17010_7637# a_16842_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2373 w_dly_sig_n[37] w_dly_sig[37] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2375 VPWR a_12835_6549# a_12751_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2376 VPWR a_9631_6575# a_9799_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2380 VGND w_dly_sig_n[23] w_dly_sig[24] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2381 VPWR a_20395_7663# a_20563_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2382 VPWR a_15979_6397# a_16147_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2385 VGND a_15503_7637# a_15461_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2386 VPWR a_16749_11445# clknet_3_6__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2388 clknet_3_0__leaf_i_stop a_9665_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2391 w_dly_sig_n[1] w_dly_sig[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2393 VPWR clknet_0_i_stop a_9389_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2394 a_21822_8207# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2396 a_20613_13481# a_19623_13109# a_20487_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2397 clknet_3_3__leaf_i_stop a_14449_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2398 VPWR w_dly_sig[10] w_dly_sig_n[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2399 clknet_3_4__leaf_i_stop a_16854_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2400 VGND clknet_3_0__leaf_i_stop a_9319_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2405 clknet_3_1__leaf_i_stop a_14817_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2406 VPWR a_11214_12671# a_11141_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2407 a_18406_7663# a_17967_7669# a_18321_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2408 VGND a_18298_11989# a_18256_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2409 o_result[45] a_20566_10636# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X2412 VGND clknet_3_2__leaf_i_stop a_10607_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2413 w_dly_sig[37] w_dly_sig_n[36] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2414 a_20157_11471# a_19991_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2415 a_14894_10901# a_14726_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2416 VPWR a_8467_9269# o_result[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2418 w_dly_sig[1] w_dly_sig_n[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2420 VPWR a_14859_11989# a_14775_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2421 VGND w_dly_sig[29] w_dly_sig_n[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2422 a_9565_8207# a_9011_8181# a_9218_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2424 VGND a_14817_7093# clknet_3_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2425 a_14637_7669# a_14471_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2426 a_16854_8207# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2429 VGND a_14767_6549# a_14725_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2430 VGND a_20563_7637# o_result[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2433 w_dly_sig[3] w_dly_sig_n[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2434 a_20211_10927# a_19513_10933# a_19954_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2435 a_9126_9269# a_8919_9269# a_9302_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2438 VPWR clknet_3_3__leaf_i_stop a_12263_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2439 w_dly_sig_n[25] w_dly_sig[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2442 a_16941_6575# w_dly_sig[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2445 VPWR w_dly_sig_n[17] w_dly_sig[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2446 VPWR a_17267_7663# a_17435_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2447 a_12337_13109# a_12171_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2449 VGND clknet_3_3__leaf_i_stop a_14011_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2453 w_dly_sig[17] w_dly_sig_n[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2455 a_17194_6549# a_17026_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2456 w_dly_sig_n[5] w_dly_sig[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2458 a_19701_9295# w_dly_sig[47] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2461 w_dly_sig_n[22] w_dly_sig[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2462 VGND w_dly_sig_n[15] w_dly_sig[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2463 clknet_3_7__leaf_i_stop a_21822_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2466 VGND w_dly_sig_n[61] w_dly_sig[62] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2469 a_18532_8041# a_18133_7669# a_18406_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2470 w_dly_sig[30] w_dly_sig_n[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2471 VGND i_stop a_16197_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2473 a_22438_13077# a_22270_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2474 VPWR a_13427_7881# a_13434_7785# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2478 a_22270_13103# a_21997_13109# a_22185_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2479 a_9302_9661# a_9055_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2482 a_16753_6581# a_16587_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2483 a_16991_12015# a_16127_12021# a_16734_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2485 a_13077_10927# w_dly_sig[38] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2489 clknet_3_4__leaf_i_stop a_16854_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2491 VGND a_17435_7637# o_result[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2494 a_16661_12015# a_16127_12021# a_16566_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2495 a_20138_10519# a_19979_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X2496 w_dly_sig_n[51] w_dly_sig[51] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2498 VPWR w_dly_sig[50] w_dly_sig_n[50] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2499 a_14174_9839# a_13901_9845# a_14089_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2500 VPWR a_16197_9813# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2502 VPWR a_20027_6575# a_20195_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2503 a_20027_6575# a_19329_6581# a_19770_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2504 o_result[29] a_12191_11739# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2508 VPWR a_22143_6575# a_22311_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2509 a_22143_6575# a_21445_6581# a_21886_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2510 a_11579_7895# a_11870_7785# a_11821_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2512 a_12199_8573# a_11417_8207# a_12115_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2515 VGND w_dly_sig_n[10] w_dly_sig[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2517 a_16891_12925# a_16109_12559# a_16807_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2518 VPWR clknet_3_3__leaf_i_stop a_13735_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2519 VPWR a_21822_8207# clknet_3_5__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2521 VPWR w_dly_sig[53] w_dly_sig_n[53] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2523 a_14449_11445# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2525 o_result[30] a_8835_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2526 VGND w_dly_sig[47] w_dly_sig_n[47] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2527 VGND w_dly_sig_n[34] w_dly_sig[35] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2529 o_result[4] a_15503_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2531 a_14300_10217# a_13901_9845# a_14174_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2533 VGND w_dly_sig[22] a_9749_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2536 a_21886_7637# a_21718_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2537 w_dly_sig[5] w_dly_sig_n[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2538 VGND w_dly_sig_n[46] w_dly_sig[47] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2542 VPWR a_16734_11989# a_16661_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2543 a_9498_13469# a_9111_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2544 a_11598_11837# a_11325_11471# a_11513_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2545 clknet_3_2__leaf_i_stop a_9389_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2546 VPWR a_11411_7895# o_result[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2547 VGND clknet_3_7__leaf_i_stop a_21831_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2549 VPWR w_dly_sig_n[21] w_dly_sig[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2551 clknet_3_6__leaf_i_stop a_16749_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2552 a_14181_12015# w_dly_sig[36] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2554 w_dly_sig_n[9] w_dly_sig[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2556 a_18555_8751# a_17857_8757# a_18298_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2559 a_9931_10357# clknet_3_2__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2560 a_9926_7637# a_9758_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2563 a_9670_12015# a_9423_12393# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2564 VGND a_11311_9269# a_11318_9569# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2568 VPWR a_17359_10749# a_17527_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2573 VPWR w_dly_sig_n[51] w_dly_sig[52] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2576 w_dly_sig_n[12] w_dly_sig[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2577 a_9374_6549# a_9206_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2578 a_11766_10901# a_11598_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2579 VPWR w_dly_sig[32] a_10117_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2580 VGND w_dly_sig[36] w_dly_sig_n[36] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2581 a_22787_7485# a_22089_7119# a_22530_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2582 a_19885_7663# w_dly_sig[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2583 VPWR w_dly_sig[32] w_dly_sig_n[32] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2584 a_9055_9295# a_8926_9569# a_8635_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2586 a_13035_13103# a_12337_13109# a_12778_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2587 a_9473_9295# a_8926_9569# a_9126_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2588 a_18555_8751# a_17691_8757# a_18298_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2589 a_14817_12393# a_13827_12021# a_14691_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2590 a_16734_8725# a_16566_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2591 a_12623_10205# a_12050_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.12 ps=1.41 w=0.42 l=0.15
X2592 VGND a_8467_9269# o_result[25] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2593 a_22553_9295# w_dly_sig[49] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2594 a_20395_7663# a_19697_7669# a_20138_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2595 w_dly_sig_n[59] w_dly_sig[59] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2596 a_16293_9295# a_16127_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2597 a_14825_8751# w_dly_sig[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2599 VPWR a_18923_9839# a_19091_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2600 a_16991_9661# a_16127_9295# a_16734_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2603 clknet_3_0__leaf_i_stop a_9665_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2607 VPWR a_14342_9813# a_14269_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2608 a_8933_6581# a_8767_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2611 a_9402_6005# a_9195_6005# a_9578_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2612 a_9494_12292# a_9287_12233# a_9670_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2613 clknet_3_3__leaf_i_stop a_14449_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2614 a_19007_9839# a_18225_9845# a_18923_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2615 a_22553_12015# w_dly_sig[64] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2616 w_dly_sig[47] w_dly_sig_n[46] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2617 clknet_3_3__leaf_i_stop a_14449_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2618 a_12889_10933# a_12723_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2621 a_9423_12393# a_9287_12233# a_9003_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2622 a_9862_10116# a_9655_10057# a_10038_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2623 a_22454_9839# a_22181_9845# a_22369_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2626 a_11269_9661# a_10859_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2629 a_10117_13481# a_9563_13321# a_9770_13380# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2630 a_20939_11837# a_20157_11471# a_20855_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2631 VGND a_19735_8475# a_19693_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2633 VPWR a_23231_9563# o_result[48] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2636 a_20395_10749# a_19531_10383# a_20138_10519# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2639 VGND w_dly_sig[30] w_dly_sig_n[30] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2640 a_22787_6397# a_22089_6031# a_22530_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2641 a_16937_7663# a_16403_7669# a_16842_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2643 a_9862_10116# a_9662_9961# a_10011_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2646 a_9551_6031# a_9331_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2648 a_9563_13321# clknet_3_2__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2649 a_14365_12559# w_dly_sig[35] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2650 w_dly_sig[48] w_dly_sig_n[47] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2651 w_dly_sig_n[4] w_dly_sig[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2653 VPWR a_20195_6549# a_20111_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2655 a_17267_7663# a_16569_7669# a_17010_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2656 o_result[47] a_22311_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2657 a_8835_12247# a_9003_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2659 VGND w_dly_sig[31] a_9841_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2660 VPWR a_18539_10901# o_result[53] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2661 a_18133_7669# a_17967_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2663 VPWR a_22587_10901# a_22503_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2664 w_dly_sig[22] w_dly_sig_n[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2666 VPWR a_9770_13380# a_9699_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2667 a_21718_8751# a_21279_8757# a_21633_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2670 a_9147_8207# a_9018_8481# a_8727_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2673 a_12870_11989# a_12702_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2675 VGND a_23047_9813# a_23005_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2677 a_13901_6581# a_13735_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2678 a_11766_10901# a_11598_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2679 VGND a_8559_8181# o_result[24] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2683 VGND w_dly_sig_n[31] w_dly_sig[32] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2685 a_22143_7663# a_21279_7669# a_21886_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2687 a_11598_10927# a_11325_10933# a_11513_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2693 a_12070_7940# a_11863_7881# a_12246_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2695 VPWR a_14449_11445# clknet_3_3__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2696 VPWR a_20138_10519# a_20072_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X2697 VPWR w_dly_sig_n[3] w_dly_sig[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2699 _64_.X a_10975_8759# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2700 VPWR a_18723_8725# a_18639_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2701 VGND w_dly_sig[34] w_dly_sig_n[34] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2703 a_9402_6005# a_9202_6305# a_9551_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2704 a_22787_7485# a_21923_7119# a_22530_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2705 clknet_0_i_stop a_16197_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2706 VGND a_16550_12671# a_16508_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2707 VPWR w_dly_sig[28] a_10485_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2708 VGND a_21822_8207# clknet_3_5__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2709 a_16692_12393# a_16293_12021# a_16566_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2711 a_12400_9813# a_12688_10057# a_12623_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.066 ps=0.745 w=0.36 l=0.15
X2712 w_dly_sig[44] w_dly_sig_n[43] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2713 a_16991_8751# a_16293_8757# a_16734_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2715 VGND w_dly_sig_n[5] w_dly_sig[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2716 a_9095_11159# a_9386_11049# a_9337_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2717 VGND a_9379_11145# a_9386_11049# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2719 a_10183_7663# a_9319_7669# a_9926_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2720 w_dly_sig[27] w_dly_sig_n[26] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2721 a_17451_6575# a_16753_6581# a_17194_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2723 VPWR a_9479_10357# o_result[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2725 a_14618_12671# a_14450_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2726 VPWR a_15319_10901# a_15235_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2727 a_21844_9129# a_21445_8757# a_21718_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2728 VGND w_dly_sig_n[19] w_dly_sig[20] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2730 a_11766_11583# a_11598_11837# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2731 a_18371_10927# a_17673_10933# a_18114_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2733 VPWR clknet_0_i_stop a_9665_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2734 a_11417_8207# a_11251_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2735 VGND a_9665_7093# clknet_3_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2737 w_dly_sig_n[28] w_dly_sig[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2738 a_21718_7663# a_21279_7669# a_21633_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2739 VGND a_14859_11989# a_14817_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2740 VPWR a_21822_8207# clknet_3_5__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2741 VGND a_17619_6549# o_result[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2742 a_9770_13380# a_9563_13321# a_9946_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2745 VPWR a_22622_9813# a_22549_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2748 clknet_3_3__leaf_i_stop a_14449_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2750 a_12246_7663# a_11999_8041# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2751 a_11447_9295# a_11311_9269# a_11027_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2752 a_16807_12925# a_15943_12559# a_16550_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2753 VGND w_dly_sig[44] w_dly_sig_n[44] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2755 VGND a_16854_8207# clknet_3_4__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2757 VPWR w_dly_sig_n[57] w_dly_sig[58] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2758 a_16991_8751# a_16127_8757# a_16734_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2760 VPWR a_14817_7093# clknet_3_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2761 a_16477_12925# a_15943_12559# a_16382_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2762 a_23063_9661# a_22365_9295# a_22806_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2764 a_10770_6397# a_10497_6031# a_10685_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2767 VPWR a_8927_11159# o_result[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2768 clknet_0_i_stop a_16197_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2770 a_11858_8319# a_11690_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2775 VPWR a_19091_9813# a_19007_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2776 VGND a_20395_7663# a_20563_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2780 VPWR a_8743_6005# o_result[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2782 VPWR a_16854_8207# clknet_3_4__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2784 clknet_3_1__leaf_i_stop a_14817_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2785 clknet_3_2__leaf_i_stop a_9389_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2787 VGND clknet_0_i_stop a_16854_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2790 a_8911_6005# a_9202_6305# a_9153_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2792 w_dly_sig_n[38] w_dly_sig[38] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2796 a_20479_7663# a_19697_7669# a_20395_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2797 VGND a_9494_12292# a_9423_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2798 VGND clknet_3_5__leaf_i_stop a_21279_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2799 w_dly_sig[19] w_dly_sig_n[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2801 w_dly_sig_n[58] w_dly_sig[58] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2805 VPWR a_22863_13077# a_22779_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2809 VPWR w_dly_sig_n[55] w_dly_sig[56] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2810 a_21844_8041# a_21445_7669# a_21718_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2813 clknet_3_2__leaf_i_stop a_9389_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2815 VGND a_15043_12827# a_15001_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2816 a_20245_12393# a_19255_12021# a_20119_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2818 VGND a_11363_6299# o_result[20] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2819 w_dly_sig[14] w_dly_sig_n[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2820 o_result[29] a_12191_11739# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2821 VPWR a_22311_7637# a_22227_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2822 VGND w_dly_sig[62] w_dly_sig_n[62] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2823 VGND a_14449_11445# clknet_3_3__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2824 a_17359_10749# a_16661_10383# a_17102_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2826 o_result[43] a_18723_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2828 a_22369_9839# w_dly_sig[50] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2829 a_11999_8041# a_11870_7785# a_11579_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2831 a_11311_9269# clknet_3_3__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2833 VGND a_12835_6549# a_12793_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2834 a_9121_6575# w_dly_sig[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2835 w_dly_sig_n[41] w_dly_sig[41] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2836 a_18130_8751# a_17691_8757# a_18045_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2840 VPWR a_22955_7387# a_22871_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2841 o_result[56] a_17159_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2842 clknet_3_0__leaf_i_stop a_9665_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2844 o_result[56] a_17159_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2846 VGND w_dly_sig_n[25] w_dly_sig[26] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2847 VGND a_17267_7663# a_17435_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2849 a_22365_12021# a_22199_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2850 VGND clknet_3_7__leaf_i_stop a_19347_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2851 VGND w_dly_sig[50] w_dly_sig_n[50] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2852 a_20337_9295# a_19347_9295# a_20211_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2853 a_21822_8207# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2855 VGND a_11363_6299# a_11321_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2856 a_12023_10927# a_11325_10933# a_11766_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2857 a_21445_6581# a_21279_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2858 VPWR a_10351_7637# a_10267_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2859 VPWR a_20379_9563# o_result[46] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2860 VPWR net1 a_10975_8759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2862 VPWR w_dly_sig_n[38] w_dly_sig[39] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2863 w_dly_sig[41] w_dly_sig_n[40] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2867 a_22362_7485# a_21923_7119# a_22277_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2873 VGND w_dly_sig[23] w_dly_sig_n[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2876 VGND w_dly_sig[19] w_dly_sig_n[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2880 VPWR a_9389_11445# clknet_3_2__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2881 a_9631_6575# a_8933_6581# a_9374_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2882 a_19421_12021# a_19255_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2883 a_21994_10927# a_21721_10933# a_21909_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2884 a_12417_8041# a_11870_7785# a_12070_7940# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2886 a_9003_12247# a_9294_12137# a_9245_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2888 a_17075_12015# a_16293_12021# a_16991_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2889 VPWR a_18555_12015# a_18723_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2890 w_dly_sig[2] w_dly_sig_n[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2891 clknet_3_4__leaf_i_stop a_16854_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2893 VPWR clknet_3_7__leaf_i_stop a_19623_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2894 VGND a_18555_12015# a_18723_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2895 VGND a_15078_8725# a_15036_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2896 a_19602_6575# a_19163_6581# a_19517_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2900 w_dly_sig_n[3] w_dly_sig[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2903 a_13805_9129# a_12815_8757# a_13679_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2904 a_18256_9129# a_17857_8757# a_18130_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2905 a_15979_6397# a_15281_6031# a_15722_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2906 VGND a_12975_7895# o_result[17] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2907 clknet_0_i_stop a_16197_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2909 a_9279_13335# a_9563_13321# a_9498_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2914 VGND a_22679_10651# a_22637_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2916 VGND a_22143_6575# a_22311_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2917 VGND a_20027_6575# a_20195_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2918 VGND a_9563_13321# a_9570_13225# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2919 w_dly_sig_n[0] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2921 VGND a_18539_10901# o_result[53] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2922 w_dly_sig_n[60] w_dly_sig[60] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2923 a_10485_10383# a_9931_10357# a_10138_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2925 a_11417_8207# a_11251_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2927 a_17857_8757# a_17691_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2930 a_14910_8751# a_14471_8757# a_14825_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2932 a_18555_12015# a_17691_12021# a_18298_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2934 VGND a_22863_13077# a_22821_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2935 a_22488_7119# a_22089_7119# a_22362_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2936 a_22362_6397# a_21923_6031# a_22277_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2938 o_result[0] a_10859_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2939 VPWR w_dly_sig[31] w_dly_sig_n[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2940 VGND a_14342_9813# a_14300_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2941 VPWR w_dly_sig[18] w_dly_sig_n[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2943 a_20096_8041# a_19697_7669# a_19970_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2944 o_result[57] a_16975_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2945 VGND a_17527_10651# o_result[54] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2947 a_15335_7663# a_14471_7669# a_15078_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2949 VGND a_21822_11471# clknet_3_7__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2952 VPWR a_12688_10057# a_12698_9961# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2953 a_10859_9269# a_11027_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2954 VGND a_20379_9563# o_result[46] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2956 w_dly_sig[32] w_dly_sig_n[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2957 VPWR a_14449_11445# clknet_3_3__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2958 VPWR w_dly_sig[26] a_9473_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2959 a_19728_6953# a_19329_6581# a_19602_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2963 VPWR a_14449_11445# clknet_3_3__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2965 a_22638_9661# a_22365_9295# a_22553_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2967 w_dly_sig[54] w_dly_sig_n[53] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2968 a_20337_11305# a_19347_10933# a_20211_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2973 clknet_0_i_stop a_16197_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2975 VPWR a_14767_6549# o_result[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2976 VPWR clknet_3_5__leaf_i_stop a_21923_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2977 VGND a_19567_8573# a_19735_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2980 VGND a_20287_11989# a_20245_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2981 a_11598_10927# a_11159_10933# a_11513_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2982 VPWR clknet_0_i_stop a_21822_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2983 a_16749_11445# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2984 VGND a_22530_7231# a_22488_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2985 VGND a_9665_7093# clknet_3_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2986 clknet_3_7__leaf_i_stop a_21822_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2988 a_14910_7663# a_14471_7669# a_14825_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2989 a_9389_11445# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2992 a_22821_13481# a_21831_13109# a_22695_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2993 a_22488_6031# a_22089_6031# a_22362_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2995 clknet_3_3__leaf_i_stop a_14449_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2996 o_result[42] a_17159_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2999 w_dly_sig_n[55] w_dly_sig[55] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3000 VGND a_16854_8207# clknet_3_4__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3001 VGND a_20138_10519# a_20076_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X3002 VPWR w_dly_sig[64] w_dly_sig_n[64] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3004 VGND a_22511_10749# a_22679_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3005 a_16566_8751# a_16127_8757# a_16481_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3007 w_dly_sig[58] w_dly_sig_n[57] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3008 VPWR a_21822_8207# clknet_3_5__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3010 a_17026_6575# a_16587_6581# a_16941_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3012 VGND a_20379_9563# a_20337_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3013 a_14089_6575# w_dly_sig[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3014 VGND a_20230_13077# a_20188_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3015 a_11513_11471# w_dly_sig[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3016 VPWR a_12283_8475# o_result[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3018 a_21445_7669# a_21279_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3020 a_20487_13103# a_19789_13109# a_20230_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3021 VPWR a_13847_8725# o_result[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3022 clknet_3_5__leaf_i_stop a_21822_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3025 a_12892_10116# a_12688_10057# a_13074_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0693 ps=0.75 w=0.42 l=0.15
X3026 VPWR a_18723_11989# o_result[58] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3028 VGND clknet_3_1__leaf_i_stop a_14471_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3030 VGND a_18723_11989# o_result[58] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3031 VPWR w_dly_sig[46] w_dly_sig_n[46] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3036 clknet_3_1__leaf_i_stop a_14817_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3038 VGND a_22530_6143# a_22488_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3043 w_dly_sig[56] w_dly_sig_n[55] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3044 VGND w_dly_sig[46] w_dly_sig_n[46] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3046 w_dly_sig[6] w_dly_sig_n[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3047 a_9331_6031# a_9202_6305# a_8911_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3048 w_dly_sig[11] w_dly_sig_n[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3049 VPWR a_15503_7637# a_15419_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3054 a_14576_12559# a_14177_12559# a_14450_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3055 a_16661_10383# a_16495_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3056 a_23005_10217# a_22015_9845# a_22879_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3057 a_16692_9129# a_16293_8757# a_16566_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3058 VGND a_11411_7895# o_result[18] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3060 clknet_3_1__leaf_i_stop a_14817_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3064 a_17152_6953# a_16753_6581# a_17026_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3065 VGND a_20598_11583# a_20556_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3066 VPWR a_22806_9407# a_22733_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3069 a_12410_6549# a_12242_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3071 clknet_3_0__leaf_i_stop a_9665_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3072 VPWR a_18999_7637# o_result[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3074 a_13169_8751# w_dly_sig[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3077 w_dly_sig[40] w_dly_sig_n[39] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3078 VPWR a_16991_12015# a_17159_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3084 a_9485_7669# a_9319_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3085 w_dly_sig_n[39] w_dly_sig[39] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3086 w_dly_sig_n[50] w_dly_sig[50] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3087 clknet_3_4__leaf_i_stop a_16854_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3088 a_16753_6581# a_16587_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3089 clknet_3_6__leaf_i_stop a_16749_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3093 VPWR a_17159_9563# a_17075_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3095 VGND a_12778_13077# a_12736_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3096 a_11969_6581# a_11803_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3099 VPWR a_9389_11445# clknet_3_2__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3100 VPWR w_dly_sig_n[54] w_dly_sig[55] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3101 a_15281_6031# a_15115_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3102 w_dly_sig[62] w_dly_sig_n[61] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3104 a_22277_7119# w_dly_sig[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3105 a_9665_7093# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3108 w_dly_sig[38] w_dly_sig_n[37] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3109 a_16854_8207# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3112 clknet_3_5__leaf_i_stop a_21822_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3114 a_9494_12292# a_9294_12137# a_9643_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3115 a_22733_9661# a_22199_9295# a_22638_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3118 VPWR w_dly_sig[43] w_dly_sig_n[43] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3119 a_17673_10933# a_17507_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3123 VGND clknet_3_5__leaf_i_stop a_21923_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3124 VPWR a_21023_11739# a_20939_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3125 a_10859_9269# a_11027_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3129 a_21994_10927# a_21555_10933# a_21909_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3130 VPWR a_16197_9813# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3131 clknet_3_3__leaf_i_stop a_14449_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3132 VPWR w_dly_sig[22] a_9749_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3133 VGND a_17451_6575# a_17619_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3134 a_9206_6575# a_8767_6581# a_9121_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3136 VPWR w_dly_sig[61] w_dly_sig_n[61] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3137 a_14910_8751# a_14637_8757# a_14825_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3139 a_16757_7663# w_dly_sig[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3140 VGND w_dly_sig_n[62] w_dly_sig[63] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3142 VPWR w_dly_sig[38] w_dly_sig_n[38] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3144 VGND a_12023_11837# a_12191_11739# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3145 clknet_3_4__leaf_i_stop a_16854_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3147 VPWR w_dly_sig_n[58] w_dly_sig[59] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3148 a_18957_8041# a_17967_7669# a_18831_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3149 a_11798_8029# a_11411_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3151 VGND w_dly_sig_n[45] w_dly_sig[46] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3153 a_17535_6575# a_16753_6581# a_17451_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3154 a_18256_12393# a_17857_12021# a_18130_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3155 a_9647_10357# a_9931_10357# a_9866_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3157 VGND a_11195_6397# a_11363_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3158 VGND a_16749_11445# clknet_3_6__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3159 a_11513_10927# w_dly_sig[39] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3160 VPWR a_9799_6549# o_result[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3161 a_16550_12671# a_16382_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3163 a_22277_6031# w_dly_sig[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3165 net1 a_855_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3167 VGND a_16807_12925# a_16975_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3168 w_dly_sig_n[11] w_dly_sig[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3170 VPWR a_14449_11445# clknet_3_3__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3172 w_dly_sig_n[23] w_dly_sig[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3173 VPWR a_14449_11445# clknet_3_3__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3174 o_result[39] a_12050_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3175 VPWR w_dly_sig[42] w_dly_sig_n[42] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3177 VGND a_21822_8207# clknet_3_5__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3179 a_10485_10383# a_9938_10657# a_10138_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3182 a_14177_12559# a_14011_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3183 a_14599_9839# a_13735_9845# a_14342_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3184 VGND clknet_3_5__leaf_i_stop a_21923_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3188 a_9332_6953# a_8933_6581# a_9206_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3189 a_14726_10927# a_14287_10933# a_14641_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3190 a_13253_12393# a_12263_12021# a_13127_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3194 VPWR a_20211_9661# a_20379_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3197 VPWR a_21822_8207# clknet_3_5__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3199 clknet_3_6__leaf_i_stop a_16749_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3202 a_21822_11471# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3203 VPWR clknet_3_6__leaf_i_stop a_16127_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3204 a_14174_6575# a_13735_6581# a_14089_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3206 a_9389_11445# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3207 VGND w_dly_sig[28] a_10485_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3210 a_8933_6581# a_8767_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3211 VGND a_12892_10116# a_12821_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0989 ps=0.995 w=0.64 l=0.15
X3213 VPWR a_14817_7093# clknet_3_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3215 a_14266_12015# a_13827_12021# a_14181_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3216 VPWR w_dly_sig[16] w_dly_sig_n[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3217 clknet_0_i_stop a_16197_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3220 a_22181_9845# a_22015_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3223 a_14821_10927# a_14287_10933# a_14726_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3230 VPWR a_16854_8207# clknet_3_4__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3231 VPWR a_17527_10651# o_result[54] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3232 VPWR a_17159_8725# a_17075_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3233 VGND w_dly_sig_n[43] w_dly_sig[44] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3236 a_11555_12925# a_10773_12559# a_11471_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3237 a_14637_7669# a_14471_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3239 a_9586_11204# a_9386_11049# a_9735_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3241 a_9371_10071# a_9662_9961# a_9613_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3242 a_8927_11159# a_9095_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3243 VGND w_dly_sig_n[26] w_dly_sig[27] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3245 a_18497_11305# a_17507_10933# a_18371_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3246 w_dly_sig[43] w_dly_sig_n[42] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3247 VPWR clknet_3_1__leaf_i_stop a_12815_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3249 o_result[58] a_18723_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3253 clknet_3_1__leaf_i_stop a_14817_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3254 clknet_3_0__leaf_i_stop a_9665_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3256 o_result[58] a_18723_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3258 a_12410_6549# a_12242_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3259 a_14300_6953# a_13901_6581# a_14174_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3261 a_12617_12015# w_dly_sig[37] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3264 VGND a_11471_12925# a_11639_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3265 VGND a_15722_6143# a_15680_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3275 a_13993_12021# a_13827_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3276 VPWR a_14894_10901# a_14821_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3278 w_dly_sig[55] w_dly_sig_n[54] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3280 VGND a_19091_9813# o_result[44] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3282 a_13901_6581# a_13735_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3284 a_22638_12015# a_22199_12021# a_22553_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3286 VPWR clknet_3_6__leaf_i_stop a_16495_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3288 VPWR a_20195_6549# o_result[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3289 VGND a_15319_10901# a_15277_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3291 w_dly_sig_n[20] w_dly_sig[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3292 VGND a_13427_7881# a_13434_7785# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3293 VGND clknet_3_5__leaf_i_stop a_22199_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3298 VPWR a_14767_9813# a_14683_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3301 VGND w_dly_sig[13] w_dly_sig_n[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3303 a_23147_9661# a_22365_9295# a_23063_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3304 a_16734_11989# a_16566_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3305 clknet_3_6__leaf_i_stop a_16749_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3306 a_20430_11837# a_20157_11471# a_20345_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3307 a_22879_9839# a_22015_9845# a_22622_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3308 a_11690_8573# a_11417_8207# a_11605_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3310 clknet_3_6__leaf_i_stop a_16749_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3313 VPWR a_16147_6299# a_16063_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3314 a_13634_7940# a_13427_7881# a_13810_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3315 VGND a_9479_10357# o_result[27] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3316 a_19701_9295# w_dly_sig[47] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3325 a_16934_10749# a_16495_10383# a_16849_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3326 VPWR a_9389_11445# clknet_3_2__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3329 VGND w_dly_sig[35] w_dly_sig_n[35] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3331 VGND a_13634_7940# a_13563_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3333 VGND w_dly_sig[57] w_dly_sig_n[57] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3335 a_18869_8207# a_18703_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3337 a_12667_6575# a_11969_6581# a_12410_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3338 a_14177_12559# a_14011_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3342 VGND w_dly_sig[2] w_dly_sig_n[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3344 VGND a_14767_6549# o_result[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3345 VGND a_20395_10749# a_20566_10636# VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3348 a_14683_6575# a_13901_6581# a_14599_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3349 VPWR clknet_3_6__leaf_i_stop a_17507_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3350 VPWR i_stop a_16197_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3352 a_21909_10927# w_dly_sig[52] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3353 VPWR a_12115_8573# a_12283_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3354 a_13810_7663# a_13563_8041# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3355 w_dly_sig[33] w_dly_sig_n[32] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3356 clknet_3_3__leaf_i_stop a_14449_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3357 a_12149_11305# a_11159_10933# a_12023_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3358 VGND w_dly_sig_n[40] w_dly_sig[41] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3359 VPWR a_13679_8751# a_13847_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3363 w_dly_sig_n[61] w_dly_sig[61] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3367 w_dly_sig_n[8] w_dly_sig[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3370 VGND a_14691_12015# a_14859_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3371 a_22162_10901# a_21994_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3374 w_dly_sig[15] w_dly_sig_n[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3377 w_dly_sig[59] w_dly_sig_n[58] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3378 VPWR a_10138_10357# a_10067_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3380 a_14641_10927# w_dly_sig[56] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3381 w_dly_sig[46] w_dly_sig_n[45] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3382 VGND w_dly_sig_n[18] w_dly_sig[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3384 VGND a_16749_11445# clknet_3_6__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3385 a_13162_10927# a_12723_10933# a_13077_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3387 VPWR a_14817_7093# clknet_3_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3391 VGND w_dly_sig[51] w_dly_sig_n[51] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3392 a_15469_6031# w_dly_sig[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3394 VGND a_9389_11445# clknet_3_2__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3395 VGND w_dly_sig_n[35] w_dly_sig[36] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3400 w_dly_sig[51] w_dly_sig_n[50] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3401 w_dly_sig_n[19] w_dly_sig[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3402 VPWR a_22311_7637# o_result[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3403 w_dly_sig_n[48] w_dly_sig[48] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3404 a_9699_13481# a_9570_13225# a_9279_13335# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3405 a_8635_9269# a_8919_9269# a_8854_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3407 w_dly_sig_n[6] w_dly_sig[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3409 w_dly_sig[23] w_dly_sig_n[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3410 VPWR w_dly_sig[26] w_dly_sig_n[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3413 o_result[3] a_15503_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3415 o_result[30] a_8835_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3416 a_13763_8751# a_12981_8757# a_13679_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3417 VPWR a_14817_7093# clknet_3_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3421 a_12705_13103# a_12171_13109# a_12610_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3422 VGND a_14434_11989# a_14392_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3423 o_result[19] a_12835_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3424 VPWR clknet_0_i_stop a_9665_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3425 a_22086_10749# a_21813_10383# a_22001_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3427 VPWR w_dly_sig[21] w_dly_sig_n[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3428 VGND a_9665_7093# clknet_3_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3429 a_12688_10057# clknet_3_3__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3431 w_dly_sig[9] w_dly_sig_n[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3433 w_dly_sig_n[42] w_dly_sig[42] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3434 a_20119_12015# a_19421_12021# a_19862_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3435 VGND a_22311_8725# a_22269_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3437 clknet_3_6__leaf_i_stop a_16749_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3440 a_21822_11471# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3441 a_11246_9295# a_10859_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3442 w_dly_sig_n[2] w_dly_sig[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3443 w_dly_sig[49] w_dly_sig_n[48] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3444 VPWR clknet_3_1__leaf_i_stop a_15115_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3445 clknet_3_2__leaf_i_stop a_9389_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3446 VGND a_16854_8207# clknet_3_4__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3448 VPWR a_23063_12015# a_23231_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3451 VGND a_23063_12015# a_23231_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3452 a_18413_9839# w_dly_sig[45] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3453 a_21997_13109# a_21831_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3454 VPWR a_12023_11837# a_12191_11739# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3455 VPWR a_17102_10495# a_17029_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3457 VGND w_dly_sig_n[27] w_dly_sig[28] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3459 VPWR w_dly_sig[24] w_dly_sig_n[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3465 VGND a_18999_7637# o_result[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3466 o_result[59] a_20287_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3471 VGND clknet_3_7__leaf_i_stop a_22015_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3472 VPWR a_16854_8207# clknet_3_4__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3474 a_18915_7663# a_18133_7669# a_18831_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3475 o_result[59] a_20287_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3477 clknet_3_5__leaf_i_stop a_21822_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3480 VPWR a_12778_13077# a_12705_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3481 a_21445_8757# a_21279_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3482 a_13143_7895# a_13434_7785# a_13385_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3483 VPWR a_16807_12925# a_16975_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3484 o_result[41] a_17159_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3488 a_12429_12021# a_12263_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3489 a_23063_12015# a_22199_12021# a_22806_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3490 VPWR a_9011_8181# a_9018_8481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3491 a_17861_10927# w_dly_sig[54] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3493 a_22806_9407# a_22638_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3495 VPWR w_dly_sig[17] w_dly_sig_n[17] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3496 clknet_3_0__leaf_i_stop a_9665_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3497 VGND a_22806_11989# a_22764_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3498 clknet_0_i_stop a_16197_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3499 w_dly_sig[27] w_dly_sig_n[26] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3500 a_22806_9407# a_22638_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3501 a_21633_7663# w_dly_sig[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3502 a_18225_9845# a_18059_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3503 a_11513_11471# w_dly_sig[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3504 net1 a_855_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3506 a_20203_12015# a_19421_12021# a_20119_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3507 VPWR w_dly_sig[33] w_dly_sig_n[33] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3508 VPWR a_16749_11445# clknet_3_6__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3509 a_20598_11583# a_20430_11837# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3510 VGND a_20855_11837# a_21023_11739# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3513 a_13634_7940# a_13434_7785# a_13783_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3514 a_18869_8207# a_18703_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3515 a_22269_6953# a_21279_6581# a_22143_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3516 a_21886_7637# a_21718_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3517 a_17029_10749# a_16495_10383# a_16934_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3519 VGND a_9195_6005# a_9202_6305# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3523 a_14269_6575# a_13735_6581# a_14174_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3524 a_20295_9661# a_19513_9295# a_20211_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3526 w_dly_sig[34] w_dly_sig_n[33] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3527 o_result[28] a_8927_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3529 VPWR a_13203_13077# o_result[33] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3530 VGND clknet_3_3__leaf_i_stop a_13827_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3532 VGND a_13203_13077# o_result[33] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3533 o_result[44] a_19091_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3536 a_11325_11471# a_11159_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3539 a_22545_11305# a_21555_10933# a_22419_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3541 VGND w_dly_sig[63] w_dly_sig_n[63] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3543 VPWR w_dly_sig_n[48] w_dly_sig[49] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3547 a_9926_7637# a_9758_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3549 a_20479_10749# a_19697_10383# a_20395_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X3552 VGND w_dly_sig_n[7] w_dly_sig[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3554 a_22365_9295# a_22199_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3555 w_dly_sig[31] w_dly_sig_n[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3556 VGND a_8919_9269# a_8926_9569# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3557 a_9665_7093# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3560 o_result[27] a_9479_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3561 VPWR w_dly_sig_n[12] w_dly_sig[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3562 VGND a_9799_6549# o_result[22] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3563 VPWR a_12870_11989# a_12797_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3564 VPWR a_12975_7895# o_result[17] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3566 w_dly_sig_n[31] w_dly_sig[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3567 a_22120_11305# a_21721_10933# a_21994_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3568 o_result[41] a_17159_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3569 clknet_3_5__leaf_i_stop a_21822_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3570 VPWR a_9402_6005# a_9331_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3572 a_8835_12247# a_9003_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3573 a_13981_8041# a_13427_7881# a_13634_7940# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3575 a_16991_9661# a_16293_9295# a_16734_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3578 a_9762_10927# a_9515_11305# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3579 VGND a_14449_11445# clknet_3_3__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3585 a_13349_8751# a_12815_8757# a_13254_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3587 VGND a_21822_11471# clknet_3_7__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3589 VPWR a_16197_9813# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3590 a_19885_7663# w_dly_sig[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3593 a_13077_10927# w_dly_sig[38] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3595 o_result[9] a_22955_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3596 VGND w_dly_sig_n[6] w_dly_sig[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3597 VGND a_22438_13077# a_22396_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3600 VPWR clknet_0_i_stop a_14449_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3601 VPWR a_8559_8181# o_result[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3602 w_dly_sig[42] w_dly_sig_n[41] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3603 clknet_3_4__leaf_i_stop a_16854_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3604 VPWR w_dly_sig[6] w_dly_sig_n[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3605 a_22695_13103# a_21997_13109# a_22438_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3606 a_11325_10933# a_11159_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3607 a_20211_10927# a_19347_10933# a_19954_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3608 a_11027_9269# a_11311_9269# a_11246_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3613 w_dly_sig_n[54] w_dly_sig[54] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3615 a_18298_8725# a_18130_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3618 VGND a_21822_8207# clknet_3_5__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3620 a_18114_10901# a_17946_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3622 a_12242_6575# a_11803_6581# a_12157_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3625 VPWR a_15078_8725# a_15005_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3627 a_9218_8181# a_9011_8181# a_9394_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3628 a_22254_10495# a_22086_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3629 a_8877_9661# a_8467_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3630 VPWR w_dly_sig_n[8] w_dly_sig[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3632 clknet_3_7__leaf_i_stop a_21822_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3634 a_9586_11204# a_9379_11145# a_9762_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3635 a_9889_10749# a_9479_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3638 VGND a_14817_7093# clknet_3_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3639 VPWR a_9665_7093# clknet_3_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3641 VGND w_dly_sig[7] w_dly_sig_n[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3642 VGND a_9389_11445# clknet_3_2__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3643 a_9515_11305# a_9379_11145# a_9095_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3644 VPWR clknet_3_7__leaf_i_stop a_21555_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3647 a_18298_8725# a_18130_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3650 a_9479_10357# a_9647_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3651 VGND a_19735_8475# o_result[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3652 a_9758_7663# a_9319_7669# a_9673_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3656 VGND a_13847_8725# o_result[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3658 VGND clknet_3_3__leaf_i_stop a_12723_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3662 VGND a_9011_8181# a_9018_8481# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3663 w_dly_sig_n[29] w_dly_sig[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3666 o_result[10] a_22955_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3667 a_19693_8207# a_18703_8207# a_19567_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3668 a_9423_12393# a_9294_12137# a_9003_12247# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3674 a_9394_8573# a_9147_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3677 VPWR w_dly_sig_n[45] w_dly_sig[46] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3678 a_19786_9661# a_19513_9295# a_19701_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3679 VGND a_15503_8725# a_15461_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3681 VPWR w_dly_sig[15] w_dly_sig_n[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3682 a_16842_7663# a_16569_7669# a_16757_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3683 a_12368_6953# a_11969_6581# a_12242_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3685 a_16849_10383# w_dly_sig[55] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3689 VPWR w_dly_sig_n[24] w_dly_sig[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3692 a_22879_9839# a_22181_9845# a_22622_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3693 a_22454_9839# a_22015_9845# a_22369_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3694 w_dly_sig_n[26] w_dly_sig[26] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3696 VPWR w_dly_sig[48] w_dly_sig_n[48] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3699 VPWR a_18555_8751# a_18723_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3701 VPWR a_20566_10636# o_result[45] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X3702 VPWR clknet_0_i_stop a_16854_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3703 a_12023_11837# a_11325_11471# a_11766_11583# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3704 a_21718_6575# a_21445_6581# a_21633_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3705 VGND a_22311_6549# o_result[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3706 VGND a_20195_6549# o_result[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3707 a_11969_6581# a_11803_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3708 VGND w_dly_sig[58] w_dly_sig_n[58] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3709 w_dly_sig[28] w_dly_sig_n[27] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3710 a_9884_8041# a_9485_7669# a_9758_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3713 VPWR w_dly_sig_n[56] w_dly_sig[57] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3714 VPWR a_20119_12015# a_20287_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3715 VPWR clknet_3_4__leaf_i_stop a_17967_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3716 a_14637_8757# a_14471_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3719 VGND a_20119_12015# a_20287_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3721 a_10497_6031# a_10331_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3722 VGND w_dly_sig[10] w_dly_sig_n[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3727 VPWR a_12191_11739# o_result[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3730 a_9287_12233# clknet_3_2__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3732 clknet_3_1__leaf_i_stop a_14817_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3733 clknet_3_0__leaf_i_stop a_9665_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3735 w_dly_sig_n[24] w_dly_sig[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3736 a_16197_9813# i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3739 VGND w_dly_sig_n[59] w_dly_sig[60] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3742 VPWR w_dly_sig_n[11] w_dly_sig[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3744 o_result[40] a_14767_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3746 VPWR a_17159_11989# o_result[56] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3747 w_dly_sig_n[62] w_dly_sig[62] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3748 a_19310_8319# a_19142_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3751 VGND a_17159_11989# o_result[56] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3753 a_15078_7637# a_14910_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3754 a_18298_11989# a_18130_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3755 a_20119_12015# a_19255_12021# a_19862_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3756 a_17577_6953# a_16587_6581# a_17451_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3757 clknet_3_1__leaf_i_stop a_14817_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3759 w_dly_sig_n[64] w_dly_sig[64] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3760 VGND clknet_0_i_stop a_14449_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3761 w_dly_sig[25] w_dly_sig_n[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3763 VGND w_dly_sig[56] w_dly_sig_n[56] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3764 VPWR a_22679_10651# a_22595_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3765 VGND a_17159_8725# a_17117_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3769 VPWR a_16749_11445# clknet_3_6__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3770 VGND a_20566_10636# a_20524_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X3771 VGND w_dly_sig_n[17] w_dly_sig[18] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3772 VPWR clknet_0_i_stop a_21822_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3775 w_dly_sig[35] w_dly_sig_n[34] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3776 VPWR a_9389_11445# clknet_3_2__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3777 o_result[9] a_22955_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3778 o_result[33] a_13203_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3780 VGND a_22955_7387# a_22913_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3781 a_17060_10383# a_16661_10383# a_16934_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3782 a_22277_6031# w_dly_sig[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3784 o_result[33] a_13203_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3785 a_12400_9813# a_12698_9961# a_12646_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0913 ps=0.855 w=0.42 l=0.15
X3786 w_dly_sig[17] w_dly_sig_n[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3787 a_21721_10933# a_21555_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3788 VGND w_dly_sig_n[42] w_dly_sig[43] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3790 w_dly_sig_n[5] w_dly_sig[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3793 a_23189_9295# a_22199_9295# a_23063_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3794 a_19789_13109# a_19623_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3795 a_9565_8207# a_9018_8481# a_9218_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3796 w_dly_sig[21] w_dly_sig_n[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3799 VPWR a_19954_9407# a_19881_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3802 VPWR a_20230_13077# a_20157_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3803 a_16293_8757# a_16127_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3805 VPWR a_22143_7663# a_22311_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3807 a_9515_11305# a_9386_11049# a_9095_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3808 VGND a_20211_10927# a_20379_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3809 a_18498_9839# a_18225_9845# a_18413_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3813 a_16734_8725# a_16566_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3815 a_13119_13103# a_12337_13109# a_13035_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3817 clknet_3_4__leaf_i_stop a_16854_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3820 a_11598_11837# a_11159_11471# a_11513_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3821 VPWR w_dly_sig[60] w_dly_sig_n[60] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3823 VPWR a_21886_6549# a_21813_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3824 a_8919_9269# clknet_3_0__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3825 a_18639_12015# a_17857_12021# a_18555_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3828 VGND a_21822_11471# clknet_3_7__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3829 VPWR a_16197_9813# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3830 clknet_3_5__leaf_i_stop a_21822_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3832 a_11471_12925# a_10773_12559# a_11214_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3833 VPWR a_20855_11837# a_21023_11739# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3834 VPWR a_11363_6299# o_result[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3835 a_13127_12015# a_12429_12021# a_12870_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3836 a_21886_8725# a_21718_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3837 o_result[10] a_22955_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3838 w_dly_sig_n[36] w_dly_sig[36] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3839 VPWR a_14449_11445# clknet_3_3__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3840 VPWR a_10183_7663# a_10351_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3841 VGND a_22955_6299# a_22913_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3842 VGND a_16975_12827# o_result[57] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3843 a_9203_10071# a_9371_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3844 VPWR w_dly_sig_n[39] w_dly_sig[40] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3845 a_19881_9661# a_19347_9295# a_19786_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3846 clknet_3_4__leaf_i_stop a_16854_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3848 a_14453_10933# a_14287_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3849 VGND a_21822_8207# clknet_3_5__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3850 a_13563_8041# a_13434_7785# a_13143_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3851 a_16566_9661# a_16127_9295# a_16481_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3853 VGND i_stop a_16197_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3858 a_12892_10116# a_12698_9961# a_13068_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.0687 ps=0.76 w=0.36 l=0.15
X3860 VPWR w_dly_sig_n[53] w_dly_sig[54] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3861 VGND a_18831_7663# a_18999_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3864 w_dly_sig[64] w_dly_sig_n[63] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3865 o_result[36] a_13295_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3866 clknet_3_7__leaf_i_stop a_21822_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3867 w_dly_sig[5] w_dly_sig_n[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3868 a_21813_6575# a_21279_6581# a_21718_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3869 a_11321_6031# a_10331_6031# a_11195_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3870 a_19517_6575# w_dly_sig[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3872 o_result[1] a_12283_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3873 VGND a_9389_11445# clknet_3_2__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3877 VPWR a_17159_8725# o_result[42] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3878 a_19513_10933# a_19347_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3882 VPWR clknet_3_4__leaf_i_stop a_16403_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3883 a_9757_6953# a_8767_6581# a_9631_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3884 VGND a_10351_7637# o_result[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3885 a_19862_11989# a_19694_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3887 w_dly_sig_n[9] w_dly_sig[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3888 o_result[17] a_12975_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3889 VPWR a_13330_10901# a_13257_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3890 w_dly_sig_n[52] w_dly_sig[52] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3891 o_result[7] a_20563_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3892 w_dly_sig_n[30] w_dly_sig[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3893 a_19694_12015# a_19421_12021# a_19609_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3894 o_result[39] a_12050_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X3896 a_13211_12015# a_12429_12021# a_13127_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3897 VGND w_dly_sig[55] w_dly_sig_n[55] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3899 a_11214_12671# a_11046_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3900 VGND a_8927_11159# o_result[28] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3901 VPWR w_dly_sig[1] w_dly_sig_n[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3902 o_result[50] a_22679_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3903 a_16692_9295# a_16293_9295# a_16566_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3905 w_dly_sig_n[12] w_dly_sig[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3906 a_12525_13103# w_dly_sig[34] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3908 a_19329_6581# a_19163_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3909 a_9485_7669# a_9319_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3912 VGND a_16749_11445# clknet_3_6__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3913 VGND a_23231_9563# o_result[48] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3915 a_11724_11305# a_11325_10933# a_11598_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3918 VPWR a_18666_9813# a_18593_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3922 a_8467_9269# a_8635_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3926 a_18413_9839# w_dly_sig[45] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3927 a_19977_13103# w_dly_sig[62] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3929 a_17026_6575# a_16753_6581# a_16941_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3931 VPWR clknet_0_i_stop a_16749_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3932 VGND w_dly_sig_n[0] w_dly_sig[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3936 a_14691_12015# a_13827_12021# a_14434_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3937 o_result[45] a_20566_10636# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X3940 a_12702_12015# a_12263_12021# a_12617_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3941 a_19057_8207# w_dly_sig[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3943 a_14361_12015# a_13827_12021# a_14266_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3944 VPWR w_dly_sig_n[2] w_dly_sig[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3945 VGND a_13422_8725# a_13380_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3946 w_dly_sig[57] w_dly_sig_n[56] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3948 a_10938_6143# a_10770_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3950 VPWR a_21822_11471# clknet_3_7__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3952 VGND a_23231_9563# a_23189_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3953 VPWR a_18539_10901# a_18455_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3954 VPWR w_dly_sig[25] w_dly_sig_n[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3955 a_15078_7637# a_14910_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3959 VGND a_9631_6575# a_9799_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3960 a_20981_11471# a_19991_11471# a_20855_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3964 a_14725_6953# a_13735_6581# a_14599_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3965 o_result[5] a_17435_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3966 w_dly_sig_n[34] w_dly_sig[34] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3967 w_dly_sig_n[40] w_dly_sig[40] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3970 VGND a_16734_9407# a_16692_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3971 a_22143_8751# a_21445_8757# a_21886_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3974 o_result[40] a_14767_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3976 VPWR w_dly_sig_n[16] w_dly_sig[17] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3978 a_18593_9839# a_18059_9845# a_18498_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3980 VPWR w_dly_sig_n[60] w_dly_sig[61] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3982 w_dly_sig[60] w_dly_sig_n[59] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3983 VGND w_dly_sig_n[1] w_dly_sig[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3984 VPWR a_19567_8573# a_19735_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3987 w_dly_sig_n[35] w_dly_sig[35] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3988 VGND w_dly_sig_n[39] w_dly_sig[40] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3991 a_13427_7881# clknet_3_1__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3992 w_dly_sig_n[57] w_dly_sig[57] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3993 w_dly_sig_n[4] w_dly_sig[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3997 w_dly_sig_n[56] w_dly_sig[56] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3998 a_22143_8751# a_21279_8757# a_21886_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4001 VPWR a_14434_11989# a_14361_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4002 VGND a_13679_8751# a_13847_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4004 VPWR i_start a_855_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4009 clknet_3_3__leaf_i_stop a_14449_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4010 a_15469_6031# w_dly_sig[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4012 VGND a_14618_12671# a_14576_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4013 a_12050_9813# a_12400_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.106 ps=0.975 w=0.65 l=0.15
X4015 VPWR w_dly_sig[31] a_9841_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4016 a_22733_12015# a_22199_12021# a_22638_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4017 VGND a_13755_10901# a_13713_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4018 VGND w_dly_sig_n[37] w_dly_sig[38] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4019 VPWR clknet_3_7__leaf_i_stop a_19531_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4020 w_dly_sig[1] w_dly_sig_n[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4021 o_result[11] a_22311_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4026 VGND a_9586_11204# a_9515_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4027 a_13074_9839# a_12821_10217# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.179 ps=1.26 w=0.42 l=0.15
X4028 w_dly_sig_n[47] w_dly_sig[47] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4030 a_22143_7663# a_21445_7669# a_21886_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4034 VGND a_18574_7637# a_18532_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4035 VPWR a_15335_7663# a_15503_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4037 w_dly_sig_n[53] w_dly_sig[53] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4040 VGND w_dly_sig_n[3] w_dly_sig[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4043 a_14875_12925# a_14011_12559# a_14618_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4044 VGND a_17527_10651# a_17485_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4045 a_17351_7663# a_16569_7669# a_17267_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4046 a_12070_7940# a_11870_7785# a_12219_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4048 w_dly_sig[36] w_dly_sig_n[35] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4049 o_result[3] a_15503_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4050 a_14545_12925# a_14011_12559# a_14450_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4051 VGND a_21822_11471# clknet_3_7__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4053 VGND clknet_0_i_stop a_9389_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4054 VGND a_21822_11471# clknet_3_7__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4055 a_10067_10383# a_9938_10657# a_9647_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4057 a_10183_7663# a_9485_7669# a_9926_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4058 o_result[26] a_9203_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4061 o_result[15] a_16147_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4063 a_9841_12393# a_9287_12233# a_9494_12292# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4064 VPWR a_22806_11989# a_22733_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4065 a_22227_6575# a_21445_6581# a_22143_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4066 VGND clknet_0_i_stop a_9665_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4071 a_13169_8751# w_dly_sig[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4073 VGND a_21822_8207# clknet_3_5__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4076 VPWR w_dly_sig[9] w_dly_sig_n[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4077 VGND a_9203_10071# o_result[26] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4078 VGND a_12688_10057# a_12698_9961# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4079 VGND clknet_3_3__leaf_i_stop a_14287_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4080 VGND a_16197_9813# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4082 VGND a_16197_9813# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4085 a_22185_13103# w_dly_sig[63] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4088 VGND a_14817_7093# clknet_3_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4089 VPWR clknet_0_i_stop a_14817_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4090 VPWR a_9665_7093# clknet_3_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4091 VPWR a_20138_7637# a_20065_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4092 a_11311_9269# clknet_3_3__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4093 a_16481_9295# w_dly_sig[42] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4094 VGND clknet_3_1__leaf_i_stop a_12815_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4096 VPWR i_stop a_16197_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4099 w_dly_sig[45] w_dly_sig_n[44] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4101 w_dly_sig[8] w_dly_sig_n[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4105 o_result[49] a_23047_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4106 w_dly_sig_n[22] w_dly_sig[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4108 VPWR a_14618_12671# a_14545_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4109 clknet_3_6__leaf_i_stop a_16749_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4110 a_12417_8041# a_11863_7881# a_12070_7940# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4111 VPWR w_dly_sig[59] w_dly_sig_n[59] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4114 VGND a_16854_8207# clknet_3_4__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4116 w_dly_sig_n[32] w_dly_sig[32] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4117 VGND w_dly_sig[1] a_11865_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4118 a_19954_9407# a_19786_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4121 a_12646_9839# a_12050_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.122 ps=1.42 w=0.42 l=0.15
X4122 a_18639_8751# a_17857_8757# a_18555_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4123 VPWR a_22311_8725# a_22227_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4128 w_dly_sig[19] w_dly_sig_n[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4129 VPWR clknet_3_7__leaf_i_stop a_19347_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4130 a_8467_9269# a_8635_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4131 VGND a_23231_11989# o_result[63] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4132 a_19970_7663# a_19697_7669# a_19885_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4134 a_22871_6397# a_22089_6031# a_22787_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4139 VGND clknet_3_3__leaf_i_stop a_12263_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4141 VGND w_dly_sig[20] w_dly_sig_n[20] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4143 VPWR w_dly_sig[25] a_9565_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4145 a_13127_12015# a_12263_12021# a_12870_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4146 a_20065_7663# a_19531_7669# a_19970_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4147 clknet_3_7__leaf_i_stop a_21822_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4148 a_17946_10927# a_17673_10933# a_17861_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4149 VPWR w_dly_sig_n[46] w_dly_sig[47] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4150 VGND a_12870_11989# a_12828_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4151 VGND a_16749_11445# clknet_3_6__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4152 a_14852_11305# a_14453_10933# a_14726_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4153 a_11690_8573# a_11251_8207# a_11605_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4154 VPWR a_16975_12827# o_result[57] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4155 VGND a_16749_11445# clknet_3_6__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4156 a_11863_7881# clknet_3_1__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4157 w_dly_sig_n[33] w_dly_sig[33] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4160 VGND w_dly_sig[49] w_dly_sig_n[49] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4164 a_19609_12015# w_dly_sig[60] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4167 a_9222_12381# a_8835_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4169 VPWR w_dly_sig[14] w_dly_sig_n[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4170 a_22419_10927# a_21721_10933# a_22162_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4174 clknet_3_2__leaf_i_stop a_9389_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4177 a_20062_13103# a_19623_13109# a_19977_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4179 a_13362_8029# a_12975_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4182 a_16849_10383# w_dly_sig[55] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4183 VGND a_18923_9839# a_19091_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4185 VPWR a_11195_6397# a_11363_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4187 o_result[32] a_11639_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4189 a_14392_12393# a_13993_12021# a_14266_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4190 VPWR clknet_3_2__leaf_i_stop a_11159_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4191 VGND a_21023_11739# o_result[60] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4194 VPWR w_dly_sig_n[47] w_dly_sig[48] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4195 VPWR a_23063_9661# a_23231_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4196 VPWR w_dly_sig[4] w_dly_sig_n[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4197 w_dly_sig_n[7] w_dly_sig[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4199 VPWR a_21822_11471# clknet_3_7__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4200 w_dly_sig_n[63] w_dly_sig[63] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4202 a_16197_9813# i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4204 a_16293_12021# a_16127_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4205 clknet_3_2__leaf_i_stop a_9389_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4206 a_19979_10749# a_19697_10383# a_19885_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X4207 a_15335_8751# a_14637_8757# a_15078_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4208 VGND w_dly_sig_n[21] w_dly_sig[22] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4210 a_10011_10205# a_9791_10217# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X4212 VGND a_20379_10901# a_20337_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4213 VPWR clknet_3_7__leaf_i_stop a_22015_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4214 VGND a_22143_7663# a_22311_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4215 w_dly_sig_n[45] w_dly_sig[45] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4216 VPWR a_16854_8207# clknet_3_4__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X4217 clknet_3_4__leaf_i_stop a_16854_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4218 a_9933_11305# a_9379_11145# a_9586_11204# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4220 a_14342_9813# a_14174_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4221 a_11816_8207# a_11417_8207# a_11690_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4223 VPWR w_dly_sig_n[23] w_dly_sig[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4225 VGND a_21886_6549# a_21844_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4229 w_dly_sig[61] w_dly_sig_n[60] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4230 a_8559_8181# a_8727_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4232 VPWR w_dly_sig_n[64] g_dly_chain_even[64].dly_stg2.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4233 o_result[50] a_22679_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4235 a_12149_11471# a_11159_11471# a_12023_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4237 clknet_3_1__leaf_i_stop a_14817_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4241 VPWR w_dly_sig[3] w_dly_sig_n[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4242 VPWR a_16991_8751# a_17159_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4246 a_15335_8751# a_14471_8757# a_15078_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4248 VPWR clknet_3_6__leaf_i_stop a_17691_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4249 a_9479_10357# a_9647_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4250 VGND a_10975_8759# _64_.X VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X4252 VGND a_10183_7663# a_10351_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4253 w_dly_sig[42] w_dly_sig_n[41] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4256 a_11667_9295# a_11447_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X4257 w_dly_sig_n[14] w_dly_sig[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4259 a_16807_12925# a_16109_12559# a_16550_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4263 w_dly_sig[24] w_dly_sig_n[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4265 a_22764_12393# a_22365_12021# a_22638_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4266 a_19701_10927# w_dly_sig[53] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4268 VPWR w_dly_sig[28] w_dly_sig_n[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4271 a_10267_7663# a_9485_7669# a_10183_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4273 o_result[14] a_17619_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4274 VGND w_dly_sig[18] w_dly_sig_n[18] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4275 VGND clknet_3_2__leaf_i_stop a_11159_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4276 a_9655_10057# clknet_3_2__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4278 a_12610_13103# a_12171_13109# a_12525_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4279 VPWR a_22162_10901# a_22089_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4282 a_15335_7663# a_14637_7669# a_15078_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4283 a_15151_10927# a_14287_10933# a_14894_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4284 w_dly_sig_n[10] w_dly_sig[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4287 VGND a_11766_10901# a_11724_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4288 a_22622_9813# a_22454_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4289 VGND a_23063_9661# a_23231_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4290 VGND a_11858_8319# a_11816_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4294 VPWR w_dly_sig[37] w_dly_sig_n[37] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4295 clknet_0_i_stop a_16197_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4298 VPWR w_dly_sig_n[32] w_dly_sig[33] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4300 o_result[25] a_8467_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4302 a_19513_9295# a_19347_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4303 a_12115_8573# a_11417_8207# a_11858_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4306 VPWR a_14599_9839# a_14767_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4307 a_22457_6397# a_21923_6031# a_22362_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4308 o_result[35] a_14859_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4309 VGND clknet_0_i_stop a_21822_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4310 VGND w_dly_sig[29] a_9933_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4311 VPWR w_dly_sig_n[15] w_dly_sig[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4313 o_result[7] a_20563_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4315 a_9111_13335# a_9279_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4316 a_9003_12247# a_9287_12233# a_9222_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4317 o_result[35] a_14859_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4319 VPWR w_dly_sig[27] a_10209_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4323 VGND a_22679_10651# o_result[50] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4324 a_19651_8573# a_18869_8207# a_19567_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4326 a_11518_9269# a_11318_9569# a_11667_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4327 VPWR a_9126_9269# a_9055_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4328 VGND clknet_0_i_stop a_21822_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4333 a_17443_10749# a_16661_10383# a_17359_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4334 a_14449_11445# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4335 a_18321_7663# w_dly_sig[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4336 a_21445_8757# a_21279_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4337 VPWR a_20566_10636# o_result[45] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4340 VGND a_16197_9813# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4341 VGND w_dly_sig_n[50] w_dly_sig[51] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4342 _64_.X a_10975_8759# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X4344 VGND a_18555_8751# a_18723_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4349 VGND a_21822_8207# clknet_3_5__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4350 VPWR clknet_3_5__leaf_i_stop a_19531_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4352 VGND a_8835_12247# o_result[30] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4355 VGND w_dly_sig_n[13] w_dly_sig[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4357 VGND i_start a_855_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4359 a_16481_12015# w_dly_sig[57] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4360 a_13262_10217# a_12688_10057# a_12892_10116# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X4362 a_21633_6575# w_dly_sig[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4364 a_16382_12925# a_16109_12559# a_16297_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4365 a_22622_9813# a_22454_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4367 clknet_3_6__leaf_i_stop a_16749_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X4369 a_13262_10217# a_12698_9961# a_12892_10116# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0662 ps=0.735 w=0.42 l=0.15
X4370 a_15554_6397# a_15115_6031# a_15469_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4371 VGND w_dly_sig[42] w_dly_sig_n[42] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4373 a_11597_12559# a_10607_12559# a_11471_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4374 VPWR a_15503_8725# a_15419_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4376 a_13288_11305# a_12889_10933# a_13162_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4377 VGND w_dly_sig[41] w_dly_sig_n[41] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4379 VPWR clknet_3_4__leaf_i_stop a_16587_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4380 a_11865_9295# a_11311_9269# a_11518_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4381 o_result[63] a_23231_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4383 o_result[63] a_23231_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4385 w_dly_sig[16] w_dly_sig_n[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4387 w_dly_sig_n[50] w_dly_sig[50] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4388 VPWR w_dly_sig[19] a_12417_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4389 VPWR a_9287_12233# a_9294_12137# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4390 w_dly_sig[50] w_dly_sig_n[49] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4393 VGND a_21886_7637# a_21844_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4394 w_dly_sig[39] w_dly_sig_n[38] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4395 clknet_3_7__leaf_i_stop a_21822_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4396 VPWR w_dly_sig_n[44] w_dly_sig[45] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4397 VPWR w_dly_sig_n[29] w_dly_sig[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4398 w_dly_sig[11] w_dly_sig_n[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4399 VPWR a_20287_11989# o_result[59] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4400 clknet_3_7__leaf_i_stop a_21822_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4403 a_9791_10217# a_9662_9961# a_9371_10071# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4404 a_19697_6575# a_19163_6581# a_19602_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4405 VGND a_20287_11989# o_result[59] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4409 clknet_3_1__leaf_i_stop a_14817_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4411 o_result[57] a_16975_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4412 a_12023_11837# a_11159_11471# a_11766_11583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4414 VPWR a_9218_8181# a_9147_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4415 a_11605_8207# w_dly_sig[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4416 o_result[17] a_12975_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4417 a_23147_12015# a_22365_12021# a_23063_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4418 a_9673_7663# w_dly_sig[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4419 a_11693_11837# a_11159_11471# a_11598_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4420 a_19885_10383# w_dly_sig[46] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X4421 a_15680_6031# a_15281_6031# a_15554_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4424 a_13068_10205# a_12821_10217# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.149 ps=1.22 w=0.42 l=0.15
X4426 a_17946_10927# a_17507_10933# a_17861_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4428 VPWR clknet_3_3__leaf_i_stop a_12171_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4429 a_22001_10383# w_dly_sig[51] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4432 o_result[37] a_13755_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4434 VPWR a_13035_13103# a_13203_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4435 VGND a_13035_13103# a_13203_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4436 VPWR a_21822_11471# clknet_3_7__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4438 o_result[60] a_21023_11739# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4439 o_result[11] a_22311_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4440 a_20138_10519# a_19979_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4441 VGND net1 w_dly_sig_n[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4445 clknet_3_2__leaf_i_stop a_9389_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4446 a_9095_11159# a_9379_11145# a_9314_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4448 VPWR clknet_3_6__leaf_i_stop a_16127_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4449 a_9665_7093# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4450 VGND a_15335_7663# a_15503_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4451 VGND w_dly_sig_n[33] w_dly_sig[34] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4452 a_8854_9295# a_8467_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4454 a_9715_6575# a_8933_6581# a_9631_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4455 clknet_3_5__leaf_i_stop a_21822_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4461 VPWR a_10859_9269# o_result[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4462 VPWR w_dly_sig_n[25] w_dly_sig[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4463 VGND w_dly_sig[43] w_dly_sig_n[43] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4466 w_dly_sig_n[16] w_dly_sig[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4468 a_13035_13103# a_12171_13109# a_12778_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4469 VPWR a_11766_11583# a_11693_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4470 VGND a_15151_10927# a_15319_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4472 a_14817_7093# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4473 a_14618_12671# a_14450_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4474 a_19237_8573# a_18703_8207# a_19142_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4475 o_result[18] a_11411_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4477 g_dly_chain_even[64].dly_stg2.Y w_dly_sig_n[64] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4478 VPWR a_22511_10749# a_22679_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4480 VGND w_dly_sig[32] a_10117_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4481 VGND a_14875_12925# a_15043_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4482 clknet_3_2__leaf_i_stop a_9389_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4483 a_11518_9269# a_11311_9269# a_11694_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4486 w_dly_sig[20] w_dly_sig_n[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4489 VGND w_dly_sig_n[30] w_dly_sig[31] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4490 o_result[25] a_8467_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4491 clknet_3_4__leaf_i_stop a_16854_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4493 VGND clknet_3_6__leaf_i_stop a_16127_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4494 VGND a_20211_9661# a_20379_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4495 w_dly_sig_n[49] w_dly_sig[49] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4496 o_result[52] a_20379_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4498 a_21909_10927# w_dly_sig[52] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4502 VPWR a_16197_9813# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 o_result[10] VGND 4.35f
C1 o_result[15] VGND 3.21f
C2 o_result[20] VGND 2.75f
C3 o_result[21] VGND 2.84f
C4 o_result[11] VGND 4.57f
C5 o_result[12] VGND 3.85f
C6 o_result[14] VGND 3.35f
C7 o_result[16] VGND 3.15f
C8 o_result[19] VGND 3.05f
C9 o_result[22] VGND 3.13f
C10 o_result[9] VGND 4.17f
C11 o_result[8] VGND 4.73f
C12 o_result[7] VGND 3.79f
C13 o_result[13] VGND 3.76f
C14 o_result[5] VGND 4.68f
C15 o_result[4] VGND 3.75f
C16 o_result[17] VGND 3.59f
C17 o_result[18] VGND 3.88f
C18 o_result[23] VGND 3.47f
C19 o_result[6] VGND 3.94f
C20 o_result[1] VGND 3.83f
C21 o_result[24] VGND 4.23f
C22 o_result[47] VGND 4.4f
C23 o_result[43] VGND 4.71f
C24 o_result[42] VGND 4.15f
C25 o_result[3] VGND 4.25f
C26 o_result[2] VGND 3.77f
C27 i_start VGND 0.9f
C28 o_result[48] VGND 4.56f
C29 o_result[46] VGND 5.32f
C30 o_result[41] VGND 4.8f
C31 o_result[0] VGND 5.24f
C32 o_result[25] VGND 4.08f
C33 o_result[49] VGND 4.21f
C34 o_result[44] VGND 5.04f
C35 o_result[40] VGND 4.32f
C36 o_result[39] VGND 6.48f
C37 o_result[26] VGND 4.51f
C38 i_stop VGND 7.17f
C39 o_result[50] VGND 4.34f
C40 o_result[45] VGND 6.9f
C41 o_result[54] VGND 4.37f
C42 o_result[27] VGND 4.63f
C43 o_result[51] VGND 5.04f
C44 o_result[52] VGND 5.34f
C45 o_result[53] VGND 4.58f
C46 o_result[55] VGND 4.09f
C47 o_result[37] VGND 3.77f
C48 o_result[38] VGND 4.33f
C49 o_result[28] VGND 4.39f
C50 o_result[60] VGND 4.05f
C51 o_result[29] VGND 4.29f
C52 o_result[63] VGND 4.1f
C53 o_result[59] VGND 3.58f
C54 o_result[58] VGND 3.5f
C55 o_result[56] VGND 3.35f
C56 o_result[35] VGND 3.46f
C57 o_result[36] VGND 3.35f
C58 o_result[30] VGND 4.27f
C59 o_result[57] VGND 3.41f
C60 o_result[34] VGND 3.13f
C61 o_result[32] VGND 3.25f
C62 o_result[62] VGND 4.24f
C63 o_result[61] VGND 3.27f
C64 o_result[33] VGND 3.16f
C65 o_result[31] VGND 3.39f
C66 VPWR VGND 2.74p
C67 a_22277_6031# VGND 0.23f $ **FLOATING
C68 a_22787_6397# VGND 0.609f $ **FLOATING
C69 a_22955_6299# VGND 0.97f $ **FLOATING
C70 a_22362_6397# VGND 0.626f $ **FLOATING
C71 a_22530_6143# VGND 0.581f $ **FLOATING
C72 a_22089_6031# VGND 1.43f $ **FLOATING
C73 a_21923_6031# VGND 1.81f $ **FLOATING
C74 a_15469_6031# VGND 0.23f $ **FLOATING
C75 a_15979_6397# VGND 0.609f $ **FLOATING
C76 a_16147_6299# VGND 0.97f $ **FLOATING
C77 a_15554_6397# VGND 0.626f $ **FLOATING
C78 a_15722_6143# VGND 0.581f $ **FLOATING
C79 a_15281_6031# VGND 1.43f $ **FLOATING
C80 a_15115_6031# VGND 1.81f $ **FLOATING
C81 a_10685_6031# VGND 0.23f $ **FLOATING
C82 a_11195_6397# VGND 0.609f $ **FLOATING
C83 a_11363_6299# VGND 0.97f $ **FLOATING
C84 a_10770_6397# VGND 0.626f $ **FLOATING
C85 a_10938_6143# VGND 0.581f $ **FLOATING
C86 a_10497_6031# VGND 1.43f $ **FLOATING
C87 a_10331_6031# VGND 1.81f $ **FLOATING
C88 a_9749_6031# VGND 0.23f $ **FLOATING
C89 w_dly_sig[22] VGND 1.72f $ **FLOATING
C90 a_9331_6031# VGND 0.581f $ **FLOATING
C91 a_9402_6005# VGND 0.626f $ **FLOATING
C92 a_9195_6005# VGND 1.81f $ **FLOATING
C93 a_9202_6305# VGND 1.43f $ **FLOATING
C94 a_8911_6005# VGND 0.609f $ **FLOATING
C95 a_8743_6005# VGND 0.97f $ **FLOATING
C96 a_21633_6575# VGND 0.23f $ **FLOATING
C97 a_19517_6575# VGND 0.23f $ **FLOATING
C98 w_dly_sig_n[14] VGND 1.37f $ **FLOATING
C99 a_16941_6575# VGND 0.23f $ **FLOATING
C100 w_dly_sig_n[16] VGND 1.37f $ **FLOATING
C101 a_14089_6575# VGND 0.23f $ **FLOATING
C102 a_12157_6575# VGND 0.23f $ **FLOATING
C103 w_dly_sig_n[21] VGND 1.56f $ **FLOATING
C104 a_9121_6575# VGND 0.23f $ **FLOATING
C105 a_22143_6575# VGND 0.609f $ **FLOATING
C106 a_22311_6549# VGND 0.97f $ **FLOATING
C107 a_21718_6575# VGND 0.626f $ **FLOATING
C108 a_21886_6549# VGND 0.581f $ **FLOATING
C109 a_21445_6581# VGND 1.43f $ **FLOATING
C110 w_dly_sig[12] VGND 1.88f $ **FLOATING
C111 a_21279_6581# VGND 1.81f $ **FLOATING
C112 w_dly_sig_n[12] VGND 1.05f $ **FLOATING
C113 a_20027_6575# VGND 0.609f $ **FLOATING
C114 a_20195_6549# VGND 0.97f $ **FLOATING
C115 a_19602_6575# VGND 0.626f $ **FLOATING
C116 a_19770_6549# VGND 0.581f $ **FLOATING
C117 a_19329_6581# VGND 1.43f $ **FLOATING
C118 a_19163_6581# VGND 1.81f $ **FLOATING
C119 w_dly_sig[13] VGND 1.96f $ **FLOATING
C120 w_dly_sig_n[13] VGND 0.821f $ **FLOATING
C121 a_17451_6575# VGND 0.609f $ **FLOATING
C122 a_17619_6549# VGND 0.97f $ **FLOATING
C123 a_17026_6575# VGND 0.626f $ **FLOATING
C124 a_17194_6549# VGND 0.581f $ **FLOATING
C125 a_16753_6581# VGND 1.43f $ **FLOATING
C126 a_16587_6581# VGND 1.81f $ **FLOATING
C127 w_dly_sig[15] VGND 1.71f $ **FLOATING
C128 w_dly_sig_n[15] VGND 0.93f $ **FLOATING
C129 w_dly_sig[16] VGND 1.69f $ **FLOATING
C130 a_14599_6575# VGND 0.609f $ **FLOATING
C131 a_14767_6549# VGND 0.97f $ **FLOATING
C132 a_14174_6575# VGND 0.626f $ **FLOATING
C133 a_14342_6549# VGND 0.581f $ **FLOATING
C134 a_13901_6581# VGND 1.43f $ **FLOATING
C135 a_13735_6581# VGND 1.81f $ **FLOATING
C136 a_12667_6575# VGND 0.609f $ **FLOATING
C137 a_12835_6549# VGND 0.97f $ **FLOATING
C138 a_12242_6575# VGND 0.626f $ **FLOATING
C139 a_12410_6549# VGND 0.581f $ **FLOATING
C140 a_11969_6581# VGND 1.43f $ **FLOATING
C141 a_11803_6581# VGND 1.81f $ **FLOATING
C142 w_dly_sig_n[20] VGND 0.782f $ **FLOATING
C143 w_dly_sig[21] VGND 1.73f $ **FLOATING
C144 a_9631_6575# VGND 0.609f $ **FLOATING
C145 a_9799_6549# VGND 0.97f $ **FLOATING
C146 a_9206_6575# VGND 0.626f $ **FLOATING
C147 a_9374_6549# VGND 0.581f $ **FLOATING
C148 a_8933_6581# VGND 1.43f $ **FLOATING
C149 a_8767_6581# VGND 1.81f $ **FLOATING
C150 a_22277_7119# VGND 0.23f $ **FLOATING
C151 a_22787_7485# VGND 0.609f $ **FLOATING
C152 a_22955_7387# VGND 0.97f $ **FLOATING
C153 a_22362_7485# VGND 0.626f $ **FLOATING
C154 a_22530_7231# VGND 0.581f $ **FLOATING
C155 a_22089_7119# VGND 1.43f $ **FLOATING
C156 a_21923_7119# VGND 1.81f $ **FLOATING
C157 w_dly_sig_n[11] VGND 1.3f $ **FLOATING
C158 w_dly_sig[20] VGND 1.69f $ **FLOATING
C159 w_dly_sig_n[9] VGND 0.782f $ **FLOATING
C160 w_dly_sig[11] VGND 2.22f $ **FLOATING
C161 w_dly_sig_n[8] VGND 0.899f $ **FLOATING
C162 w_dly_sig_n[7] VGND 0.86f $ **FLOATING
C163 a_14817_7093# VGND 4.03f $ **FLOATING
C164 w_dly_sig[17] VGND 1.84f $ **FLOATING
C165 w_dly_sig_n[17] VGND 0.782f $ **FLOATING
C166 w_dly_sig_n[18] VGND 1.17f $ **FLOATING
C167 w_dly_sig_n[19] VGND 0.813f $ **FLOATING
C168 a_9665_7093# VGND 4.03f $ **FLOATING
C169 w_dly_sig_n[22] VGND 1.52f $ **FLOATING
C170 a_21633_7663# VGND 0.23f $ **FLOATING
C171 a_19885_7663# VGND 0.23f $ **FLOATING
C172 a_18321_7663# VGND 0.23f $ **FLOATING
C173 a_16757_7663# VGND 0.23f $ **FLOATING
C174 a_14825_7663# VGND 0.23f $ **FLOATING
C175 a_13981_8041# VGND 0.23f $ **FLOATING
C176 a_12417_8041# VGND 0.23f $ **FLOATING
C177 a_9673_7663# VGND 0.23f $ **FLOATING
C178 a_22143_7663# VGND 0.609f $ **FLOATING
C179 a_22311_7637# VGND 0.97f $ **FLOATING
C180 a_21718_7663# VGND 0.626f $ **FLOATING
C181 a_21886_7637# VGND 0.581f $ **FLOATING
C182 a_21445_7669# VGND 1.43f $ **FLOATING
C183 w_dly_sig[9] VGND 2.11f $ **FLOATING
C184 a_21279_7669# VGND 1.81f $ **FLOATING
C185 a_20395_7663# VGND 0.609f $ **FLOATING
C186 a_20563_7637# VGND 0.97f $ **FLOATING
C187 a_19970_7663# VGND 0.626f $ **FLOATING
C188 a_20138_7637# VGND 0.581f $ **FLOATING
C189 a_19697_7669# VGND 1.43f $ **FLOATING
C190 w_dly_sig[8] VGND 1.95f $ **FLOATING
C191 a_19531_7669# VGND 1.81f $ **FLOATING
C192 a_18831_7663# VGND 0.609f $ **FLOATING
C193 a_18999_7637# VGND 0.97f $ **FLOATING
C194 a_18406_7663# VGND 0.626f $ **FLOATING
C195 a_18574_7637# VGND 0.581f $ **FLOATING
C196 a_18133_7669# VGND 1.43f $ **FLOATING
C197 w_dly_sig[14] VGND 1.83f $ **FLOATING
C198 a_17967_7669# VGND 1.81f $ **FLOATING
C199 a_17267_7663# VGND 0.609f $ **FLOATING
C200 a_17435_7637# VGND 0.97f $ **FLOATING
C201 a_16842_7663# VGND 0.626f $ **FLOATING
C202 a_17010_7637# VGND 0.581f $ **FLOATING
C203 a_16569_7669# VGND 1.43f $ **FLOATING
C204 a_16403_7669# VGND 1.81f $ **FLOATING
C205 a_15335_7663# VGND 0.609f $ **FLOATING
C206 a_15503_7637# VGND 0.97f $ **FLOATING
C207 a_14910_7663# VGND 0.626f $ **FLOATING
C208 a_15078_7637# VGND 0.581f $ **FLOATING
C209 a_14637_7669# VGND 1.43f $ **FLOATING
C210 a_14471_7669# VGND 1.81f $ **FLOATING
C211 w_dly_sig[18] VGND 1.65f $ **FLOATING
C212 a_13563_8041# VGND 0.581f $ **FLOATING
C213 a_13634_7940# VGND 0.626f $ **FLOATING
C214 a_13434_7785# VGND 1.43f $ **FLOATING
C215 a_13427_7881# VGND 1.81f $ **FLOATING
C216 a_13143_7895# VGND 0.609f $ **FLOATING
C217 a_12975_7895# VGND 0.97f $ **FLOATING
C218 w_dly_sig[19] VGND 1.88f $ **FLOATING
C219 a_11999_8041# VGND 0.581f $ **FLOATING
C220 a_12070_7940# VGND 0.626f $ **FLOATING
C221 a_11870_7785# VGND 1.43f $ **FLOATING
C222 a_11863_7881# VGND 1.81f $ **FLOATING
C223 a_11579_7895# VGND 0.609f $ **FLOATING
C224 a_11411_7895# VGND 0.97f $ **FLOATING
C225 a_10183_7663# VGND 0.609f $ **FLOATING
C226 a_10351_7637# VGND 0.97f $ **FLOATING
C227 a_9758_7663# VGND 0.626f $ **FLOATING
C228 a_9926_7637# VGND 0.581f $ **FLOATING
C229 a_9485_7669# VGND 1.43f $ **FLOATING
C230 a_9319_7669# VGND 1.81f $ **FLOATING
C231 w_dly_sig_n[23] VGND 0.813f $ **FLOATING
C232 w_dly_sig[23] VGND 2.13f $ **FLOATING
C233 w_dly_sig_n[10] VGND 1.34f $ **FLOATING
C234 a_19057_8207# VGND 0.23f $ **FLOATING
C235 a_21822_8207# VGND 4.03f $ **FLOATING
C236 w_dly_sig[10] VGND 1.94f $ **FLOATING
C237 a_19567_8573# VGND 0.609f $ **FLOATING
C238 a_19735_8475# VGND 0.97f $ **FLOATING
C239 a_19142_8573# VGND 0.626f $ **FLOATING
C240 a_19310_8319# VGND 0.581f $ **FLOATING
C241 a_18869_8207# VGND 1.43f $ **FLOATING
C242 w_dly_sig[7] VGND 2.21f $ **FLOATING
C243 a_18703_8207# VGND 1.81f $ **FLOATING
C244 w_dly_sig_n[6] VGND 1.81f $ **FLOATING
C245 w_dly_sig_n[5] VGND 1.15f $ **FLOATING
C246 a_11605_8207# VGND 0.23f $ **FLOATING
C247 a_16854_8207# VGND 4.03f $ **FLOATING
C248 w_dly_sig[6] VGND 1.58f $ **FLOATING
C249 w_dly_sig[5] VGND 1.76f $ **FLOATING
C250 w_dly_sig_n[4] VGND 0.782f $ **FLOATING
C251 w_dly_sig_n[3] VGND 0.938f $ **FLOATING
C252 a_12115_8573# VGND 0.609f $ **FLOATING
C253 a_12283_8475# VGND 0.97f $ **FLOATING
C254 a_11690_8573# VGND 0.626f $ **FLOATING
C255 a_11858_8319# VGND 0.581f $ **FLOATING
C256 a_11417_8207# VGND 1.43f $ **FLOATING
C257 a_11251_8207# VGND 1.81f $ **FLOATING
C258 a_9565_8207# VGND 0.23f $ **FLOATING
C259 a_9147_8207# VGND 0.581f $ **FLOATING
C260 a_9218_8181# VGND 0.626f $ **FLOATING
C261 a_9011_8181# VGND 1.81f $ **FLOATING
C262 a_9018_8481# VGND 1.43f $ **FLOATING
C263 a_8727_8181# VGND 0.609f $ **FLOATING
C264 a_8559_8181# VGND 0.97f $ **FLOATING
C265 a_21633_8751# VGND 0.23f $ **FLOATING
C266 a_18045_8751# VGND 0.23f $ **FLOATING
C267 a_16481_8751# VGND 0.23f $ **FLOATING
C268 a_14825_8751# VGND 0.23f $ **FLOATING
C269 a_13169_8751# VGND 0.23f $ **FLOATING
C270 _64_.X VGND 0.226f $ **FLOATING
C271 w_dly_sig_n[24] VGND 1.4f $ **FLOATING
C272 a_22143_8751# VGND 0.609f $ **FLOATING
C273 a_22311_8725# VGND 0.97f $ **FLOATING
C274 a_21718_8751# VGND 0.626f $ **FLOATING
C275 a_21886_8725# VGND 0.581f $ **FLOATING
C276 a_21445_8757# VGND 1.43f $ **FLOATING
C277 a_21279_8757# VGND 1.81f $ **FLOATING
C278 a_18555_8751# VGND 0.609f $ **FLOATING
C279 a_18723_8725# VGND 0.97f $ **FLOATING
C280 a_18130_8751# VGND 0.626f $ **FLOATING
C281 a_18298_8725# VGND 0.581f $ **FLOATING
C282 a_17857_8757# VGND 1.43f $ **FLOATING
C283 a_17691_8757# VGND 1.81f $ **FLOATING
C284 a_16991_8751# VGND 0.609f $ **FLOATING
C285 a_17159_8725# VGND 0.97f $ **FLOATING
C286 a_16566_8751# VGND 0.626f $ **FLOATING
C287 a_16734_8725# VGND 0.581f $ **FLOATING
C288 a_16293_8757# VGND 1.43f $ **FLOATING
C289 a_16127_8757# VGND 1.81f $ **FLOATING
C290 clknet_3_4__leaf_i_stop VGND 9.75f $ **FLOATING
C291 a_15335_8751# VGND 0.609f $ **FLOATING
C292 a_15503_8725# VGND 0.97f $ **FLOATING
C293 a_14910_8751# VGND 0.626f $ **FLOATING
C294 a_15078_8725# VGND 0.581f $ **FLOATING
C295 a_14637_8757# VGND 1.43f $ **FLOATING
C296 w_dly_sig[4] VGND 1.73f $ **FLOATING
C297 a_14471_8757# VGND 1.81f $ **FLOATING
C298 a_13679_8751# VGND 0.609f $ **FLOATING
C299 a_13847_8725# VGND 0.97f $ **FLOATING
C300 a_13254_8751# VGND 0.626f $ **FLOATING
C301 a_13422_8725# VGND 0.581f $ **FLOATING
C302 a_12981_8757# VGND 1.43f $ **FLOATING
C303 w_dly_sig[3] VGND 1.9f $ **FLOATING
C304 a_12815_8757# VGND 1.81f $ **FLOATING
C305 clknet_3_1__leaf_i_stop VGND 8.27f $ **FLOATING
C306 w_dly_sig_n[2] VGND 0.899f $ **FLOATING
C307 w_dly_sig[2] VGND 1.69f $ **FLOATING
C308 w_dly_sig_n[1] VGND 0.782f $ **FLOATING
C309 a_10975_8759# VGND 0.648f $ **FLOATING
C310 w_dly_sig_n[0] VGND 0.782f $ **FLOATING
C311 net1 VGND 5.34f $ **FLOATING
C312 w_dly_sig[24] VGND 2.1f $ **FLOATING
C313 w_dly_sig[25] VGND 2.03f $ **FLOATING
C314 w_dly_sig_n[25] VGND 0.782f $ **FLOATING
C315 a_855_8751# VGND 0.524f $ **FLOATING
C316 a_22553_9295# VGND 0.23f $ **FLOATING
C317 a_23063_9661# VGND 0.609f $ **FLOATING
C318 a_23231_9563# VGND 0.97f $ **FLOATING
C319 a_22638_9661# VGND 0.626f $ **FLOATING
C320 a_22806_9407# VGND 0.581f $ **FLOATING
C321 a_22365_9295# VGND 1.43f $ **FLOATING
C322 a_22199_9295# VGND 1.81f $ **FLOATING
C323 clknet_3_5__leaf_i_stop VGND 8.8f $ **FLOATING
C324 w_dly_sig_n[48] VGND 1.15f $ **FLOATING
C325 a_19701_9295# VGND 0.23f $ **FLOATING
C326 w_dly_sig[49] VGND 2f $ **FLOATING
C327 w_dly_sig[48] VGND 1.54f $ **FLOATING
C328 w_dly_sig_n[47] VGND 0.782f $ **FLOATING
C329 a_20211_9661# VGND 0.609f $ **FLOATING
C330 a_20379_9563# VGND 0.97f $ **FLOATING
C331 a_19786_9661# VGND 0.626f $ **FLOATING
C332 a_19954_9407# VGND 0.581f $ **FLOATING
C333 a_19513_9295# VGND 1.43f $ **FLOATING
C334 w_dly_sig[47] VGND 1.92f $ **FLOATING
C335 a_19347_9295# VGND 1.81f $ **FLOATING
C336 a_16481_9295# VGND 0.23f $ **FLOATING
C337 w_dly_sig[44] VGND 1.56f $ **FLOATING
C338 w_dly_sig_n[43] VGND 1.79f $ **FLOATING
C339 w_dly_sig_n[44] VGND 0.93f $ **FLOATING
C340 a_16991_9661# VGND 0.609f $ **FLOATING
C341 a_17159_9563# VGND 0.97f $ **FLOATING
C342 a_16566_9661# VGND 0.626f $ **FLOATING
C343 a_16734_9407# VGND 0.581f $ **FLOATING
C344 a_16293_9295# VGND 1.43f $ **FLOATING
C345 a_16127_9295# VGND 1.81f $ **FLOATING
C346 w_dly_sig[43] VGND 1.99f $ **FLOATING
C347 w_dly_sig_n[40] VGND 1.02f $ **FLOATING
C348 a_11865_9295# VGND 0.23f $ **FLOATING
C349 w_dly_sig[1] VGND 1.97f $ **FLOATING
C350 a_11447_9295# VGND 0.581f $ **FLOATING
C351 a_11518_9269# VGND 0.626f $ **FLOATING
C352 a_11311_9269# VGND 1.81f $ **FLOATING
C353 a_11318_9569# VGND 1.43f $ **FLOATING
C354 a_11027_9269# VGND 0.609f $ **FLOATING
C355 a_10859_9269# VGND 0.97f $ **FLOATING
C356 clknet_3_0__leaf_i_stop VGND 9.61f $ **FLOATING
C357 a_9473_9295# VGND 0.23f $ **FLOATING
C358 w_dly_sig[26] VGND 1.72f $ **FLOATING
C359 a_9055_9295# VGND 0.581f $ **FLOATING
C360 a_9126_9269# VGND 0.626f $ **FLOATING
C361 a_8919_9269# VGND 1.81f $ **FLOATING
C362 a_8926_9569# VGND 1.43f $ **FLOATING
C363 a_8635_9269# VGND 0.609f $ **FLOATING
C364 a_8467_9269# VGND 0.97f $ **FLOATING
C365 a_22369_9839# VGND 0.23f $ **FLOATING
C366 w_dly_sig_n[46] VGND 1.17f $ **FLOATING
C367 a_18413_9839# VGND 0.23f $ **FLOATING
C368 w_dly_sig_n[42] VGND 1.01f $ **FLOATING
C369 a_14089_9839# VGND 0.23f $ **FLOATING
C370 a_13262_10217# VGND 0.216f $ **FLOATING
C371 a_10209_10217# VGND 0.23f $ **FLOATING
C372 w_dly_sig_n[49] VGND 1.73f $ **FLOATING
C373 a_22879_9839# VGND 0.609f $ **FLOATING
C374 a_23047_9813# VGND 0.97f $ **FLOATING
C375 a_22454_9839# VGND 0.626f $ **FLOATING
C376 a_22622_9813# VGND 0.581f $ **FLOATING
C377 a_22181_9845# VGND 1.43f $ **FLOATING
C378 a_22015_9845# VGND 1.81f $ **FLOATING
C379 w_dly_sig_n[50] VGND 0.813f $ **FLOATING
C380 w_dly_sig[50] VGND 2.29f $ **FLOATING
C381 w_dly_sig_n[45] VGND 1.36f $ **FLOATING
C382 a_18923_9839# VGND 0.609f $ **FLOATING
C383 a_19091_9813# VGND 0.97f $ **FLOATING
C384 a_18498_9839# VGND 0.626f $ **FLOATING
C385 a_18666_9813# VGND 0.581f $ **FLOATING
C386 a_18225_9845# VGND 1.43f $ **FLOATING
C387 w_dly_sig[45] VGND 1.85f $ **FLOATING
C388 a_18059_9845# VGND 1.81f $ **FLOATING
C389 a_16197_9813# VGND 4.03f $ **FLOATING
C390 w_dly_sig[42] VGND 1.91f $ **FLOATING
C391 w_dly_sig_n[41] VGND 1.39f $ **FLOATING
C392 a_14599_9839# VGND 0.609f $ **FLOATING
C393 a_14767_9813# VGND 0.97f $ **FLOATING
C394 a_14174_9839# VGND 0.626f $ **FLOATING
C395 a_14342_9813# VGND 0.581f $ **FLOATING
C396 a_13901_9845# VGND 1.43f $ **FLOATING
C397 w_dly_sig[41] VGND 1.77f $ **FLOATING
C398 a_13735_9845# VGND 1.81f $ **FLOATING
C399 w_dly_sig[40] VGND 2.1f $ **FLOATING
C400 a_12821_10217# VGND 0.587f $ **FLOATING
C401 a_12892_10116# VGND 0.627f $ **FLOATING
C402 a_12698_9961# VGND 1.39f $ **FLOATING
C403 a_12688_10057# VGND 1.77f $ **FLOATING
C404 a_12400_9813# VGND 0.599f $ **FLOATING
C405 a_12050_9813# VGND 1.41f $ **FLOATING
C406 a_9791_10217# VGND 0.581f $ **FLOATING
C407 a_9862_10116# VGND 0.626f $ **FLOATING
C408 a_9662_9961# VGND 1.43f $ **FLOATING
C409 a_9655_10057# VGND 1.81f $ **FLOATING
C410 a_9371_10071# VGND 0.609f $ **FLOATING
C411 a_9203_10071# VGND 0.97f $ **FLOATING
C412 w_dly_sig[27] VGND 1.87f $ **FLOATING
C413 w_dly_sig_n[26] VGND 1.18f $ **FLOATING
C414 a_22001_10383# VGND 0.23f $ **FLOATING
C415 a_22511_10749# VGND 0.609f $ **FLOATING
C416 a_22679_10651# VGND 0.97f $ **FLOATING
C417 a_22086_10749# VGND 0.626f $ **FLOATING
C418 a_22254_10495# VGND 0.581f $ **FLOATING
C419 a_21813_10383# VGND 1.43f $ **FLOATING
C420 a_21647_10383# VGND 1.81f $ **FLOATING
C421 a_19885_10383# VGND 0.216f $ **FLOATING
C422 w_dly_sig[51] VGND 1.51f $ **FLOATING
C423 a_20395_10749# VGND 0.599f $ **FLOATING
C424 a_20566_10636# VGND 1.41f $ **FLOATING
C425 a_19979_10749# VGND 0.627f $ **FLOATING
C426 a_20138_10519# VGND 0.587f $ **FLOATING
C427 a_19697_10383# VGND 1.39f $ **FLOATING
C428 w_dly_sig[46] VGND 1.52f $ **FLOATING
C429 a_19531_10383# VGND 1.77f $ **FLOATING
C430 a_16849_10383# VGND 0.23f $ **FLOATING
C431 a_17359_10749# VGND 0.609f $ **FLOATING
C432 a_17527_10651# VGND 0.97f $ **FLOATING
C433 a_16934_10749# VGND 0.626f $ **FLOATING
C434 a_17102_10495# VGND 0.581f $ **FLOATING
C435 a_16661_10383# VGND 1.43f $ **FLOATING
C436 a_16495_10383# VGND 1.81f $ **FLOATING
C437 w_dly_sig_n[39] VGND 0.991f $ **FLOATING
C438 a_10485_10383# VGND 0.23f $ **FLOATING
C439 a_10067_10383# VGND 0.581f $ **FLOATING
C440 a_10138_10357# VGND 0.626f $ **FLOATING
C441 a_9931_10357# VGND 1.81f $ **FLOATING
C442 a_9938_10657# VGND 1.43f $ **FLOATING
C443 a_9647_10357# VGND 0.609f $ **FLOATING
C444 a_9479_10357# VGND 0.97f $ **FLOATING
C445 w_dly_sig_n[27] VGND 1.02f $ **FLOATING
C446 w_dly_sig[28] VGND 1.83f $ **FLOATING
C447 a_21909_10927# VGND 0.23f $ **FLOATING
C448 a_19701_10927# VGND 0.23f $ **FLOATING
C449 a_17861_10927# VGND 0.23f $ **FLOATING
C450 a_14641_10927# VGND 0.23f $ **FLOATING
C451 a_13077_10927# VGND 0.23f $ **FLOATING
C452 a_11513_10927# VGND 0.23f $ **FLOATING
C453 a_9933_11305# VGND 0.23f $ **FLOATING
C454 w_dly_sig_n[51] VGND 1.67f $ **FLOATING
C455 a_22419_10927# VGND 0.609f $ **FLOATING
C456 a_22587_10901# VGND 0.97f $ **FLOATING
C457 a_21994_10927# VGND 0.626f $ **FLOATING
C458 a_22162_10901# VGND 0.581f $ **FLOATING
C459 a_21721_10933# VGND 1.43f $ **FLOATING
C460 a_21555_10933# VGND 1.81f $ **FLOATING
C461 w_dly_sig[52] VGND 1.96f $ **FLOATING
C462 w_dly_sig_n[52] VGND 0.821f $ **FLOATING
C463 a_20211_10927# VGND 0.609f $ **FLOATING
C464 a_20379_10901# VGND 0.97f $ **FLOATING
C465 a_19786_10927# VGND 0.626f $ **FLOATING
C466 a_19954_10901# VGND 0.581f $ **FLOATING
C467 a_19513_10933# VGND 1.43f $ **FLOATING
C468 w_dly_sig[53] VGND 2.26f $ **FLOATING
C469 a_19347_10933# VGND 1.81f $ **FLOATING
C470 w_dly_sig_n[53] VGND 0.965f $ **FLOATING
C471 a_18371_10927# VGND 0.609f $ **FLOATING
C472 a_18539_10901# VGND 0.97f $ **FLOATING
C473 a_17946_10927# VGND 0.626f $ **FLOATING
C474 a_18114_10901# VGND 0.581f $ **FLOATING
C475 a_17673_10933# VGND 1.43f $ **FLOATING
C476 a_17507_10933# VGND 1.81f $ **FLOATING
C477 w_dly_sig[54] VGND 2.14f $ **FLOATING
C478 w_dly_sig_n[54] VGND 0.782f $ **FLOATING
C479 w_dly_sig_n[55] VGND 0.813f $ **FLOATING
C480 w_dly_sig[55] VGND 1.82f $ **FLOATING
C481 a_15151_10927# VGND 0.609f $ **FLOATING
C482 a_15319_10901# VGND 0.97f $ **FLOATING
C483 a_14726_10927# VGND 0.626f $ **FLOATING
C484 a_14894_10901# VGND 0.581f $ **FLOATING
C485 a_14453_10933# VGND 1.43f $ **FLOATING
C486 w_dly_sig[56] VGND 2.6f $ **FLOATING
C487 a_14287_10933# VGND 1.81f $ **FLOATING
C488 a_13587_10927# VGND 0.609f $ **FLOATING
C489 a_13755_10901# VGND 0.97f $ **FLOATING
C490 a_13162_10927# VGND 0.626f $ **FLOATING
C491 a_13330_10901# VGND 0.581f $ **FLOATING
C492 a_12889_10933# VGND 1.43f $ **FLOATING
C493 w_dly_sig[38] VGND 1.68f $ **FLOATING
C494 a_12723_10933# VGND 1.81f $ **FLOATING
C495 a_12023_10927# VGND 0.609f $ **FLOATING
C496 a_12191_10901# VGND 0.97f $ **FLOATING
C497 a_11598_10927# VGND 0.626f $ **FLOATING
C498 a_11766_10901# VGND 0.581f $ **FLOATING
C499 a_11325_10933# VGND 1.43f $ **FLOATING
C500 a_11159_10933# VGND 1.81f $ **FLOATING
C501 a_9515_11305# VGND 0.581f $ **FLOATING
C502 a_9586_11204# VGND 0.626f $ **FLOATING
C503 a_9386_11049# VGND 1.43f $ **FLOATING
C504 a_9379_11145# VGND 1.81f $ **FLOATING
C505 a_9095_11159# VGND 0.609f $ **FLOATING
C506 a_8927_11159# VGND 0.97f $ **FLOATING
C507 w_dly_sig_n[28] VGND 1.05f $ **FLOATING
C508 a_20345_11471# VGND 0.23f $ **FLOATING
C509 a_21822_11471# VGND 4.03f $ **FLOATING
C510 a_20855_11837# VGND 0.609f $ **FLOATING
C511 a_21023_11739# VGND 0.97f $ **FLOATING
C512 a_20430_11837# VGND 0.626f $ **FLOATING
C513 a_20598_11583# VGND 0.581f $ **FLOATING
C514 a_20157_11471# VGND 1.43f $ **FLOATING
C515 a_19991_11471# VGND 1.81f $ **FLOATING
C516 w_dly_sig[39] VGND 2.94f $ **FLOATING
C517 w_dly_sig_n[37] VGND 1.18f $ **FLOATING
C518 a_11513_11471# VGND 0.23f $ **FLOATING
C519 w_dly_sig_n[60] VGND 0.938f $ **FLOATING
C520 a_16749_11445# VGND 4.03f $ **FLOATING
C521 a_14449_11445# VGND 4.03f $ **FLOATING
C522 w_dly_sig_n[38] VGND 1.85f $ **FLOATING
C523 a_12023_11837# VGND 0.609f $ **FLOATING
C524 a_12191_11739# VGND 0.97f $ **FLOATING
C525 a_11598_11837# VGND 0.626f $ **FLOATING
C526 a_11766_11583# VGND 0.581f $ **FLOATING
C527 a_11325_11471# VGND 1.43f $ **FLOATING
C528 a_11159_11471# VGND 1.81f $ **FLOATING
C529 clknet_0_i_stop VGND 19.1f $ **FLOATING
C530 a_9389_11445# VGND 4.03f $ **FLOATING
C531 w_dly_sig_n[29] VGND 0.782f $ **FLOATING
C532 w_dly_sig[29] VGND 2.04f $ **FLOATING
C533 a_22553_12015# VGND 0.23f $ **FLOATING
C534 a_19609_12015# VGND 0.23f $ **FLOATING
C535 a_18045_12015# VGND 0.23f $ **FLOATING
C536 a_16481_12015# VGND 0.23f $ **FLOATING
C537 w_dly_sig_n[57] VGND 1.21f $ **FLOATING
C538 a_14181_12015# VGND 0.23f $ **FLOATING
C539 a_12617_12015# VGND 0.23f $ **FLOATING
C540 a_9841_12393# VGND 0.23f $ **FLOATING
C541 a_23063_12015# VGND 0.609f $ **FLOATING
C542 a_23231_11989# VGND 0.97f $ **FLOATING
C543 a_22638_12015# VGND 0.626f $ **FLOATING
C544 a_22806_11989# VGND 0.581f $ **FLOATING
C545 a_22365_12021# VGND 1.43f $ **FLOATING
C546 a_22199_12021# VGND 1.81f $ **FLOATING
C547 a_20119_12015# VGND 0.609f $ **FLOATING
C548 a_20287_11989# VGND 0.97f $ **FLOATING
C549 a_19694_12015# VGND 0.626f $ **FLOATING
C550 a_19862_11989# VGND 0.581f $ **FLOATING
C551 a_19421_12021# VGND 1.43f $ **FLOATING
C552 w_dly_sig[60] VGND 1.81f $ **FLOATING
C553 a_19255_12021# VGND 1.81f $ **FLOATING
C554 a_18555_12015# VGND 0.609f $ **FLOATING
C555 a_18723_11989# VGND 0.97f $ **FLOATING
C556 a_18130_12015# VGND 0.626f $ **FLOATING
C557 a_18298_11989# VGND 0.581f $ **FLOATING
C558 a_17857_12021# VGND 1.43f $ **FLOATING
C559 a_17691_12021# VGND 1.81f $ **FLOATING
C560 a_16991_12015# VGND 0.609f $ **FLOATING
C561 a_17159_11989# VGND 0.97f $ **FLOATING
C562 a_16566_12015# VGND 0.626f $ **FLOATING
C563 a_16734_11989# VGND 0.581f $ **FLOATING
C564 a_16293_12021# VGND 1.43f $ **FLOATING
C565 a_16127_12021# VGND 1.81f $ **FLOATING
C566 w_dly_sig[57] VGND 1.54f $ **FLOATING
C567 w_dly_sig_n[56] VGND 1.39f $ **FLOATING
C568 a_14691_12015# VGND 0.609f $ **FLOATING
C569 a_14859_11989# VGND 0.97f $ **FLOATING
C570 a_14266_12015# VGND 0.626f $ **FLOATING
C571 a_14434_11989# VGND 0.581f $ **FLOATING
C572 a_13993_12021# VGND 1.43f $ **FLOATING
C573 w_dly_sig[36] VGND 1.83f $ **FLOATING
C574 a_13827_12021# VGND 1.81f $ **FLOATING
C575 a_13127_12015# VGND 0.609f $ **FLOATING
C576 a_13295_11989# VGND 0.97f $ **FLOATING
C577 a_12702_12015# VGND 0.626f $ **FLOATING
C578 a_12870_11989# VGND 0.581f $ **FLOATING
C579 a_12429_12021# VGND 1.43f $ **FLOATING
C580 a_12263_12021# VGND 1.81f $ **FLOATING
C581 a_9423_12393# VGND 0.581f $ **FLOATING
C582 a_9494_12292# VGND 0.626f $ **FLOATING
C583 a_9294_12137# VGND 1.43f $ **FLOATING
C584 a_9287_12233# VGND 1.81f $ **FLOATING
C585 a_9003_12247# VGND 0.609f $ **FLOATING
C586 a_8835_12247# VGND 0.97f $ **FLOATING
C587 g_dly_chain_even[64].dly_stg2.Y VGND 0.238f $ **FLOATING
C588 w_dly_sig[64] VGND 1.52f $ **FLOATING
C589 w_dly_sig_n[59] VGND 1.41f $ **FLOATING
C590 a_16297_12559# VGND 0.23f $ **FLOATING
C591 w_dly_sig_n[64] VGND 1.13f $ **FLOATING
C592 w_dly_sig_n[63] VGND 0.93f $ **FLOATING
C593 w_dly_sig_n[61] VGND 0.782f $ **FLOATING
C594 w_dly_sig[61] VGND 2.04f $ **FLOATING
C595 w_dly_sig[59] VGND 1.52f $ **FLOATING
C596 w_dly_sig_n[58] VGND 0.782f $ **FLOATING
C597 a_16807_12925# VGND 0.609f $ **FLOATING
C598 a_16975_12827# VGND 0.97f $ **FLOATING
C599 a_16382_12925# VGND 0.626f $ **FLOATING
C600 a_16550_12671# VGND 0.581f $ **FLOATING
C601 a_16109_12559# VGND 1.43f $ **FLOATING
C602 w_dly_sig[58] VGND 2.14f $ **FLOATING
C603 a_15943_12559# VGND 1.81f $ **FLOATING
C604 clknet_3_6__leaf_i_stop VGND 10.2f $ **FLOATING
C605 a_14365_12559# VGND 0.23f $ **FLOATING
C606 a_14875_12925# VGND 0.609f $ **FLOATING
C607 a_15043_12827# VGND 0.97f $ **FLOATING
C608 a_14450_12925# VGND 0.626f $ **FLOATING
C609 a_14618_12671# VGND 0.581f $ **FLOATING
C610 a_14177_12559# VGND 1.43f $ **FLOATING
C611 a_14011_12559# VGND 1.81f $ **FLOATING
C612 w_dly_sig_n[35] VGND 1.21f $ **FLOATING
C613 w_dly_sig[37] VGND 1.82f $ **FLOATING
C614 a_10961_12559# VGND 0.23f $ **FLOATING
C615 w_dly_sig[35] VGND 1.62f $ **FLOATING
C616 w_dly_sig_n[34] VGND 0.93f $ **FLOATING
C617 w_dly_sig_n[36] VGND 1.23f $ **FLOATING
C618 w_dly_sig_n[33] VGND 1.33f $ **FLOATING
C619 a_11471_12925# VGND 0.609f $ **FLOATING
C620 a_11639_12827# VGND 0.97f $ **FLOATING
C621 a_11046_12925# VGND 0.626f $ **FLOATING
C622 a_11214_12671# VGND 0.581f $ **FLOATING
C623 a_10773_12559# VGND 1.43f $ **FLOATING
C624 a_10607_12559# VGND 1.81f $ **FLOATING
C625 w_dly_sig[33] VGND 1.72f $ **FLOATING
C626 w_dly_sig_n[30] VGND 1.3f $ **FLOATING
C627 w_dly_sig_n[32] VGND 0.998f $ **FLOATING
C628 w_dly_sig_n[31] VGND 1.32f $ **FLOATING
C629 w_dly_sig[30] VGND 2.63f $ **FLOATING
C630 w_dly_sig[31] VGND 1.98f $ **FLOATING
C631 a_22185_13103# VGND 0.23f $ **FLOATING
C632 a_19977_13103# VGND 0.23f $ **FLOATING
C633 a_12525_13103# VGND 0.23f $ **FLOATING
C634 a_10117_13481# VGND 0.23f $ **FLOATING
C635 a_22695_13103# VGND 0.609f $ **FLOATING
C636 a_22863_13077# VGND 0.97f $ **FLOATING
C637 a_22270_13103# VGND 0.626f $ **FLOATING
C638 a_22438_13077# VGND 0.581f $ **FLOATING
C639 a_21997_13109# VGND 1.43f $ **FLOATING
C640 w_dly_sig[63] VGND 1.95f $ **FLOATING
C641 a_21831_13109# VGND 1.81f $ **FLOATING
C642 w_dly_sig_n[62] VGND 0.782f $ **FLOATING
C643 a_20487_13103# VGND 0.609f $ **FLOATING
C644 a_20655_13077# VGND 0.97f $ **FLOATING
C645 a_20062_13103# VGND 0.626f $ **FLOATING
C646 a_20230_13077# VGND 0.581f $ **FLOATING
C647 a_19789_13109# VGND 1.43f $ **FLOATING
C648 w_dly_sig[62] VGND 2.34f $ **FLOATING
C649 a_19623_13109# VGND 1.81f $ **FLOATING
C650 clknet_3_7__leaf_i_stop VGND 13.4f $ **FLOATING
C651 a_13035_13103# VGND 0.609f $ **FLOATING
C652 a_13203_13077# VGND 0.97f $ **FLOATING
C653 a_12610_13103# VGND 0.626f $ **FLOATING
C654 a_12778_13077# VGND 0.581f $ **FLOATING
C655 a_12337_13109# VGND 1.43f $ **FLOATING
C656 w_dly_sig[34] VGND 1.6f $ **FLOATING
C657 a_12171_13109# VGND 1.81f $ **FLOATING
C658 clknet_3_3__leaf_i_stop VGND 10.3f $ **FLOATING
C659 clknet_3_2__leaf_i_stop VGND 8.17f $ **FLOATING
C660 w_dly_sig[32] VGND 1.79f $ **FLOATING
C661 a_9699_13481# VGND 0.581f $ **FLOATING
C662 a_9770_13380# VGND 0.626f $ **FLOATING
C663 a_9570_13225# VGND 1.43f $ **FLOATING
C664 a_9563_13321# VGND 1.81f $ **FLOATING
C665 a_9279_13335# VGND 0.609f $ **FLOATING
C666 a_9111_13335# VGND 0.97f $ **FLOATING
.ends
