magic
tech sky130A
magscale 1 2
timestamp 1710678572
<< viali >>
rect 10701 18853 10735 18887
rect 1409 18785 1443 18819
rect 6561 18785 6595 18819
rect 7205 18785 7239 18819
rect 7849 18785 7883 18819
rect 8585 18785 8619 18819
rect 9689 18785 9723 18819
rect 9873 18785 9907 18819
rect 9965 18785 9999 18819
rect 10241 18785 10275 18819
rect 10517 18785 10551 18819
rect 10609 18785 10643 18819
rect 11161 18785 11195 18819
rect 11417 18785 11451 18819
rect 13912 18785 13946 18819
rect 16129 18785 16163 18819
rect 16396 18785 16430 18819
rect 19248 18785 19282 18819
rect 20821 18785 20855 18819
rect 20913 18785 20947 18819
rect 21281 18785 21315 18819
rect 22017 18785 22051 18819
rect 22293 18785 22327 18819
rect 22845 18785 22879 18819
rect 24970 18785 25004 18819
rect 27813 18785 27847 18819
rect 28457 18785 28491 18819
rect 30757 18785 30791 18819
rect 1133 18717 1167 18751
rect 9597 18717 9631 18751
rect 13645 18717 13679 18751
rect 18981 18717 19015 18751
rect 25237 18717 25271 18751
rect 21373 18649 21407 18683
rect 21925 18649 21959 18683
rect 22201 18649 22235 18683
rect 857 18581 891 18615
rect 8493 18581 8527 18615
rect 10149 18581 10183 18615
rect 10425 18581 10459 18615
rect 12541 18581 12575 18615
rect 15025 18581 15059 18615
rect 17509 18581 17543 18615
rect 20361 18581 20395 18615
rect 22753 18581 22787 18615
rect 23857 18581 23891 18615
rect 31033 18581 31067 18615
rect 9505 18377 9539 18411
rect 12909 18377 12943 18411
rect 14197 18377 14231 18411
rect 21005 18377 21039 18411
rect 22753 18377 22787 18411
rect 23029 18377 23063 18411
rect 8493 18309 8527 18343
rect 11621 18309 11655 18343
rect 13921 18309 13955 18343
rect 7021 18241 7055 18275
rect 7573 18241 7607 18275
rect 7849 18241 7883 18275
rect 9965 18241 9999 18275
rect 14565 18241 14599 18275
rect 17141 18241 17175 18275
rect 857 18173 891 18207
rect 7113 18173 7147 18207
rect 7481 18173 7515 18207
rect 7941 18173 7975 18207
rect 8217 18173 8251 18207
rect 8585 18173 8619 18207
rect 8861 18173 8895 18207
rect 8953 18173 8987 18207
rect 9321 18173 9355 18207
rect 9597 18173 9631 18207
rect 9873 18173 9907 18207
rect 11713 18173 11747 18207
rect 11897 18173 11931 18207
rect 11989 18173 12023 18207
rect 12265 18173 12299 18207
rect 12357 18173 12391 18207
rect 13001 18173 13035 18207
rect 13737 18173 13771 18207
rect 13829 18173 13863 18207
rect 14105 18173 14139 18207
rect 14821 18173 14855 18207
rect 16773 18173 16807 18207
rect 17049 18173 17083 18207
rect 19349 18173 19383 18207
rect 19625 18173 19659 18207
rect 19901 18173 19935 18207
rect 20177 18173 20211 18207
rect 20729 18173 20763 18207
rect 21097 18173 21131 18207
rect 22385 18173 22419 18207
rect 22845 18173 22879 18207
rect 23121 18173 23155 18207
rect 23397 18173 23431 18207
rect 23489 18173 23523 18207
rect 24041 18173 24075 18207
rect 24409 18173 24443 18207
rect 24961 18173 24995 18207
rect 9781 18105 9815 18139
rect 10210 18105 10244 18139
rect 12173 18105 12207 18139
rect 17408 18105 17442 18139
rect 19809 18105 19843 18139
rect 20085 18105 20119 18139
rect 22293 18105 22327 18139
rect 23305 18105 23339 18139
rect 24869 18105 24903 18139
rect 8125 18037 8159 18071
rect 9229 18037 9263 18071
rect 11345 18037 11379 18071
rect 12449 18037 12483 18071
rect 13645 18037 13679 18071
rect 15945 18037 15979 18071
rect 16681 18037 16715 18071
rect 16957 18037 16991 18071
rect 18521 18037 18555 18071
rect 19257 18037 19291 18071
rect 19533 18037 19567 18071
rect 20637 18037 20671 18071
rect 23581 18037 23615 18071
rect 23949 18037 23983 18071
rect 24317 18037 24351 18071
rect 6745 17833 6779 17867
rect 7389 17833 7423 17867
rect 12265 17833 12299 17867
rect 12817 17833 12851 17867
rect 13093 17833 13127 17867
rect 13369 17833 13403 17867
rect 16221 17833 16255 17867
rect 24317 17833 24351 17867
rect 24593 17833 24627 17867
rect 25513 17833 25547 17867
rect 7665 17765 7699 17799
rect 8554 17765 8588 17799
rect 13890 17765 13924 17799
rect 22394 17765 22428 17799
rect 23866 17765 23900 17799
rect 25237 17765 25271 17799
rect 25789 17765 25823 17799
rect 6561 17697 6595 17731
rect 6837 17697 6871 17731
rect 7113 17697 7147 17731
rect 7481 17697 7515 17731
rect 7757 17697 7791 17731
rect 7849 17697 7883 17731
rect 12357 17697 12391 17731
rect 12633 17697 12667 17731
rect 12909 17697 12943 17731
rect 13185 17697 13219 17731
rect 13277 17697 13311 17731
rect 13645 17697 13679 17731
rect 16313 17697 16347 17731
rect 16661 17697 16695 17731
rect 17877 17697 17911 17731
rect 18613 17697 18647 17731
rect 19073 17697 19107 17731
rect 19349 17697 19383 17731
rect 19441 17697 19475 17731
rect 19717 17697 19751 17731
rect 22661 17697 22695 17731
rect 24409 17697 24443 17731
rect 24685 17697 24719 17731
rect 25329 17697 25363 17731
rect 25605 17697 25639 17731
rect 25881 17697 25915 17731
rect 26065 17697 26099 17731
rect 26157 17697 26191 17731
rect 8309 17629 8343 17663
rect 12541 17629 12575 17663
rect 16405 17629 16439 17663
rect 18705 17629 18739 17663
rect 18981 17629 19015 17663
rect 24133 17629 24167 17663
rect 17969 17561 18003 17595
rect 6469 17493 6503 17527
rect 7021 17493 7055 17527
rect 7941 17493 7975 17527
rect 9689 17493 9723 17527
rect 15025 17493 15059 17527
rect 17785 17493 17819 17527
rect 19257 17493 19291 17527
rect 19533 17493 19567 17527
rect 19809 17493 19843 17527
rect 21281 17493 21315 17527
rect 22753 17493 22787 17527
rect 6745 17289 6779 17323
rect 7297 17289 7331 17323
rect 11805 17289 11839 17323
rect 12081 17289 12115 17323
rect 19441 17289 19475 17323
rect 25053 17289 25087 17323
rect 25329 17289 25363 17323
rect 5089 17221 5123 17255
rect 16129 17221 16163 17255
rect 19717 17221 19751 17255
rect 20269 17221 20303 17255
rect 12633 17153 12667 17187
rect 14749 17153 14783 17187
rect 17877 17153 17911 17187
rect 21741 17153 21775 17187
rect 857 17085 891 17119
rect 3709 17085 3743 17119
rect 5549 17085 5583 17119
rect 5825 17085 5859 17119
rect 6101 17085 6135 17119
rect 6377 17085 6411 17119
rect 6837 17085 6871 17119
rect 7113 17085 7147 17119
rect 7389 17085 7423 17119
rect 9689 17085 9723 17119
rect 11897 17085 11931 17119
rect 12173 17085 12207 17119
rect 12265 17085 12299 17119
rect 12541 17085 12575 17119
rect 12817 17085 12851 17119
rect 15005 17085 15039 17119
rect 17621 17085 17655 17119
rect 19349 17085 19383 17119
rect 19625 17085 19659 17119
rect 20085 17085 20119 17119
rect 20177 17085 20211 17119
rect 20453 17085 20487 17119
rect 20729 17085 20763 17119
rect 21189 17085 21223 17119
rect 21465 17085 21499 17119
rect 25145 17085 25179 17119
rect 25421 17085 25455 17119
rect 25697 17085 25731 17119
rect 25789 17085 25823 17119
rect 26065 17085 26099 17119
rect 27721 17085 27755 17119
rect 3976 17017 4010 17051
rect 6009 17017 6043 17051
rect 6285 17017 6319 17051
rect 9934 17017 9968 17051
rect 20545 17017 20579 17051
rect 20821 17017 20855 17051
rect 21986 17017 22020 17051
rect 26157 17017 26191 17051
rect 27454 17017 27488 17051
rect 5457 16949 5491 16983
rect 5733 16949 5767 16983
rect 7021 16949 7055 16983
rect 11069 16949 11103 16983
rect 12357 16949 12391 16983
rect 12909 16949 12943 16983
rect 16497 16949 16531 16983
rect 19993 16949 20027 16983
rect 21097 16949 21131 16983
rect 21557 16949 21591 16983
rect 23121 16949 23155 16983
rect 25605 16949 25639 16983
rect 25881 16949 25915 16983
rect 26341 16949 26375 16983
rect 5273 16745 5307 16779
rect 11805 16745 11839 16779
rect 12173 16745 12207 16779
rect 12449 16745 12483 16779
rect 20085 16745 20119 16779
rect 25697 16745 25731 16779
rect 25973 16745 26007 16779
rect 27169 16745 27203 16779
rect 5549 16677 5583 16711
rect 13430 16677 13464 16711
rect 18052 16677 18086 16711
rect 27997 16677 28031 16711
rect 2053 16609 2087 16643
rect 3249 16609 3283 16643
rect 3709 16609 3743 16643
rect 3801 16609 3835 16643
rect 3893 16609 3927 16643
rect 4261 16609 4295 16643
rect 4537 16609 4571 16643
rect 4813 16609 4847 16643
rect 4905 16609 4939 16643
rect 5365 16609 5399 16643
rect 5641 16609 5675 16643
rect 6009 16609 6043 16643
rect 6193 16609 6227 16643
rect 6285 16609 6319 16643
rect 6377 16609 6411 16643
rect 6633 16609 6667 16643
rect 8033 16609 8067 16643
rect 8289 16609 8323 16643
rect 10149 16609 10183 16643
rect 11253 16609 11287 16643
rect 11529 16609 11563 16643
rect 11713 16609 11747 16643
rect 12081 16609 12115 16643
rect 12357 16609 12391 16643
rect 17785 16609 17819 16643
rect 19901 16609 19935 16643
rect 20177 16609 20211 16643
rect 20453 16599 20487 16633
rect 20729 16609 20763 16643
rect 21281 16609 21315 16643
rect 21741 16609 21775 16643
rect 22017 16609 22051 16643
rect 22201 16609 22235 16643
rect 22293 16609 22327 16643
rect 23581 16609 23615 16643
rect 23848 16609 23882 16643
rect 25789 16609 25823 16643
rect 26065 16609 26099 16643
rect 26801 16609 26835 16643
rect 27261 16609 27295 16643
rect 27353 16609 27387 16643
rect 27445 16609 27479 16643
rect 27813 16609 27847 16643
rect 28089 16609 28123 16643
rect 29754 16609 29788 16643
rect 13185 16541 13219 16575
rect 27721 16541 27755 16575
rect 30021 16541 30055 16575
rect 19809 16473 19843 16507
rect 20361 16473 20395 16507
rect 21373 16473 21407 16507
rect 1961 16405 1995 16439
rect 3341 16405 3375 16439
rect 3617 16405 3651 16439
rect 4169 16405 4203 16439
rect 4445 16405 4479 16439
rect 5917 16405 5951 16439
rect 7757 16405 7791 16439
rect 9413 16405 9447 16439
rect 10241 16405 10275 16439
rect 11161 16405 11195 16439
rect 11437 16405 11471 16439
rect 14565 16405 14599 16439
rect 19165 16405 19199 16439
rect 20821 16405 20855 16439
rect 21649 16405 21683 16439
rect 21925 16405 21959 16439
rect 24961 16405 24995 16439
rect 26893 16405 26927 16439
rect 28641 16405 28675 16439
rect 1869 16201 1903 16235
rect 11069 16201 11103 16235
rect 11437 16201 11471 16235
rect 19349 16201 19383 16235
rect 19625 16201 19659 16235
rect 26893 16201 26927 16235
rect 27629 16201 27663 16235
rect 28733 16201 28767 16235
rect 29101 16201 29135 16235
rect 2421 16133 2455 16167
rect 9781 16133 9815 16167
rect 20085 16133 20119 16167
rect 20361 16133 20395 16167
rect 23489 16133 23523 16167
rect 8401 16065 8435 16099
rect 17509 16065 17543 16099
rect 26709 16065 26743 16099
rect 29377 16065 29411 16099
rect 1685 15997 1719 16031
rect 1961 15997 1995 16031
rect 2053 15997 2087 16031
rect 2145 15997 2179 16031
rect 2513 15997 2547 16031
rect 2789 15997 2823 16031
rect 2973 15997 3007 16031
rect 3065 15997 3099 16031
rect 3525 15997 3559 16031
rect 3617 15997 3651 16031
rect 4997 15997 5031 16031
rect 8657 15997 8691 16031
rect 9873 15997 9907 16031
rect 10333 15997 10367 16031
rect 10609 15997 10643 16031
rect 10885 15997 10919 16031
rect 10977 15997 11011 16031
rect 11529 15997 11563 16031
rect 11989 15997 12023 16031
rect 14657 15997 14691 16031
rect 17253 15997 17287 16031
rect 18889 15997 18923 16031
rect 19165 15997 19199 16031
rect 19449 15997 19483 16031
rect 19725 15997 19759 16031
rect 19993 15997 20027 16031
rect 20453 15997 20487 16031
rect 20729 15997 20763 16031
rect 20821 15997 20855 16031
rect 21281 15997 21315 16031
rect 21557 15997 21591 16031
rect 22109 15997 22143 16031
rect 22376 15997 22410 16031
rect 25237 15997 25271 16031
rect 26985 15997 27019 16031
rect 27537 15997 27571 16031
rect 27997 15997 28031 16031
rect 28273 15997 28307 16031
rect 28549 15997 28583 16031
rect 28825 15997 28859 16031
rect 29193 15997 29227 16031
rect 29469 15997 29503 16031
rect 1593 15929 1627 15963
rect 3433 15929 3467 15963
rect 5242 15929 5276 15963
rect 10517 15929 10551 15963
rect 10793 15929 10827 15963
rect 12234 15929 12268 15963
rect 14924 15929 14958 15963
rect 24992 15929 25026 15963
rect 26442 15929 26476 15963
rect 28181 15929 28215 15963
rect 2697 15861 2731 15895
rect 3709 15861 3743 15895
rect 6377 15861 6411 15895
rect 9965 15861 9999 15895
rect 10241 15861 10275 15895
rect 13369 15861 13403 15895
rect 16037 15861 16071 15895
rect 16129 15861 16163 15895
rect 18797 15861 18831 15895
rect 19073 15861 19107 15895
rect 20637 15861 20671 15895
rect 20913 15861 20947 15895
rect 21189 15861 21223 15895
rect 21465 15861 21499 15895
rect 23857 15861 23891 15895
rect 25329 15861 25363 15895
rect 27905 15861 27939 15895
rect 28457 15861 28491 15895
rect 9229 15657 9263 15691
rect 10057 15657 10091 15691
rect 10609 15657 10643 15691
rect 19073 15657 19107 15691
rect 28181 15657 28215 15691
rect 28457 15657 28491 15691
rect 2942 15589 2976 15623
rect 6714 15589 6748 15623
rect 18521 15589 18555 15623
rect 19616 15589 19650 15623
rect 22170 15589 22204 15623
rect 27546 15589 27580 15623
rect 1317 15521 1351 15555
rect 1593 15521 1627 15555
rect 1869 15521 1903 15555
rect 1961 15521 1995 15555
rect 2237 15521 2271 15555
rect 4169 15521 4203 15555
rect 4425 15521 4459 15555
rect 6469 15521 6503 15555
rect 9321 15521 9355 15555
rect 9597 15521 9631 15555
rect 9689 15521 9723 15555
rect 10149 15521 10183 15555
rect 10425 15521 10459 15555
rect 10517 15521 10551 15555
rect 11529 15521 11563 15555
rect 11785 15521 11819 15555
rect 13645 15521 13679 15555
rect 13901 15521 13935 15555
rect 15301 15521 15335 15555
rect 15577 15521 15611 15555
rect 16865 15521 16899 15555
rect 17141 15521 17175 15555
rect 17417 15521 17451 15555
rect 17693 15521 17727 15555
rect 18337 15521 18371 15555
rect 18613 15521 18647 15555
rect 18889 15521 18923 15555
rect 19165 15521 19199 15555
rect 21005 15521 21039 15555
rect 21925 15521 21959 15555
rect 24312 15521 24346 15555
rect 24409 15521 24443 15555
rect 24501 15521 24535 15555
rect 24629 15521 24663 15555
rect 24777 15521 24811 15555
rect 28273 15521 28307 15555
rect 28549 15521 28583 15555
rect 28825 15511 28859 15545
rect 29101 15521 29135 15555
rect 29201 15519 29235 15553
rect 29561 15521 29595 15555
rect 29817 15521 29851 15555
rect 2697 15453 2731 15487
rect 10333 15453 10367 15487
rect 17325 15453 17359 15487
rect 17601 15453 17635 15487
rect 18245 15453 18279 15487
rect 19349 15453 19383 15487
rect 27813 15453 27847 15487
rect 28733 15453 28767 15487
rect 9781 15385 9815 15419
rect 29285 15385 29319 15419
rect 1225 15317 1259 15351
rect 1501 15317 1535 15351
rect 1777 15317 1811 15351
rect 2053 15317 2087 15351
rect 2329 15317 2363 15351
rect 4077 15317 4111 15351
rect 5549 15317 5583 15351
rect 7849 15317 7883 15351
rect 9505 15317 9539 15351
rect 12909 15317 12943 15351
rect 15025 15317 15059 15351
rect 15209 15317 15243 15351
rect 15485 15317 15519 15351
rect 16773 15317 16807 15351
rect 17049 15317 17083 15351
rect 18797 15317 18831 15351
rect 20729 15317 20763 15351
rect 20913 15317 20947 15351
rect 23305 15317 23339 15351
rect 24133 15317 24167 15351
rect 26433 15317 26467 15351
rect 29009 15317 29043 15351
rect 30941 15317 30975 15351
rect 1961 15113 1995 15147
rect 9321 15113 9355 15147
rect 14749 15113 14783 15147
rect 15577 15113 15611 15147
rect 19257 15113 19291 15147
rect 25237 15113 25271 15147
rect 28733 15113 28767 15147
rect 29929 15113 29963 15147
rect 8217 15045 8251 15079
rect 11437 15045 11471 15079
rect 15301 15045 15335 15079
rect 24501 15045 24535 15079
rect 28457 15045 28491 15079
rect 29101 15045 29135 15079
rect 6837 14977 6871 15011
rect 15025 14977 15059 15011
rect 16221 14977 16255 15011
rect 20729 14977 20763 15011
rect 1777 14909 1811 14943
rect 2053 14909 2087 14943
rect 2145 14909 2179 14943
rect 4629 14909 4663 14943
rect 9413 14909 9447 14943
rect 9689 14909 9723 14943
rect 9781 14909 9815 14943
rect 10057 14909 10091 14943
rect 11989 14909 12023 14943
rect 12256 14909 12290 14943
rect 14289 14909 14323 14943
rect 14565 14909 14599 14943
rect 14841 14909 14875 14943
rect 15117 14909 15151 14943
rect 15393 14909 15427 14943
rect 15669 14909 15703 14943
rect 15761 14909 15795 14943
rect 15853 14909 15887 14943
rect 16488 14909 16522 14943
rect 17693 14909 17727 14943
rect 17877 14909 17911 14943
rect 18061 14909 18095 14943
rect 18705 14909 18739 14943
rect 18889 14909 18923 14943
rect 18981 14909 19015 14943
rect 19073 14909 19107 14943
rect 20996 14909 21030 14943
rect 23857 14909 23891 14943
rect 23950 14909 23984 14943
rect 24133 14909 24167 14943
rect 24363 14909 24397 14943
rect 26617 14909 26651 14943
rect 28549 14909 28583 14943
rect 28825 14909 28859 14943
rect 29193 14909 29227 14943
rect 29469 14909 29503 14943
rect 29561 14909 29595 14943
rect 29837 14909 29871 14943
rect 4874 14841 4908 14875
rect 7082 14841 7116 14875
rect 9873 14841 9907 14875
rect 10324 14841 10358 14875
rect 17969 14841 18003 14875
rect 24225 14841 24259 14875
rect 26372 14841 26406 14875
rect 1685 14773 1719 14807
rect 2237 14773 2271 14807
rect 6009 14773 6043 14807
rect 9597 14773 9631 14807
rect 13369 14773 13403 14807
rect 14197 14773 14231 14807
rect 14473 14773 14507 14807
rect 17601 14773 17635 14807
rect 18245 14773 18279 14807
rect 22109 14773 22143 14807
rect 29377 14773 29411 14807
rect 29653 14773 29687 14807
rect 4169 14569 4203 14603
rect 7941 14569 7975 14603
rect 9413 14569 9447 14603
rect 10517 14569 10551 14603
rect 15393 14569 15427 14603
rect 20913 14569 20947 14603
rect 26801 14569 26835 14603
rect 27445 14569 27479 14603
rect 28825 14569 28859 14603
rect 29377 14569 29411 14603
rect 30941 14569 30975 14603
rect 3034 14501 3068 14535
rect 13737 14501 13771 14535
rect 13953 14501 13987 14535
rect 21465 14501 21499 14535
rect 22201 14501 22235 14535
rect 22339 14501 22373 14535
rect 23213 14501 23247 14535
rect 23673 14501 23707 14535
rect 24837 14501 24871 14535
rect 25053 14501 25087 14535
rect 27721 14501 27755 14535
rect 28273 14501 28307 14535
rect 29806 14501 29840 14535
rect 22523 14467 22557 14501
rect 22983 14467 23017 14501
rect 23443 14467 23477 14501
rect 1409 14433 1443 14467
rect 1685 14433 1719 14467
rect 1961 14433 1995 14467
rect 2237 14433 2271 14467
rect 2513 14433 2547 14467
rect 4629 14433 4663 14467
rect 5089 14433 5123 14467
rect 5825 14433 5859 14467
rect 5917 14433 5951 14467
rect 6193 14433 6227 14467
rect 6561 14433 6595 14467
rect 6817 14433 6851 14467
rect 9505 14433 9539 14467
rect 9597 14433 9631 14467
rect 10057 14433 10091 14467
rect 10333 14433 10367 14467
rect 10425 14433 10459 14467
rect 10977 14433 11011 14467
rect 11244 14433 11278 14467
rect 12633 14433 12667 14467
rect 13093 14433 13127 14467
rect 13185 14433 13219 14467
rect 13621 14433 13655 14467
rect 14197 14433 14231 14467
rect 14749 14433 14783 14467
rect 15117 14433 15151 14467
rect 15209 14433 15243 14467
rect 15301 14433 15335 14467
rect 16589 14433 16623 14467
rect 16845 14433 16879 14467
rect 19540 14433 19574 14467
rect 19789 14433 19823 14467
rect 23949 14433 23983 14467
rect 24042 14433 24076 14467
rect 24225 14433 24259 14467
rect 24317 14433 24351 14467
rect 24455 14433 24489 14467
rect 26433 14433 26467 14467
rect 26525 14433 26559 14467
rect 26893 14433 26927 14467
rect 27537 14433 27571 14467
rect 27629 14433 27663 14467
rect 27905 14433 27939 14467
rect 28365 14433 28399 14467
rect 28641 14433 28675 14467
rect 28733 14433 28767 14467
rect 29009 14433 29043 14467
rect 29469 14433 29503 14467
rect 1593 14365 1627 14399
rect 2789 14365 2823 14399
rect 13001 14365 13035 14399
rect 13277 14365 13311 14399
rect 29561 14365 29595 14399
rect 1317 14297 1351 14331
rect 2145 14297 2179 14331
rect 2421 14297 2455 14331
rect 9689 14297 9723 14331
rect 9965 14297 9999 14331
rect 12541 14297 12575 14331
rect 13553 14297 13587 14331
rect 1869 14229 1903 14263
rect 4721 14229 4755 14263
rect 4997 14229 5031 14263
rect 6285 14229 6319 14263
rect 10241 14229 10275 14263
rect 12357 14229 12391 14263
rect 13921 14229 13955 14263
rect 14105 14229 14139 14263
rect 14289 14229 14323 14263
rect 14841 14229 14875 14263
rect 17969 14229 18003 14263
rect 22477 14229 22511 14263
rect 22661 14229 22695 14263
rect 22845 14229 22879 14263
rect 23029 14229 23063 14263
rect 23305 14229 23339 14263
rect 23489 14229 23523 14263
rect 24593 14229 24627 14263
rect 24685 14229 24719 14263
rect 24869 14229 24903 14263
rect 27997 14229 28031 14263
rect 28549 14229 28583 14263
rect 29101 14229 29135 14263
rect 1501 14025 1535 14059
rect 4353 14025 4387 14059
rect 6469 14025 6503 14059
rect 6745 14025 6779 14059
rect 12909 14025 12943 14059
rect 13829 14025 13863 14059
rect 14289 14025 14323 14059
rect 15761 14025 15795 14059
rect 16405 14025 16439 14059
rect 17325 14025 17359 14059
rect 18889 14025 18923 14059
rect 20177 14025 20211 14059
rect 20637 14025 20671 14059
rect 22109 14025 22143 14059
rect 23121 14025 23155 14059
rect 23213 14025 23247 14059
rect 24041 14025 24075 14059
rect 26801 14025 26835 14059
rect 27629 14025 27663 14059
rect 27905 14025 27939 14059
rect 29377 14025 29411 14059
rect 3065 13957 3099 13991
rect 7941 13957 7975 13991
rect 9781 13957 9815 13991
rect 15945 13957 15979 13991
rect 19073 13957 19107 13991
rect 19441 13957 19475 13991
rect 19533 13957 19567 13991
rect 20453 13957 20487 13991
rect 21281 13957 21315 13991
rect 23029 13957 23063 13991
rect 24593 13957 24627 13991
rect 27077 13957 27111 13991
rect 1225 13889 1259 13923
rect 1685 13889 1719 13923
rect 5365 13889 5399 13923
rect 8401 13889 8435 13923
rect 14841 13889 14875 13923
rect 19625 13889 19659 13923
rect 27353 13889 27387 13923
rect 1317 13821 1351 13855
rect 1409 13821 1443 13855
rect 1952 13821 1986 13855
rect 4169 13831 4203 13865
rect 4261 13821 4295 13855
rect 4537 13821 4571 13855
rect 4629 13821 4663 13855
rect 4813 13821 4847 13855
rect 4905 13821 4939 13855
rect 5273 13821 5307 13855
rect 5641 13821 5675 13855
rect 5917 13821 5951 13855
rect 6377 13821 6411 13855
rect 6829 13815 6863 13849
rect 6929 13821 6963 13855
rect 7481 13821 7515 13855
rect 7665 13821 7699 13855
rect 7757 13821 7791 13855
rect 7849 13823 7883 13857
rect 9873 13821 9907 13855
rect 11621 13821 11655 13855
rect 13277 13821 13311 13855
rect 13369 13821 13403 13855
rect 15300 13799 15334 13833
rect 19717 13821 19751 13855
rect 19901 13821 19935 13855
rect 21005 13821 21039 13855
rect 21097 13821 21131 13855
rect 21465 13821 21499 13855
rect 21649 13821 21683 13855
rect 21741 13821 21775 13855
rect 22753 13821 22787 13855
rect 23489 13821 23523 13855
rect 25717 13821 25751 13855
rect 25973 13821 26007 13855
rect 26065 13821 26099 13855
rect 26157 13821 26191 13855
rect 26433 13821 26467 13855
rect 26709 13821 26743 13855
rect 26985 13821 27019 13855
rect 27261 13821 27295 13855
rect 27537 13821 27571 13855
rect 27997 13821 28031 13855
rect 29009 13821 29043 13855
rect 29469 13821 29503 13855
rect 15807 13787 15841 13821
rect 24087 13787 24121 13821
rect 8646 13753 8680 13787
rect 10140 13753 10174 13787
rect 11805 13753 11839 13787
rect 12633 13753 12667 13787
rect 12725 13753 12759 13787
rect 12941 13753 12975 13787
rect 13645 13753 13679 13787
rect 14105 13753 14139 13787
rect 14321 13753 14355 13787
rect 14999 13753 15033 13787
rect 15092 13753 15126 13787
rect 15209 13753 15243 13787
rect 15485 13753 15519 13787
rect 15577 13753 15611 13787
rect 16221 13753 16255 13787
rect 17509 13753 17543 13787
rect 18705 13753 18739 13787
rect 20361 13753 20395 13787
rect 20621 13753 20655 13787
rect 20821 13753 20855 13787
rect 21925 13753 21959 13787
rect 23857 13753 23891 13787
rect 4077 13685 4111 13719
rect 5733 13685 5767 13719
rect 6009 13685 6043 13719
rect 7021 13685 7055 13719
rect 7389 13685 7423 13719
rect 11253 13685 11287 13719
rect 11529 13685 11563 13719
rect 13093 13685 13127 13719
rect 13845 13685 13879 13719
rect 14013 13685 14047 13719
rect 14473 13685 14507 13719
rect 16426 13685 16460 13719
rect 16589 13685 16623 13719
rect 17141 13685 17175 13719
rect 17309 13685 17343 13719
rect 18905 13685 18939 13719
rect 19165 13685 19199 13719
rect 19993 13685 20027 13719
rect 20161 13685 20195 13719
rect 22130 13685 22164 13719
rect 22293 13685 22327 13719
rect 23397 13685 23431 13719
rect 24225 13685 24259 13719
rect 26525 13685 26559 13719
rect 29101 13685 29135 13719
rect 1133 13481 1167 13515
rect 4077 13481 4111 13515
rect 4905 13481 4939 13515
rect 5181 13481 5215 13515
rect 9873 13481 9907 13515
rect 10149 13481 10183 13515
rect 13921 13481 13955 13515
rect 16773 13481 16807 13515
rect 23489 13481 23523 13515
rect 24593 13481 24627 13515
rect 24869 13481 24903 13515
rect 26525 13481 26559 13515
rect 26801 13481 26835 13515
rect 28457 13481 28491 13515
rect 8125 13413 8159 13447
rect 11713 13413 11747 13447
rect 11929 13413 11963 13447
rect 17877 13413 17911 13447
rect 17969 13413 18003 13447
rect 18949 13413 18983 13447
rect 19165 13413 19199 13447
rect 19809 13413 19843 13447
rect 28098 13413 28132 13447
rect 29570 13413 29604 13447
rect 1041 13345 1075 13379
rect 1317 13345 1351 13379
rect 1941 13345 1975 13379
rect 4169 13345 4203 13379
rect 4445 13345 4479 13379
rect 4537 13345 4571 13379
rect 4813 13345 4847 13379
rect 5089 13345 5123 13379
rect 5825 13345 5859 13379
rect 6081 13345 6115 13379
rect 7297 13345 7331 13379
rect 8493 13345 8527 13379
rect 9689 13345 9723 13379
rect 9965 13345 9999 13379
rect 10057 13345 10091 13379
rect 11621 13345 11655 13379
rect 12173 13345 12207 13379
rect 13185 13345 13219 13379
rect 13369 13345 13403 13379
rect 14105 13345 14139 13379
rect 14289 13345 14323 13379
rect 14565 13345 14599 13379
rect 16681 13345 16715 13379
rect 16957 13345 16991 13379
rect 17049 13345 17083 13379
rect 17601 13345 17635 13379
rect 17694 13345 17728 13379
rect 18066 13345 18100 13379
rect 19441 13345 19475 13379
rect 20545 13345 20579 13379
rect 21465 13345 21499 13379
rect 22376 13345 22410 13379
rect 24501 13345 24535 13379
rect 24961 13345 24995 13379
rect 25237 13345 25271 13379
rect 25329 13345 25363 13379
rect 26433 13345 26467 13379
rect 26709 13345 26743 13379
rect 28365 13345 28399 13379
rect 1685 13277 1719 13311
rect 4629 13277 4663 13311
rect 8401 13277 8435 13311
rect 13001 13277 13035 13311
rect 19257 13277 19291 13311
rect 21281 13277 21315 13311
rect 22109 13277 22143 13311
rect 26065 13277 26099 13311
rect 29837 13277 29871 13311
rect 3065 13209 3099 13243
rect 13553 13209 13587 13243
rect 14473 13209 14507 13243
rect 18797 13209 18831 13243
rect 19625 13209 19659 13243
rect 1409 13141 1443 13175
rect 4353 13141 4387 13175
rect 7205 13141 7239 13175
rect 9597 13141 9631 13175
rect 11529 13141 11563 13175
rect 11897 13141 11931 13175
rect 12081 13141 12115 13175
rect 13461 13141 13495 13175
rect 13645 13141 13679 13175
rect 14381 13141 14415 13175
rect 14841 13141 14875 13175
rect 17141 13141 17175 13175
rect 17417 13141 17451 13175
rect 18245 13141 18279 13175
rect 18981 13141 19015 13175
rect 21649 13141 21683 13175
rect 25145 13141 25179 13175
rect 26985 13141 27019 13175
rect 4445 12937 4479 12971
rect 9321 12937 9355 12971
rect 11989 12937 12023 12971
rect 13185 12937 13219 12971
rect 14013 12937 14047 12971
rect 14289 12937 14323 12971
rect 16703 12937 16737 12971
rect 18889 12937 18923 12971
rect 19257 12937 19291 12971
rect 24777 12937 24811 12971
rect 25053 12937 25087 12971
rect 30757 12937 30791 12971
rect 13369 12869 13403 12903
rect 13829 12869 13863 12903
rect 19717 12869 19751 12903
rect 9873 12801 9907 12835
rect 21465 12801 21499 12835
rect 23213 12801 23247 12835
rect 1041 12733 1075 12767
rect 1133 12733 1167 12767
rect 1317 12733 1351 12767
rect 1685 12733 1719 12767
rect 4261 12733 4295 12767
rect 4353 12733 4387 12767
rect 4629 12733 4663 12767
rect 6101 12733 6135 12767
rect 6193 12733 6227 12767
rect 6469 12733 6503 12767
rect 7849 12733 7883 12767
rect 8125 12733 8159 12767
rect 9229 12733 9263 12767
rect 9689 12733 9723 12767
rect 12449 12733 12483 12767
rect 13553 12733 13587 12767
rect 13737 12733 13771 12767
rect 13921 12733 13955 12767
rect 14933 12733 14967 12767
rect 15200 12733 15234 12767
rect 17647 12733 17681 12767
rect 17785 12733 17819 12767
rect 17877 12733 17911 12767
rect 18005 12733 18039 12767
rect 18153 12733 18187 12767
rect 19257 12733 19291 12767
rect 19441 12733 19475 12767
rect 19533 12733 19567 12767
rect 19809 12733 19843 12767
rect 20177 12733 20211 12767
rect 20453 12733 20487 12767
rect 20545 12733 20579 12767
rect 20913 12733 20947 12767
rect 21166 12733 21200 12767
rect 22957 12733 22991 12767
rect 24041 12733 24075 12767
rect 24409 12733 24443 12767
rect 24869 12733 24903 12767
rect 24961 12733 24995 12767
rect 26709 12733 26743 12767
rect 29009 12733 29043 12767
rect 29377 12733 29411 12767
rect 29633 12733 29667 12767
rect 1930 12665 1964 12699
rect 6009 12665 6043 12699
rect 7205 12665 7239 12699
rect 9597 12665 9631 12699
rect 10118 12665 10152 12699
rect 11805 12665 11839 12699
rect 13001 12665 13035 12699
rect 16497 12665 16531 12699
rect 16697 12665 16731 12699
rect 18797 12665 18831 12699
rect 24133 12665 24167 12699
rect 24501 12665 24535 12699
rect 26442 12665 26476 12699
rect 26801 12665 26835 12699
rect 27537 12665 27571 12699
rect 1409 12597 1443 12631
rect 3065 12597 3099 12631
rect 4169 12597 4203 12631
rect 4721 12597 4755 12631
rect 6285 12597 6319 12631
rect 7757 12597 7791 12631
rect 8033 12597 8067 12631
rect 11253 12597 11287 12631
rect 12015 12597 12049 12631
rect 12173 12597 12207 12631
rect 12357 12597 12391 12631
rect 13201 12597 13235 12631
rect 16313 12597 16347 12631
rect 16865 12597 16899 12631
rect 17509 12597 17543 12631
rect 19993 12597 20027 12631
rect 21833 12597 21867 12631
rect 25329 12597 25363 12631
rect 29101 12597 29135 12631
rect 1777 12393 1811 12427
rect 3985 12393 4019 12427
rect 5641 12393 5675 12427
rect 6837 12393 6871 12427
rect 9413 12393 9447 12427
rect 9965 12393 9999 12427
rect 12265 12393 12299 12427
rect 18061 12393 18095 12427
rect 23397 12393 23431 12427
rect 23581 12393 23615 12427
rect 6469 12325 6503 12359
rect 6561 12325 6595 12359
rect 7634 12325 7668 12359
rect 11989 12325 12023 12359
rect 13001 12325 13035 12359
rect 13201 12325 13235 12359
rect 14381 12325 14415 12359
rect 17575 12325 17609 12359
rect 17785 12325 17819 12359
rect 23029 12325 23063 12359
rect 23121 12325 23155 12359
rect 25513 12325 25547 12359
rect 1593 12247 1627 12281
rect 1869 12257 1903 12291
rect 1961 12257 1995 12291
rect 3893 12257 3927 12291
rect 4528 12257 4562 12291
rect 6193 12257 6227 12291
rect 6286 12257 6320 12291
rect 6699 12257 6733 12291
rect 7197 12255 7231 12289
rect 9321 12257 9355 12291
rect 9597 12257 9631 12291
rect 9689 12257 9723 12291
rect 9873 12257 9907 12291
rect 10149 12257 10183 12291
rect 11897 12257 11931 12291
rect 12173 12257 12207 12291
rect 14197 12257 14231 12291
rect 15301 12257 15335 12291
rect 15449 12257 15483 12291
rect 15577 12257 15611 12291
rect 15669 12257 15703 12291
rect 15807 12257 15841 12291
rect 16957 12257 16991 12291
rect 17141 12257 17175 12291
rect 17325 12257 17359 12291
rect 17693 12257 17727 12291
rect 17877 12257 17911 12291
rect 19349 12257 19383 12291
rect 19441 12257 19475 12291
rect 19625 12257 19659 12291
rect 19993 12257 20027 12291
rect 20246 12257 20280 12291
rect 22661 12257 22695 12291
rect 22753 12257 22787 12291
rect 22846 12257 22880 12291
rect 23218 12257 23252 12291
rect 23489 12257 23523 12291
rect 24041 12257 24075 12291
rect 24133 12257 24167 12291
rect 24317 12257 24351 12291
rect 24685 12257 24719 12291
rect 24938 12257 24972 12291
rect 28017 12257 28051 12291
rect 28273 12257 28307 12291
rect 29570 12257 29604 12291
rect 29837 12257 29871 12291
rect 29929 12257 29963 12291
rect 2053 12189 2087 12223
rect 4261 12189 4295 12223
rect 7389 12189 7423 12223
rect 10241 12189 10275 12223
rect 14013 12189 14047 12223
rect 17417 12189 17451 12223
rect 20545 12189 20579 12223
rect 8769 12121 8803 12155
rect 15945 12121 15979 12155
rect 22569 12121 22603 12155
rect 26893 12121 26927 12155
rect 28457 12121 28491 12155
rect 1501 12053 1535 12087
rect 7113 12053 7147 12087
rect 13185 12053 13219 12087
rect 13369 12053 13403 12087
rect 16589 12053 16623 12087
rect 16865 12053 16899 12087
rect 17049 12053 17083 12087
rect 30021 12053 30055 12087
rect 1225 11849 1259 11883
rect 9413 11849 9447 11883
rect 9689 11849 9723 11883
rect 14657 11849 14691 11883
rect 16589 11849 16623 11883
rect 18061 11849 18095 11883
rect 26157 11849 26191 11883
rect 28365 11849 28399 11883
rect 28641 11849 28675 11883
rect 29561 11849 29595 11883
rect 4813 11781 4847 11815
rect 11805 11781 11839 11815
rect 17049 11781 17083 11815
rect 23029 11781 23063 11815
rect 23949 11781 23983 11815
rect 24685 11781 24719 11815
rect 949 11713 983 11747
rect 1685 11713 1719 11747
rect 3433 11713 3467 11747
rect 16773 11713 16807 11747
rect 18153 11713 18187 11747
rect 20085 11713 20119 11747
rect 21649 11713 21683 11747
rect 23581 11713 23615 11747
rect 24593 11713 24627 11747
rect 1041 11645 1075 11679
rect 1133 11645 1167 11679
rect 1409 11645 1443 11679
rect 3700 11645 3734 11679
rect 5641 11645 5675 11679
rect 5734 11645 5768 11679
rect 5917 11645 5951 11679
rect 6009 11645 6043 11679
rect 6147 11645 6181 11679
rect 7481 11645 7515 11679
rect 7574 11645 7608 11679
rect 7849 11645 7883 11679
rect 7987 11645 8021 11679
rect 9229 11645 9263 11679
rect 9321 11645 9355 11679
rect 9781 11645 9815 11679
rect 9965 11645 9999 11679
rect 11897 11645 11931 11679
rect 11989 11645 12023 11679
rect 13553 11645 13587 11679
rect 13737 11645 13771 11679
rect 13829 11645 13863 11679
rect 13921 11645 13955 11679
rect 14841 11645 14875 11679
rect 15025 11645 15059 11679
rect 15143 11645 15177 11679
rect 15301 11645 15335 11679
rect 16865 11645 16899 11679
rect 18061 11645 18095 11679
rect 18337 11645 18371 11679
rect 18705 11645 18739 11679
rect 18889 11645 18923 11679
rect 19073 11645 19107 11679
rect 19441 11645 19475 11679
rect 19694 11645 19728 11679
rect 20361 11645 20395 11679
rect 20545 11645 20579 11679
rect 20729 11645 20763 11679
rect 21097 11645 21131 11679
rect 21350 11645 21384 11679
rect 22109 11645 22143 11679
rect 22201 11645 22235 11679
rect 22477 11645 22511 11679
rect 22569 11645 22603 11679
rect 22845 11645 22879 11679
rect 22937 11645 22971 11679
rect 23213 11645 23247 11679
rect 23305 11645 23339 11679
rect 23673 11645 23707 11679
rect 24133 11645 24167 11679
rect 24317 11645 24351 11679
rect 26065 11645 26099 11679
rect 27537 11645 27571 11679
rect 28273 11645 28307 11679
rect 28733 11645 28767 11679
rect 29009 11645 29043 11679
rect 29469 11645 29503 11679
rect 30941 11645 30975 11679
rect 1930 11577 1964 11611
rect 7757 11577 7791 11611
rect 10232 11577 10266 11611
rect 12256 11577 12290 11611
rect 14933 11577 14967 11611
rect 16589 11577 16623 11611
rect 24225 11577 24259 11611
rect 24455 11577 24489 11611
rect 25820 11577 25854 11611
rect 27270 11577 27304 11611
rect 30674 11577 30708 11611
rect 1501 11509 1535 11543
rect 3065 11509 3099 11543
rect 6285 11509 6319 11543
rect 8125 11509 8159 11543
rect 9137 11509 9171 11543
rect 11345 11509 11379 11543
rect 13369 11509 13403 11543
rect 14105 11509 14139 11543
rect 18521 11509 18555 11543
rect 22753 11509 22787 11543
rect 29101 11509 29135 11543
rect 29377 11509 29411 11543
rect 6469 11305 6503 11339
rect 9045 11305 9079 11339
rect 16221 11305 16255 11339
rect 17325 11305 17359 11339
rect 23029 11305 23063 11339
rect 27261 11305 27295 11339
rect 28365 11305 28399 11339
rect 29193 11305 29227 11339
rect 29561 11305 29595 11339
rect 5365 11237 5399 11271
rect 5457 11237 5491 11271
rect 6193 11237 6227 11271
rect 7288 11237 7322 11271
rect 8769 11237 8803 11271
rect 14442 11237 14476 11271
rect 16957 11237 16991 11271
rect 20576 11237 20610 11271
rect 1317 11169 1351 11203
rect 1573 11169 1607 11203
rect 3341 11169 3375 11203
rect 3608 11169 3642 11203
rect 5273 11169 5307 11203
rect 5641 11169 5675 11203
rect 5825 11169 5859 11203
rect 5918 11169 5952 11203
rect 6101 11169 6135 11203
rect 6331 11169 6365 11203
rect 8493 11169 8527 11203
rect 8677 11169 8711 11203
rect 8861 11169 8895 11203
rect 9413 11169 9447 11203
rect 9689 11169 9723 11203
rect 9965 11169 9999 11203
rect 10241 11169 10275 11203
rect 10517 11169 10551 11203
rect 10793 11169 10827 11203
rect 11253 11169 11287 11203
rect 11437 11169 11471 11203
rect 11529 11169 11563 11203
rect 11897 11169 11931 11203
rect 12165 11169 12199 11203
rect 12449 11169 12483 11203
rect 12541 11169 12575 11203
rect 14197 11169 14231 11203
rect 16405 11169 16439 11203
rect 16589 11169 16623 11203
rect 16681 11169 16715 11203
rect 16819 11169 16853 11203
rect 17049 11169 17083 11203
rect 17187 11169 17221 11203
rect 17417 11169 17451 11203
rect 17601 11169 17635 11203
rect 17877 11169 17911 11203
rect 18153 11169 18187 11203
rect 18406 11169 18440 11203
rect 20821 11169 20855 11203
rect 22394 11169 22428 11203
rect 22661 11169 22695 11203
rect 22753 11169 22787 11203
rect 24153 11169 24187 11203
rect 24409 11169 24443 11203
rect 25513 11169 25547 11203
rect 26893 11169 26927 11203
rect 27169 11169 27203 11203
rect 27445 11169 27479 11203
rect 27905 11169 27939 11203
rect 28181 11169 28215 11203
rect 28273 11169 28307 11203
rect 28549 11169 28583 11203
rect 28825 11169 28859 11203
rect 29101 11169 29135 11203
rect 30674 11169 30708 11203
rect 30941 11169 30975 11203
rect 7021 11101 7055 11135
rect 10701 11101 10735 11135
rect 11805 11101 11839 11135
rect 12357 11101 12391 11135
rect 12633 11101 12667 11135
rect 18705 11101 18739 11135
rect 22845 11101 22879 11135
rect 26985 11101 27019 11135
rect 5089 11033 5123 11067
rect 8401 11033 8435 11067
rect 9321 11033 9355 11067
rect 9597 11033 9631 11067
rect 9873 11033 9907 11067
rect 11161 11033 11195 11067
rect 15577 11033 15611 11067
rect 27537 11033 27571 11067
rect 27813 11033 27847 11067
rect 28089 11033 28123 11067
rect 2697 10965 2731 10999
rect 4721 10965 4755 10999
rect 10149 10965 10183 10999
rect 10425 10965 10459 10999
rect 12081 10965 12115 10999
rect 19441 10965 19475 10999
rect 21281 10965 21315 10999
rect 25605 10965 25639 10999
rect 28641 10965 28675 10999
rect 28917 10965 28951 10999
rect 1593 10761 1627 10795
rect 5549 10761 5583 10795
rect 9873 10761 9907 10795
rect 12725 10761 12759 10795
rect 14289 10761 14323 10795
rect 14749 10761 14783 10795
rect 15209 10761 15243 10795
rect 15669 10761 15703 10795
rect 16589 10761 16623 10795
rect 16865 10761 16899 10795
rect 17509 10761 17543 10795
rect 18337 10761 18371 10795
rect 20361 10761 20395 10795
rect 21465 10761 21499 10795
rect 25053 10761 25087 10795
rect 25697 10761 25731 10795
rect 25973 10761 26007 10795
rect 26433 10761 26467 10795
rect 27261 10761 27295 10795
rect 27813 10761 27847 10795
rect 28089 10761 28123 10795
rect 28365 10761 28399 10795
rect 28733 10761 28767 10795
rect 29469 10761 29503 10795
rect 15853 10693 15887 10727
rect 18889 10693 18923 10727
rect 10701 10625 10735 10659
rect 22293 10625 22327 10659
rect 30481 10625 30515 10659
rect 1685 10557 1719 10591
rect 1777 10557 1811 10591
rect 2053 10557 2087 10591
rect 4261 10557 4295 10591
rect 4997 10557 5031 10591
rect 5273 10557 5307 10591
rect 5365 10557 5399 10591
rect 6653 10557 6687 10591
rect 8401 10557 8435 10591
rect 8585 10557 8619 10591
rect 8769 10557 8803 10591
rect 9505 10557 9539 10591
rect 9597 10557 9631 10591
rect 9965 10557 9999 10591
rect 10333 10557 10367 10591
rect 10793 10557 10827 10591
rect 15945 10557 15979 10591
rect 16038 10557 16072 10591
rect 16313 10557 16347 10591
rect 16410 10557 16444 10591
rect 18705 10557 18739 10591
rect 19717 10557 19751 10591
rect 19810 10557 19844 10591
rect 20085 10557 20119 10591
rect 20223 10557 20257 10591
rect 21373 10557 21407 10591
rect 21649 10557 21683 10591
rect 21925 10557 21959 10591
rect 22560 10557 22594 10591
rect 25145 10557 25179 10591
rect 25513 10557 25547 10591
rect 25789 10557 25823 10591
rect 25881 10557 25915 10591
rect 26341 10557 26375 10591
rect 26617 10557 26651 10591
rect 27077 10557 27111 10591
rect 27169 10557 27203 10591
rect 27629 10557 27663 10591
rect 27721 10557 27755 10591
rect 27997 10557 28031 10591
rect 28457 10557 28491 10591
rect 28825 10557 28859 10591
rect 29101 10557 29135 10591
rect 29193 10557 29227 10591
rect 29377 10557 29411 10591
rect 29745 10557 29779 10591
rect 29837 10557 29871 10591
rect 30941 10557 30975 10591
rect 5181 10489 5215 10523
rect 6920 10489 6954 10523
rect 8677 10489 8711 10523
rect 12541 10489 12575 10523
rect 12757 10489 12791 10523
rect 14473 10489 14507 10523
rect 14565 10489 14599 10523
rect 14765 10489 14799 10523
rect 15025 10489 15059 10523
rect 15485 10489 15519 10523
rect 16221 10489 16255 10523
rect 16681 10489 16715 10523
rect 16897 10489 16931 10523
rect 17601 10489 17635 10523
rect 18153 10489 18187 10523
rect 19993 10489 20027 10523
rect 21741 10489 21775 10523
rect 26709 10489 26743 10523
rect 26985 10489 27019 10523
rect 1869 10421 1903 10455
rect 2145 10421 2179 10455
rect 4169 10421 4203 10455
rect 8033 10421 8067 10455
rect 8953 10421 8987 10455
rect 10241 10421 10275 10455
rect 12909 10421 12943 10455
rect 14105 10421 14139 10455
rect 14273 10421 14307 10455
rect 14933 10421 14967 10455
rect 15225 10421 15259 10455
rect 15393 10421 15427 10455
rect 15695 10421 15729 10455
rect 17049 10421 17083 10455
rect 18358 10421 18392 10455
rect 18521 10421 18555 10455
rect 22017 10421 22051 10455
rect 23673 10421 23707 10455
rect 27537 10421 27571 10455
rect 19625 10217 19659 10251
rect 21557 10217 21591 10251
rect 21833 10217 21867 10251
rect 22109 10217 22143 10251
rect 22937 10217 22971 10251
rect 23857 10217 23891 10251
rect 26893 10217 26927 10251
rect 30941 10217 30975 10251
rect 3709 10149 3743 10183
rect 4537 10149 4571 10183
rect 4813 10149 4847 10183
rect 9588 10149 9622 10183
rect 13369 10149 13403 10183
rect 13585 10149 13619 10183
rect 16129 10149 16163 10183
rect 22385 10149 22419 10183
rect 25513 10149 25547 10183
rect 28006 10149 28040 10183
rect 28917 10149 28951 10183
rect 29644 10149 29678 10183
rect 1225 10081 1259 10115
rect 1501 10081 1535 10115
rect 1869 10081 1903 10115
rect 2125 10081 2159 10115
rect 3341 10081 3375 10115
rect 3433 10081 3467 10115
rect 3801 10081 3835 10115
rect 3893 10081 3927 10115
rect 4169 10081 4203 10115
rect 4445 10081 4479 10115
rect 4721 10081 4755 10115
rect 7205 10081 7239 10115
rect 7665 10081 7699 10115
rect 9321 10081 9355 10115
rect 11897 10081 11931 10115
rect 12153 10081 12187 10115
rect 14013 10081 14047 10115
rect 14197 10081 14231 10115
rect 14289 10081 14323 10115
rect 15393 10081 15427 10115
rect 15577 10081 15611 10115
rect 17969 10081 18003 10115
rect 18153 10081 18187 10115
rect 18337 10081 18371 10115
rect 18705 10081 18739 10115
rect 18958 10081 18992 10115
rect 19533 10081 19567 10115
rect 20749 10081 20783 10115
rect 21005 10081 21039 10115
rect 21649 10081 21683 10115
rect 21741 10081 21775 10115
rect 22201 10081 22235 10115
rect 22293 10081 22327 10115
rect 22569 10081 22603 10115
rect 22845 10081 22879 10115
rect 23581 10081 23615 10115
rect 23949 10081 23983 10115
rect 25421 10081 25455 10115
rect 25789 10081 25823 10115
rect 28733 10081 28767 10115
rect 28825 10081 28859 10115
rect 29285 10081 29319 10115
rect 30849 10081 30883 10115
rect 15117 10013 15151 10047
rect 15209 10013 15243 10047
rect 25697 10013 25731 10047
rect 28273 10013 28307 10047
rect 29377 10013 29411 10047
rect 3985 9945 4019 9979
rect 4261 9945 4295 9979
rect 10701 9945 10735 9979
rect 13277 9945 13311 9979
rect 17417 9945 17451 9979
rect 23213 9945 23247 9979
rect 23489 9945 23523 9979
rect 1317 9877 1351 9911
rect 1593 9877 1627 9911
rect 3249 9877 3283 9911
rect 7297 9877 7331 9911
rect 7573 9877 7607 9911
rect 13553 9877 13587 9911
rect 13737 9877 13771 9911
rect 14381 9877 14415 9911
rect 14473 9877 14507 9911
rect 14749 9877 14783 9911
rect 14841 9877 14875 9911
rect 15301 9877 15335 9911
rect 22661 9877 22695 9911
rect 23673 9877 23707 9911
rect 28641 9877 28675 9911
rect 29193 9877 29227 9911
rect 30757 9877 30791 9911
rect 1869 9673 1903 9707
rect 3801 9673 3835 9707
rect 4077 9673 4111 9707
rect 4353 9673 4387 9707
rect 13829 9673 13863 9707
rect 14657 9673 14691 9707
rect 15117 9673 15151 9707
rect 16589 9673 16623 9707
rect 16681 9673 16715 9707
rect 16957 9673 16991 9707
rect 17141 9673 17175 9707
rect 17509 9673 17543 9707
rect 19165 9673 19199 9707
rect 22109 9673 22143 9707
rect 22661 9673 22695 9707
rect 30021 9673 30055 9707
rect 30297 9673 30331 9707
rect 7573 9605 7607 9639
rect 12817 9605 12851 9639
rect 14013 9605 14047 9639
rect 15577 9605 15611 9639
rect 19625 9605 19659 9639
rect 21189 9605 21223 9639
rect 21833 9605 21867 9639
rect 29101 9605 29135 9639
rect 29653 9605 29687 9639
rect 12633 9537 12667 9571
rect 13921 9537 13955 9571
rect 14749 9537 14783 9571
rect 15209 9537 15243 9571
rect 20177 9537 20211 9571
rect 25697 9537 25731 9571
rect 30573 9537 30607 9571
rect 1409 9469 1443 9503
rect 1593 9469 1627 9503
rect 1685 9469 1719 9503
rect 1777 9469 1811 9503
rect 2053 9469 2087 9503
rect 2329 9469 2363 9503
rect 3525 9469 3559 9503
rect 3893 9469 3927 9503
rect 4169 9469 4203 9503
rect 4261 9469 4295 9503
rect 4905 9469 4939 9503
rect 5161 9469 5195 9503
rect 6837 9469 6871 9503
rect 6929 9469 6963 9503
rect 7389 9469 7423 9503
rect 7665 9469 7699 9503
rect 7757 9469 7791 9503
rect 8033 9469 8067 9503
rect 8401 9469 8435 9503
rect 8657 9469 8691 9503
rect 10885 9469 10919 9503
rect 11152 9469 11186 9503
rect 12357 9469 12391 9503
rect 12725 9469 12759 9503
rect 13553 9469 13587 9503
rect 14841 9469 14875 9503
rect 15393 9469 15427 9503
rect 15952 9469 15986 9503
rect 16038 9469 16072 9503
rect 16310 9469 16344 9503
rect 16429 9469 16463 9503
rect 17049 9469 17083 9503
rect 17417 9469 17451 9503
rect 17693 9469 17727 9503
rect 17785 9469 17819 9503
rect 19349 9469 19383 9503
rect 19441 9469 19475 9503
rect 19717 9469 19751 9503
rect 19993 9469 20027 9503
rect 20085 9469 20119 9503
rect 20269 9469 20303 9503
rect 20453 9469 20487 9503
rect 20545 9469 20579 9503
rect 20638 9469 20672 9503
rect 20913 9469 20947 9503
rect 21010 9469 21044 9503
rect 21925 9469 21959 9503
rect 22201 9469 22235 9503
rect 22293 9469 22327 9503
rect 22569 9469 22603 9503
rect 24133 9469 24167 9503
rect 24317 9469 24351 9503
rect 24501 9469 24535 9503
rect 24869 9469 24903 9503
rect 25122 9469 25156 9503
rect 27169 9469 27203 9503
rect 29193 9469 29227 9503
rect 29469 9469 29503 9503
rect 29745 9469 29779 9503
rect 30113 9469 30147 9503
rect 30389 9469 30423 9503
rect 30481 9469 30515 9503
rect 13093 9401 13127 9435
rect 14565 9401 14599 9435
rect 15117 9401 15151 9435
rect 16221 9401 16255 9435
rect 19165 9401 19199 9435
rect 20821 9401 20855 9435
rect 26902 9401 26936 9435
rect 29377 9401 29411 9435
rect 1317 9333 1351 9367
rect 2145 9333 2179 9367
rect 2421 9333 2455 9367
rect 3433 9333 3467 9367
rect 6285 9333 6319 9367
rect 6745 9333 6779 9367
rect 7021 9333 7055 9367
rect 7297 9333 7331 9367
rect 7849 9333 7883 9367
rect 8125 9333 8159 9367
rect 9781 9333 9815 9367
rect 12265 9333 12299 9367
rect 12449 9333 12483 9367
rect 13645 9333 13679 9367
rect 14289 9333 14323 9367
rect 15025 9333 15059 9367
rect 17279 9333 17313 9367
rect 22385 9333 22419 9367
rect 25789 9333 25823 9367
rect 1317 9129 1351 9163
rect 3249 9129 3283 9163
rect 3801 9129 3835 9163
rect 5641 9129 5675 9163
rect 10241 9129 10275 9163
rect 11529 9129 11563 9163
rect 15025 9129 15059 9163
rect 20545 9129 20579 9163
rect 21925 9129 21959 9163
rect 22201 9129 22235 9163
rect 23857 9129 23891 9163
rect 24593 9129 24627 9163
rect 25027 9129 25061 9163
rect 25487 9129 25521 9163
rect 26525 9129 26559 9163
rect 30941 9129 30975 9163
rect 2697 9061 2731 9095
rect 7297 9061 7331 9095
rect 9106 9061 9140 9095
rect 11161 9061 11195 9095
rect 11377 9061 11411 9095
rect 14381 9061 14415 9095
rect 16405 9061 16439 9095
rect 18505 9061 18539 9095
rect 18705 9061 18739 9095
rect 20039 9061 20073 9095
rect 20177 9061 20211 9095
rect 25237 9061 25271 9095
rect 25697 9061 25731 9095
rect 1133 8993 1167 9027
rect 1409 8993 1443 9027
rect 1685 8993 1719 9027
rect 1961 8993 1995 9027
rect 2145 8993 2179 9027
rect 2237 8993 2271 9027
rect 2605 8993 2639 9027
rect 2881 8993 2915 9027
rect 3157 8993 3191 9027
rect 3433 8993 3467 9027
rect 3893 8993 3927 9027
rect 4077 8993 4111 9027
rect 4169 8993 4203 9027
rect 4517 8993 4551 9027
rect 7113 8993 7147 9027
rect 7389 8993 7423 9027
rect 7665 8993 7699 9027
rect 7757 8993 7791 9027
rect 11805 8993 11839 9027
rect 13001 8993 13035 9027
rect 13185 8993 13219 9027
rect 13277 8993 13311 9027
rect 14657 8993 14691 9027
rect 15117 8993 15151 9027
rect 16313 8993 16347 9027
rect 16497 8993 16531 9027
rect 16635 8993 16669 9027
rect 16773 8993 16807 9027
rect 17141 8993 17175 9027
rect 18061 8993 18095 9027
rect 18245 8993 18279 9027
rect 20269 8993 20303 9027
rect 20361 8993 20395 9027
rect 22017 8993 22051 9027
rect 22109 8993 22143 9027
rect 22733 8993 22767 9027
rect 24685 8993 24719 9027
rect 27649 8993 27683 9027
rect 27905 8993 27939 9027
rect 28365 8993 28399 9027
rect 28825 8993 28859 9027
rect 29101 8993 29135 9027
rect 29377 8993 29411 9027
rect 29561 8993 29595 9027
rect 29817 8993 29851 9027
rect 1593 8925 1627 8959
rect 2973 8925 3007 8959
rect 3525 8925 3559 8959
rect 4261 8925 4295 8959
rect 8861 8925 8895 8959
rect 11989 8925 12023 8959
rect 17509 8925 17543 8959
rect 19901 8925 19935 8959
rect 22477 8925 22511 8959
rect 1041 8857 1075 8891
rect 1869 8857 1903 8891
rect 11621 8857 11655 8891
rect 13461 8857 13495 8891
rect 14749 8857 14783 8891
rect 14841 8857 14875 8891
rect 16129 8857 16163 8891
rect 24225 8857 24259 8891
rect 7021 8789 7055 8823
rect 7573 8789 7607 8823
rect 7849 8789 7883 8823
rect 11345 8789 11379 8823
rect 13277 8789 13311 8823
rect 17325 8789 17359 8823
rect 17785 8789 17819 8823
rect 17877 8789 17911 8823
rect 17969 8789 18003 8823
rect 18337 8789 18371 8823
rect 18521 8789 18555 8823
rect 23949 8789 23983 8823
rect 24317 8789 24351 8823
rect 24409 8789 24443 8823
rect 24869 8789 24903 8823
rect 25053 8789 25087 8823
rect 25329 8789 25363 8823
rect 25513 8789 25547 8823
rect 28457 8789 28491 8823
rect 28733 8789 28767 8823
rect 29009 8789 29043 8823
rect 29285 8789 29319 8823
rect 1685 8585 1719 8619
rect 2145 8585 2179 8619
rect 2421 8585 2455 8619
rect 2697 8585 2731 8619
rect 5825 8585 5859 8619
rect 7113 8585 7147 8619
rect 12541 8585 12575 8619
rect 13001 8585 13035 8619
rect 14289 8585 14323 8619
rect 14565 8585 14599 8619
rect 15209 8585 15243 8619
rect 15853 8585 15887 8619
rect 17049 8585 17083 8619
rect 17233 8585 17267 8619
rect 17693 8585 17727 8619
rect 19717 8585 19751 8619
rect 19993 8585 20027 8619
rect 23489 8585 23523 8619
rect 23673 8585 23707 8619
rect 24317 8585 24351 8619
rect 26525 8585 26559 8619
rect 29377 8585 29411 8619
rect 9781 8517 9815 8551
rect 11805 8517 11839 8551
rect 12633 8517 12667 8551
rect 13921 8517 13955 8551
rect 14013 8517 14047 8551
rect 14749 8517 14783 8551
rect 15301 8517 15335 8551
rect 19349 8517 19383 8551
rect 19809 8517 19843 8551
rect 14933 8449 14967 8483
rect 24225 8449 24259 8483
rect 27905 8449 27939 8483
rect 1593 8381 1627 8415
rect 2053 8381 2087 8415
rect 2513 8381 2547 8415
rect 2605 8381 2639 8415
rect 4445 8381 4479 8415
rect 6377 8381 6411 8415
rect 6561 8381 6595 8415
rect 6653 8381 6687 8415
rect 6929 8381 6963 8415
rect 7021 8381 7055 8415
rect 7481 8381 7515 8415
rect 7573 8381 7607 8415
rect 8401 8381 8435 8415
rect 8657 8381 8691 8415
rect 10425 8381 10459 8415
rect 12265 8381 12299 8415
rect 12449 8381 12483 8415
rect 12725 8381 12759 8415
rect 13553 8381 13587 8415
rect 13829 8381 13863 8415
rect 15393 8381 15427 8415
rect 15485 8381 15519 8415
rect 15672 8381 15706 8415
rect 16037 8381 16071 8415
rect 16221 8381 16255 8415
rect 16681 8381 16715 8415
rect 16865 8381 16899 8415
rect 17417 8381 17451 8415
rect 17509 8381 17543 8415
rect 18981 8381 19015 8415
rect 19165 8381 19199 8415
rect 19257 8381 19291 8415
rect 19441 8381 19475 8415
rect 22385 8381 22419 8415
rect 23857 8381 23891 8415
rect 24133 8381 24167 8415
rect 24593 8381 24627 8415
rect 26249 8381 26283 8415
rect 28825 8381 28859 8415
rect 29193 8381 29227 8415
rect 29469 8381 29503 8415
rect 29745 8381 29779 8415
rect 30021 8381 30055 8415
rect 30113 8381 30147 8415
rect 30573 8381 30607 8415
rect 30665 8381 30699 8415
rect 4712 8313 4746 8347
rect 6285 8313 6319 8347
rect 10670 8313 10704 8347
rect 14381 8313 14415 8347
rect 17233 8313 17267 8347
rect 20177 8313 20211 8347
rect 22118 8313 22152 8347
rect 23305 8313 23339 8347
rect 25982 8313 26016 8347
rect 27660 8313 27694 8347
rect 28733 8313 28767 8347
rect 29929 8313 29963 8347
rect 6837 8245 6871 8279
rect 7389 8245 7423 8279
rect 7665 8245 7699 8279
rect 13645 8245 13679 8279
rect 14581 8245 14615 8279
rect 19967 8245 20001 8279
rect 21005 8245 21039 8279
rect 23505 8245 23539 8279
rect 24501 8245 24535 8279
rect 24869 8245 24903 8279
rect 29101 8245 29135 8279
rect 29653 8245 29687 8279
rect 30205 8245 30239 8279
rect 30481 8245 30515 8279
rect 30757 8245 30791 8279
rect 3617 8041 3651 8075
rect 6193 8041 6227 8075
rect 13185 8041 13219 8075
rect 13645 8041 13679 8075
rect 16129 8041 16163 8075
rect 16681 8041 16715 8075
rect 17785 8041 17819 8075
rect 18613 8041 18647 8075
rect 18781 8041 18815 8075
rect 19349 8041 19383 8075
rect 19517 8041 19551 8075
rect 20269 8041 20303 8075
rect 20437 8041 20471 8075
rect 22017 8041 22051 8075
rect 22293 8041 22327 8075
rect 22569 8041 22603 8075
rect 24409 8041 24443 8075
rect 30941 8041 30975 8075
rect 3954 7973 3988 8007
rect 8094 7973 8128 8007
rect 13277 7973 13311 8007
rect 13477 7973 13511 8007
rect 18981 7973 19015 8007
rect 19717 7973 19751 8007
rect 20177 7973 20211 8007
rect 20637 7973 20671 8007
rect 28917 7973 28951 8007
rect 29806 7973 29840 8007
rect 19947 7939 19981 7973
rect 2504 7905 2538 7939
rect 3709 7905 3743 7939
rect 5641 7905 5675 7939
rect 5825 7905 5859 7939
rect 6285 7905 6319 7939
rect 7297 7905 7331 7939
rect 7573 7905 7607 7939
rect 11233 7905 11267 7939
rect 12449 7905 12483 7939
rect 12633 7905 12667 7939
rect 14013 7905 14047 7939
rect 14197 7905 14231 7939
rect 15301 7895 15335 7929
rect 15485 7905 15519 7939
rect 16865 7905 16899 7939
rect 18153 7905 18187 7939
rect 18521 7905 18555 7939
rect 21557 7905 21591 7939
rect 21649 7905 21683 7939
rect 22109 7905 22143 7939
rect 22385 7905 22419 7939
rect 22477 7905 22511 7939
rect 23285 7905 23319 7939
rect 26249 7905 26283 7939
rect 27822 7905 27856 7939
rect 28089 7905 28123 7939
rect 28733 7905 28767 7939
rect 28825 7905 28859 7939
rect 29101 7905 29135 7939
rect 2237 7837 2271 7871
rect 6561 7837 6595 7871
rect 7849 7837 7883 7871
rect 10977 7837 11011 7871
rect 14381 7837 14415 7871
rect 16589 7837 16623 7871
rect 17049 7837 17083 7871
rect 17325 7837 17359 7871
rect 23029 7837 23063 7871
rect 25421 7837 25455 7871
rect 29561 7837 29595 7871
rect 5089 7769 5123 7803
rect 12357 7769 12391 7803
rect 16313 7769 16347 7803
rect 17601 7769 17635 7803
rect 19809 7769 19843 7803
rect 26709 7769 26743 7803
rect 5549 7701 5583 7735
rect 5917 7701 5951 7735
rect 7481 7701 7515 7735
rect 9229 7701 9263 7735
rect 12725 7701 12759 7735
rect 12817 7701 12851 7735
rect 12909 7701 12943 7735
rect 13461 7701 13495 7735
rect 15117 7701 15151 7735
rect 18797 7701 18831 7735
rect 19533 7701 19567 7735
rect 19993 7701 20027 7735
rect 20453 7701 20487 7735
rect 21465 7701 21499 7735
rect 21741 7701 21775 7735
rect 28641 7701 28675 7735
rect 29193 7701 29227 7735
rect 2513 7497 2547 7531
rect 11621 7497 11655 7531
rect 11805 7497 11839 7531
rect 13093 7497 13127 7531
rect 13277 7497 13311 7531
rect 14565 7497 14599 7531
rect 19165 7497 19199 7531
rect 21649 7497 21683 7531
rect 21925 7497 21959 7531
rect 22201 7497 22235 7531
rect 22477 7497 22511 7531
rect 26157 7497 26191 7531
rect 28549 7497 28583 7531
rect 30297 7497 30331 7531
rect 30941 7497 30975 7531
rect 6285 7429 6319 7463
rect 8125 7429 8159 7463
rect 15301 7429 15335 7463
rect 16497 7429 16531 7463
rect 18061 7429 18095 7463
rect 24685 7429 24719 7463
rect 6745 7361 6779 7395
rect 8953 7361 8987 7395
rect 14933 7361 14967 7395
rect 15853 7361 15887 7395
rect 27537 7361 27571 7395
rect 27997 7361 28031 7395
rect 29101 7361 29135 7395
rect 1133 7293 1167 7327
rect 4169 7293 4203 7327
rect 5825 7293 5859 7327
rect 6009 7293 6043 7327
rect 6101 7293 6135 7327
rect 6377 7293 6411 7327
rect 6469 7293 6503 7327
rect 8861 7293 8895 7327
rect 10425 7293 10459 7327
rect 14289 7293 14323 7327
rect 15945 7293 15979 7327
rect 16037 7293 16071 7327
rect 16681 7293 16715 7327
rect 17233 7293 17267 7327
rect 17325 7293 17359 7327
rect 17417 7293 17451 7327
rect 20289 7293 20323 7327
rect 20545 7293 20579 7327
rect 21189 7295 21223 7329
rect 21465 7293 21499 7327
rect 21557 7293 21591 7327
rect 22017 7293 22051 7327
rect 22293 7293 22327 7327
rect 22385 7293 22419 7327
rect 23673 7293 23707 7327
rect 26065 7293 26099 7327
rect 28089 7293 28123 7327
rect 28733 7293 28767 7327
rect 29193 7293 29227 7327
rect 29469 7293 29503 7327
rect 30473 7293 30507 7327
rect 30573 7293 30607 7327
rect 30849 7293 30883 7327
rect 13139 7259 13173 7293
rect 1400 7225 1434 7259
rect 4436 7225 4470 7259
rect 6990 7225 7024 7259
rect 9198 7225 9232 7259
rect 11161 7225 11195 7259
rect 11437 7225 11471 7259
rect 12909 7225 12943 7259
rect 14381 7225 14415 7259
rect 15117 7225 15151 7259
rect 15485 7225 15519 7259
rect 15669 7225 15703 7259
rect 17785 7225 17819 7259
rect 22937 7225 22971 7259
rect 25820 7225 25854 7259
rect 27292 7225 27326 7259
rect 5549 7157 5583 7191
rect 5733 7157 5767 7191
rect 6561 7157 6595 7191
rect 8769 7157 8803 7191
rect 10333 7157 10367 7191
rect 11637 7157 11671 7191
rect 14105 7157 14139 7191
rect 14581 7157 14615 7191
rect 14749 7157 14783 7191
rect 21097 7157 21131 7191
rect 21373 7157 21407 7191
rect 29285 7157 29319 7191
rect 30665 7157 30699 7191
rect 8677 6953 8711 6987
rect 12751 6953 12785 6987
rect 14749 6953 14783 6987
rect 16589 6953 16623 6987
rect 19517 6953 19551 6987
rect 27537 6953 27571 6987
rect 27813 6953 27847 6987
rect 30113 6953 30147 6987
rect 7297 6885 7331 6919
rect 12541 6885 12575 6919
rect 14565 6885 14599 6919
rect 17417 6885 17451 6919
rect 19717 6885 19751 6919
rect 26433 6885 26467 6919
rect 27261 6885 27295 6919
rect 2145 6817 2179 6851
rect 2401 6817 2435 6851
rect 5825 6817 5859 6851
rect 6285 6817 6319 6851
rect 7481 6817 7515 6851
rect 7573 6817 7607 6851
rect 7665 6817 7699 6851
rect 8309 6817 8343 6851
rect 8585 6817 8619 6851
rect 9045 6817 9079 6851
rect 9321 6817 9355 6851
rect 11233 6817 11267 6851
rect 13645 6817 13679 6851
rect 13829 6817 13863 6851
rect 14197 6817 14231 6851
rect 15209 6817 15243 6851
rect 15301 6817 15335 6851
rect 15485 6817 15519 6851
rect 16221 6817 16255 6851
rect 17693 6817 17727 6851
rect 18153 6817 18187 6851
rect 18521 6817 18555 6851
rect 18981 6817 19015 6851
rect 21557 6817 21591 6851
rect 22017 6817 22051 6851
rect 22293 6817 22327 6851
rect 22569 6817 22603 6851
rect 23958 6817 23992 6851
rect 26249 6817 26283 6851
rect 27629 6817 27663 6851
rect 27905 6817 27939 6851
rect 28273 6817 28307 6851
rect 28457 6817 28491 6851
rect 28733 6817 28767 6851
rect 29101 6817 29135 6851
rect 29745 6817 29779 6851
rect 29837 6817 29871 6851
rect 30205 6817 30239 6851
rect 30849 6817 30883 6851
rect 6561 6749 6595 6783
rect 10977 6749 11011 6783
rect 13093 6749 13127 6783
rect 18889 6749 18923 6783
rect 21925 6749 21959 6783
rect 22477 6749 22511 6783
rect 24225 6749 24259 6783
rect 5917 6681 5951 6715
rect 6193 6681 6227 6715
rect 7757 6681 7791 6715
rect 9413 6681 9447 6715
rect 12357 6681 12391 6715
rect 12909 6681 12943 6715
rect 15025 6681 15059 6715
rect 17601 6681 17635 6715
rect 22201 6681 22235 6715
rect 28549 6681 28583 6715
rect 3525 6613 3559 6647
rect 8401 6613 8435 6647
rect 9137 6613 9171 6647
rect 12725 6613 12759 6647
rect 13369 6613 13403 6647
rect 13461 6613 13495 6647
rect 13553 6613 13587 6647
rect 15117 6613 15151 6647
rect 16589 6613 16623 6647
rect 16773 6613 16807 6647
rect 19349 6613 19383 6647
rect 19533 6613 19567 6647
rect 21649 6613 21683 6647
rect 22845 6613 22879 6647
rect 26157 6613 26191 6647
rect 28181 6613 28215 6647
rect 28825 6613 28859 6647
rect 29285 6613 29319 6647
rect 30665 6613 30699 6647
rect 6193 6409 6227 6443
rect 6561 6409 6595 6443
rect 8493 6409 8527 6443
rect 9597 6409 9631 6443
rect 10517 6409 10551 6443
rect 12909 6409 12943 6443
rect 13093 6409 13127 6443
rect 14013 6409 14047 6443
rect 14289 6409 14323 6443
rect 14565 6409 14599 6443
rect 19441 6409 19475 6443
rect 22109 6409 22143 6443
rect 22937 6409 22971 6443
rect 23213 6409 23247 6443
rect 23489 6409 23523 6443
rect 24225 6409 24259 6443
rect 28733 6409 28767 6443
rect 31033 6409 31067 6443
rect 2513 6341 2547 6375
rect 6837 6341 6871 6375
rect 14749 6341 14783 6375
rect 15945 6341 15979 6375
rect 19073 6341 19107 6375
rect 22661 6341 22695 6375
rect 24501 6341 24535 6375
rect 24777 6341 24811 6375
rect 27813 6341 27847 6375
rect 28089 6341 28123 6375
rect 8217 6273 8251 6307
rect 10977 6273 11011 6307
rect 15669 6273 15703 6307
rect 15761 6273 15795 6307
rect 18705 6273 18739 6307
rect 26433 6273 26467 6307
rect 26709 6273 26743 6307
rect 949 6205 983 6239
rect 1205 6205 1239 6239
rect 2605 6205 2639 6239
rect 2881 6205 2915 6239
rect 3709 6205 3743 6239
rect 4077 6205 4111 6239
rect 4353 6205 4387 6239
rect 4445 6205 4479 6239
rect 6285 6205 6319 6239
rect 6469 6205 6503 6239
rect 7961 6205 7995 6239
rect 8401 6205 8435 6239
rect 8677 6205 8711 6239
rect 8953 6205 8987 6239
rect 9229 6205 9263 6239
rect 9505 6205 9539 6239
rect 9965 6205 9999 6239
rect 10149 6205 10183 6239
rect 10425 6205 10459 6239
rect 10701 6205 10735 6239
rect 13553 6205 13587 6239
rect 13737 6205 13771 6239
rect 13829 6205 13863 6239
rect 13921 6205 13955 6239
rect 15559 6205 15593 6239
rect 17325 6205 17359 6239
rect 17417 6205 17451 6239
rect 17693 6205 17727 6239
rect 17969 6205 18003 6239
rect 18113 6205 18147 6239
rect 18889 6205 18923 6239
rect 20565 6205 20599 6239
rect 20821 6205 20855 6239
rect 21925 6205 21959 6239
rect 22017 6205 22051 6239
rect 22477 6205 22511 6239
rect 22753 6205 22787 6239
rect 22845 6205 22879 6239
rect 23305 6205 23339 6239
rect 23581 6205 23615 6239
rect 24041 6205 24075 6239
rect 24317 6205 24351 6239
rect 24409 6205 24443 6239
rect 24869 6205 24903 6239
rect 24961 6205 24995 6239
rect 25421 6205 25455 6239
rect 25697 6205 25731 6239
rect 25973 6205 26007 6239
rect 26249 6205 26283 6239
rect 26341 6205 26375 6239
rect 26801 6205 26835 6239
rect 27077 6205 27111 6239
rect 27353 6205 27387 6239
rect 27629 6205 27663 6239
rect 27721 6205 27755 6239
rect 28181 6205 28215 6239
rect 28457 6207 28491 6241
rect 28825 6205 28859 6239
rect 29561 6205 29595 6239
rect 29653 6205 29687 6239
rect 29909 6205 29943 6239
rect 12955 6171 12989 6205
rect 4690 6137 4724 6171
rect 8769 6137 8803 6171
rect 9873 6137 9907 6171
rect 10241 6137 10275 6171
rect 10793 6137 10827 6171
rect 11222 6137 11256 6171
rect 12725 6137 12759 6171
rect 14381 6137 14415 6171
rect 14597 6137 14631 6171
rect 17141 6137 17175 6171
rect 17877 6137 17911 6171
rect 21189 6137 21223 6171
rect 25053 6137 25087 6171
rect 25329 6137 25363 6171
rect 25881 6137 25915 6171
rect 26157 6137 26191 6171
rect 26985 6137 27019 6171
rect 27261 6137 27295 6171
rect 27537 6137 27571 6171
rect 2329 6069 2363 6103
rect 2789 6069 2823 6103
rect 3617 6069 3651 6103
rect 3985 6069 4019 6103
rect 4261 6069 4295 6103
rect 5825 6069 5859 6103
rect 9045 6069 9079 6103
rect 9321 6069 9355 6103
rect 12357 6069 12391 6103
rect 17417 6069 17451 6103
rect 18262 6069 18296 6103
rect 22385 6069 22419 6103
rect 23949 6069 23983 6103
rect 25605 6069 25639 6103
rect 28365 6069 28399 6103
rect 29377 6069 29411 6103
rect 2789 5865 2823 5899
rect 4629 5865 4663 5899
rect 4905 5865 4939 5899
rect 7205 5865 7239 5899
rect 10333 5865 10367 5899
rect 14197 5865 14231 5899
rect 19073 5865 19107 5899
rect 19691 5865 19725 5899
rect 20161 5865 20195 5899
rect 20611 5865 20645 5899
rect 23949 5865 23983 5899
rect 25421 5865 25455 5899
rect 28641 5865 28675 5899
rect 29101 5865 29135 5899
rect 30941 5865 30975 5899
rect 5181 5797 5215 5831
rect 12081 5797 12115 5831
rect 14105 5797 14139 5831
rect 15025 5797 15059 5831
rect 18061 5797 18095 5831
rect 19241 5797 19275 5831
rect 19441 5797 19475 5831
rect 19901 5797 19935 5831
rect 20361 5797 20395 5831
rect 20821 5797 20855 5831
rect 23167 5797 23201 5831
rect 1041 5729 1075 5763
rect 1133 5729 1167 5763
rect 1389 5729 1423 5763
rect 2881 5729 2915 5763
rect 3157 5729 3191 5763
rect 3249 5729 3283 5763
rect 3516 5729 3550 5763
rect 4997 5729 5031 5763
rect 5273 5729 5307 5763
rect 5825 5729 5859 5763
rect 6081 5729 6115 5763
rect 7481 5729 7515 5763
rect 7849 5729 7883 5763
rect 9689 5729 9723 5763
rect 9965 5729 9999 5763
rect 10425 5729 10459 5763
rect 12429 5729 12463 5763
rect 14933 5729 14967 5763
rect 15117 5729 15151 5763
rect 16497 5729 16531 5763
rect 16865 5729 16899 5763
rect 17233 5729 17267 5763
rect 17785 5729 17819 5763
rect 21281 5729 21315 5763
rect 21548 5729 21582 5763
rect 23305 5729 23339 5763
rect 23397 5729 23431 5763
rect 23488 5751 23522 5785
rect 23857 5729 23891 5763
rect 24501 5729 24535 5763
rect 24593 5729 24627 5763
rect 24869 5729 24903 5763
rect 25237 5729 25271 5763
rect 25513 5729 25547 5763
rect 26525 5729 26559 5763
rect 26617 5729 26651 5763
rect 28201 5729 28235 5763
rect 28457 5729 28491 5763
rect 28733 5729 28767 5763
rect 29193 5729 29227 5763
rect 30501 5729 30535 5763
rect 30757 5729 30791 5763
rect 30849 5729 30883 5763
rect 949 5661 983 5695
rect 11345 5661 11379 5695
rect 12173 5661 12207 5695
rect 23029 5661 23063 5695
rect 23673 5661 23707 5695
rect 24777 5661 24811 5695
rect 25145 5661 25179 5695
rect 2513 5593 2547 5627
rect 9873 5593 9907 5627
rect 13553 5593 13587 5627
rect 18429 5593 18463 5627
rect 19533 5593 19567 5627
rect 27077 5593 27111 5627
rect 29377 5593 29411 5627
rect 3065 5525 3099 5559
rect 7389 5525 7423 5559
rect 7757 5525 7791 5559
rect 9597 5525 9631 5559
rect 17877 5525 17911 5559
rect 18061 5525 18095 5559
rect 19257 5525 19291 5559
rect 19717 5525 19751 5559
rect 19993 5525 20027 5559
rect 20177 5525 20211 5559
rect 20453 5525 20487 5559
rect 20637 5525 20671 5559
rect 22661 5525 22695 5559
rect 1409 5321 1443 5355
rect 1961 5321 1995 5355
rect 2513 5321 2547 5355
rect 4813 5321 4847 5355
rect 5365 5321 5399 5355
rect 6193 5321 6227 5355
rect 7021 5321 7055 5355
rect 9413 5321 9447 5355
rect 9689 5321 9723 5355
rect 10241 5321 10275 5355
rect 13185 5321 13219 5355
rect 14289 5321 14323 5355
rect 14473 5321 14507 5355
rect 15945 5321 15979 5355
rect 18889 5321 18923 5355
rect 19717 5321 19751 5355
rect 19809 5321 19843 5355
rect 20269 5321 20303 5355
rect 20637 5321 20671 5355
rect 20729 5321 20763 5355
rect 23857 5321 23891 5355
rect 25329 5321 25363 5355
rect 28457 5321 28491 5355
rect 28733 5321 28767 5355
rect 30573 5321 30607 5355
rect 4261 5253 4295 5287
rect 5089 5253 5123 5287
rect 8585 5253 8619 5287
rect 11989 5253 12023 5287
rect 13369 5253 13403 5287
rect 15301 5253 15335 5287
rect 16957 5253 16991 5287
rect 2237 5185 2271 5219
rect 8861 5185 8895 5219
rect 9965 5185 9999 5219
rect 10609 5185 10643 5219
rect 19441 5185 19475 5219
rect 19901 5185 19935 5219
rect 22569 5185 22603 5219
rect 23213 5185 23247 5219
rect 25237 5185 25271 5219
rect 29009 5185 29043 5219
rect 1501 5117 1535 5151
rect 1685 5117 1719 5151
rect 1777 5117 1811 5151
rect 2053 5117 2087 5151
rect 2329 5117 2363 5151
rect 2421 5117 2455 5151
rect 2697 5117 2731 5151
rect 3801 5117 3835 5151
rect 4077 5117 4111 5151
rect 4353 5117 4387 5151
rect 4905 5117 4939 5151
rect 5181 5117 5215 5151
rect 5457 5117 5491 5151
rect 5549 5117 5583 5151
rect 5641 5117 5675 5151
rect 6009 5117 6043 5151
rect 6285 5117 6319 5151
rect 6469 5117 6503 5151
rect 6561 5117 6595 5151
rect 6837 5117 6871 5151
rect 7113 5117 7147 5151
rect 7389 5117 7423 5151
rect 7665 5117 7699 5151
rect 7941 5117 7975 5151
rect 8125 5117 8159 5151
rect 8217 5117 8251 5151
rect 8677 5117 8711 5151
rect 8953 5117 8987 5151
rect 9229 5117 9263 5151
rect 9321 5117 9355 5151
rect 9781 5117 9815 5151
rect 10057 5117 10091 5151
rect 10149 5117 10183 5151
rect 15577 5117 15611 5151
rect 15761 5117 15795 5151
rect 16129 5117 16163 5151
rect 17509 5117 17543 5151
rect 17601 5117 17635 5151
rect 19993 5117 20027 5151
rect 20177 5117 20211 5151
rect 20545 5117 20579 5151
rect 21005 5117 21039 5151
rect 22753 5117 22787 5151
rect 23075 5117 23109 5151
rect 24970 5117 25004 5151
rect 26709 5117 26743 5151
rect 28549 5117 28583 5151
rect 28825 5117 28859 5151
rect 29276 5117 29310 5151
rect 30665 5117 30699 5151
rect 30757 5117 30791 5151
rect 3709 5049 3743 5083
rect 3985 5049 4019 5083
rect 6745 5049 6779 5083
rect 7573 5049 7607 5083
rect 10854 5049 10888 5083
rect 13001 5049 13035 5083
rect 14105 5049 14139 5083
rect 15025 5049 15059 5083
rect 17233 5049 17267 5083
rect 18873 5049 18907 5083
rect 19073 5049 19107 5083
rect 22845 5049 22879 5083
rect 22937 5049 22971 5083
rect 26464 5049 26498 5083
rect 30849 5049 30883 5083
rect 2789 4981 2823 5015
rect 5917 4981 5951 5015
rect 7297 4981 7331 5015
rect 7849 4981 7883 5015
rect 9137 4981 9171 5015
rect 13211 4981 13245 5015
rect 14315 4981 14349 5015
rect 15485 4981 15519 5015
rect 16313 4981 16347 5015
rect 16773 4981 16807 5015
rect 17325 4981 17359 5015
rect 18705 4981 18739 5015
rect 20913 4981 20947 5015
rect 30389 4981 30423 5015
rect 1777 4777 1811 4811
rect 7205 4777 7239 4811
rect 8677 4777 8711 4811
rect 11463 4777 11497 4811
rect 12081 4777 12115 4811
rect 13645 4777 13679 4811
rect 14105 4777 14139 4811
rect 14841 4777 14875 4811
rect 15004 4777 15038 4811
rect 18613 4777 18647 4811
rect 18981 4777 19015 4811
rect 19625 4777 19659 4811
rect 20361 4777 20395 4811
rect 21005 4777 21039 4811
rect 23029 4777 23063 4811
rect 29469 4777 29503 4811
rect 3770 4709 3804 4743
rect 7542 4709 7576 4743
rect 9496 4709 9530 4743
rect 11253 4709 11287 4743
rect 11713 4709 11747 4743
rect 12173 4709 12207 4743
rect 12389 4709 12423 4743
rect 13159 4709 13193 4743
rect 13369 4709 13403 4743
rect 13737 4709 13771 4743
rect 13953 4709 13987 4743
rect 15209 4709 15243 4743
rect 16681 4709 16715 4743
rect 20269 4709 20303 4743
rect 21916 4709 21950 4743
rect 29101 4709 29135 4743
rect 11943 4675 11977 4709
rect 1041 4641 1075 4675
rect 1225 4641 1259 4675
rect 1317 4641 1351 4675
rect 1409 4641 1443 4675
rect 1869 4641 1903 4675
rect 2053 4641 2087 4675
rect 2309 4641 2343 4675
rect 5825 4641 5859 4675
rect 6081 4641 6115 4675
rect 13277 4641 13311 4675
rect 13461 4641 13495 4675
rect 15485 4641 15519 4675
rect 17141 4641 17175 4675
rect 17325 4641 17359 4675
rect 17877 4641 17911 4675
rect 18061 4641 18095 4675
rect 18153 4641 18187 4675
rect 18889 4641 18923 4675
rect 19165 4641 19199 4675
rect 20085 4641 20119 4675
rect 21097 4641 21131 4675
rect 21649 4641 21683 4675
rect 27730 4641 27764 4675
rect 28917 4641 28951 4675
rect 29009 4641 29043 4675
rect 30582 4641 30616 4675
rect 30849 4641 30883 4675
rect 3525 4573 3559 4607
rect 7297 4573 7331 4607
rect 9229 4573 9263 4607
rect 13001 4573 13035 4607
rect 15301 4573 15335 4607
rect 17509 4573 17543 4607
rect 19901 4573 19935 4607
rect 27997 4573 28031 4607
rect 28825 4573 28859 4607
rect 4905 4505 4939 4539
rect 10609 4505 10643 4539
rect 11621 4505 11655 4539
rect 18245 4505 18279 4539
rect 949 4437 983 4471
rect 1501 4437 1535 4471
rect 3433 4437 3467 4471
rect 11437 4437 11471 4471
rect 11897 4437 11931 4471
rect 12357 4437 12391 4471
rect 12541 4437 12575 4471
rect 13921 4437 13955 4471
rect 15025 4437 15059 4471
rect 15669 4437 15703 4471
rect 16589 4437 16623 4471
rect 16957 4437 16991 4471
rect 18337 4437 18371 4471
rect 19257 4437 19291 4471
rect 19349 4437 19383 4471
rect 20637 4437 20671 4471
rect 20729 4437 20763 4471
rect 20821 4437 20855 4471
rect 26617 4437 26651 4471
rect 2053 4233 2087 4267
rect 11713 4233 11747 4267
rect 14473 4233 14507 4267
rect 15108 4233 15142 4267
rect 15301 4233 15335 4267
rect 15577 4233 15611 4267
rect 16773 4233 16807 4267
rect 17785 4233 17819 4267
rect 18061 4233 18095 4267
rect 18245 4233 18279 4267
rect 20085 4233 20119 4267
rect 21557 4233 21591 4267
rect 21741 4233 21775 4267
rect 22753 4233 22787 4267
rect 23029 4233 23063 4267
rect 23213 4233 23247 4267
rect 24041 4233 24075 4267
rect 24317 4233 24351 4267
rect 24501 4233 24535 4267
rect 24777 4233 24811 4267
rect 30757 4233 30791 4267
rect 1777 4165 1811 4199
rect 10977 4165 11011 4199
rect 14657 4165 14691 4199
rect 15761 4165 15795 4199
rect 17325 4165 17359 4199
rect 19901 4165 19935 4199
rect 23857 4165 23891 4199
rect 29377 4165 29411 4199
rect 30205 4165 30239 4199
rect 17417 4097 17451 4131
rect 1501 4029 1535 4063
rect 1593 4029 1627 4063
rect 1869 4029 1903 4063
rect 1961 4029 1995 4063
rect 2237 4029 2271 4063
rect 2697 4029 2731 4063
rect 3617 4029 3651 4063
rect 5641 4029 5675 4063
rect 9597 4029 9631 4063
rect 9853 4029 9887 4063
rect 17049 4029 17083 4063
rect 17233 4029 17267 4063
rect 17509 4029 17543 4063
rect 20361 4029 20395 4063
rect 26157 4029 26191 4063
rect 27997 4029 28031 4063
rect 28457 4029 28491 4063
rect 29193 4029 29227 4063
rect 29285 4029 29319 4063
rect 29561 4029 29595 4063
rect 29837 4029 29871 4063
rect 30113 4029 30147 4063
rect 30389 4029 30423 4063
rect 30665 4029 30699 4063
rect 22707 3995 22741 4029
rect 3862 3961 3896 3995
rect 5886 3961 5920 3995
rect 11529 3961 11563 3995
rect 11745 3961 11779 3995
rect 14289 3961 14323 3995
rect 14505 3961 14539 3995
rect 14933 3961 14967 3995
rect 15133 3961 15167 3995
rect 15393 3961 15427 3995
rect 16957 3961 16991 3995
rect 17877 3961 17911 3995
rect 20064 3961 20098 3995
rect 20269 3961 20303 3995
rect 21925 3961 21959 3995
rect 22937 3961 22971 3995
rect 23397 3961 23431 3995
rect 24225 3961 24259 3995
rect 24685 3961 24719 3995
rect 25912 3961 25946 3995
rect 27730 3961 27764 3995
rect 28549 3961 28583 3995
rect 29101 3961 29135 3995
rect 2329 3893 2363 3927
rect 2605 3893 2639 3927
rect 4997 3893 5031 3927
rect 7021 3893 7055 3927
rect 11897 3893 11931 3927
rect 15593 3893 15627 3927
rect 16589 3893 16623 3927
rect 16757 3893 16791 3927
rect 18077 3893 18111 3927
rect 20545 3893 20579 3927
rect 21725 3893 21759 3927
rect 22569 3893 22603 3927
rect 23187 3893 23221 3927
rect 24015 3893 24049 3927
rect 24485 3893 24519 3927
rect 26617 3893 26651 3927
rect 29653 3893 29687 3927
rect 29929 3893 29963 3927
rect 30481 3893 30515 3927
rect 1961 3689 1995 3723
rect 2513 3689 2547 3723
rect 4169 3689 4203 3723
rect 12751 3689 12785 3723
rect 13829 3689 13863 3723
rect 14825 3689 14859 3723
rect 15117 3689 15151 3723
rect 15285 3689 15319 3723
rect 16513 3689 16547 3723
rect 16681 3689 16715 3723
rect 17249 3689 17283 3723
rect 17417 3689 17451 3723
rect 18889 3689 18923 3723
rect 19349 3689 19383 3723
rect 20269 3689 20303 3723
rect 21281 3689 21315 3723
rect 21741 3689 21775 3723
rect 21909 3689 21943 3723
rect 23505 3689 23539 3723
rect 23673 3689 23707 3723
rect 24593 3689 24627 3723
rect 27261 3689 27295 3723
rect 27537 3689 27571 3723
rect 27813 3689 27847 3723
rect 28733 3689 28767 3723
rect 29009 3689 29043 3723
rect 29377 3689 29411 3723
rect 2237 3621 2271 3655
rect 12541 3621 12575 3655
rect 13027 3621 13061 3655
rect 13461 3621 13495 3655
rect 13677 3621 13711 3655
rect 14197 3621 14231 3655
rect 14413 3621 14447 3655
rect 15025 3621 15059 3655
rect 15485 3621 15519 3655
rect 16313 3621 16347 3655
rect 17049 3621 17083 3655
rect 19041 3621 19075 3655
rect 19257 3621 19291 3655
rect 19512 3621 19546 3655
rect 19717 3621 19751 3655
rect 19901 3621 19935 3655
rect 20101 3621 20135 3655
rect 21449 3621 21483 3655
rect 21649 3621 21683 3655
rect 22109 3621 22143 3655
rect 23305 3621 23339 3655
rect 25706 3621 25740 3655
rect 29806 3621 29840 3655
rect 13231 3587 13265 3621
rect 1317 3553 1351 3587
rect 1409 3553 1443 3587
rect 1593 3553 1627 3587
rect 2053 3553 2087 3587
rect 2329 3553 2363 3587
rect 2421 3553 2455 3587
rect 3056 3553 3090 3587
rect 6561 3553 6595 3587
rect 6828 3553 6862 3587
rect 8289 3553 8323 3587
rect 26801 3553 26835 3587
rect 26893 3553 26927 3587
rect 27169 3553 27203 3587
rect 27445 3553 27479 3587
rect 27721 3553 27755 3587
rect 28365 3553 28399 3587
rect 28457 3553 28491 3587
rect 28825 3553 28859 3587
rect 29101 3553 29135 3587
rect 29285 3553 29319 3587
rect 2789 3485 2823 3519
rect 8033 3485 8067 3519
rect 25973 3485 26007 3519
rect 29561 3485 29595 3519
rect 9413 3417 9447 3451
rect 12909 3417 12943 3451
rect 13369 3417 13403 3451
rect 14565 3417 14599 3451
rect 14657 3417 14691 3451
rect 1685 3349 1719 3383
rect 7941 3349 7975 3383
rect 12725 3349 12759 3383
rect 13185 3349 13219 3383
rect 13645 3349 13679 3383
rect 14381 3349 14415 3383
rect 14841 3349 14875 3383
rect 15301 3349 15335 3383
rect 16497 3349 16531 3383
rect 17233 3349 17267 3383
rect 19073 3349 19107 3383
rect 19533 3349 19567 3383
rect 20085 3349 20119 3383
rect 21465 3349 21499 3383
rect 21925 3349 21959 3383
rect 23489 3349 23523 3383
rect 30941 3349 30975 3383
rect 2973 3145 3007 3179
rect 8217 3145 8251 3179
rect 12633 3145 12667 3179
rect 13001 3145 13035 3179
rect 13185 3145 13219 3179
rect 14933 3145 14967 3179
rect 17141 3145 17175 3179
rect 18705 3145 18739 3179
rect 21557 3145 21591 3179
rect 23305 3145 23339 3179
rect 23857 3145 23891 3179
rect 29101 3145 29135 3179
rect 29929 3145 29963 3179
rect 10977 3077 11011 3111
rect 26617 3077 26651 3111
rect 27169 3077 27203 3111
rect 27445 3077 27479 3111
rect 1869 2943 1903 2977
rect 2145 2941 2179 2975
rect 2329 2941 2363 2975
rect 2789 2941 2823 2975
rect 2881 2941 2915 2975
rect 3893 2941 3927 2975
rect 5365 2941 5399 2975
rect 6837 2941 6871 2975
rect 9597 2941 9631 2975
rect 11253 2941 11287 2975
rect 13553 2941 13587 2975
rect 15761 2941 15795 2975
rect 20085 2941 20119 2975
rect 20177 2941 20211 2975
rect 21925 2941 21959 2975
rect 25237 2941 25271 2975
rect 25329 2941 25363 2975
rect 25605 2941 25639 2975
rect 26065 2941 26099 2975
rect 26157 2941 26191 2975
rect 26525 2941 26559 2975
rect 26801 2941 26835 2975
rect 27077 2941 27111 2975
rect 28825 2941 28859 2975
rect 29009 2941 29043 2975
rect 29837 2941 29871 2975
rect 31033 2941 31067 2975
rect 1777 2873 1811 2907
rect 2053 2873 2087 2907
rect 4138 2873 4172 2907
rect 5610 2873 5644 2907
rect 7082 2873 7116 2907
rect 9864 2873 9898 2907
rect 11498 2873 11532 2907
rect 12817 2873 12851 2907
rect 13033 2873 13067 2907
rect 13820 2873 13854 2907
rect 16028 2873 16062 2907
rect 19818 2873 19852 2907
rect 20422 2873 20456 2907
rect 22192 2873 22226 2907
rect 24970 2873 25004 2907
rect 26249 2873 26283 2907
rect 26893 2873 26927 2907
rect 28580 2873 28614 2907
rect 2421 2805 2455 2839
rect 2697 2805 2731 2839
rect 5273 2805 5307 2839
rect 6745 2805 6779 2839
rect 25421 2805 25455 2839
rect 25697 2805 25731 2839
rect 25973 2805 26007 2839
rect 2421 2601 2455 2635
rect 10793 2601 10827 2635
rect 13001 2601 13035 2635
rect 14473 2601 14507 2635
rect 15945 2601 15979 2635
rect 17969 2601 18003 2635
rect 19533 2601 19567 2635
rect 20269 2601 20303 2635
rect 24041 2601 24075 2635
rect 26617 2601 26651 2635
rect 27261 2601 27295 2635
rect 27537 2601 27571 2635
rect 26157 2533 26191 2567
rect 26893 2533 26927 2567
rect 2513 2465 2547 2499
rect 2605 2465 2639 2499
rect 3065 2465 3099 2499
rect 3157 2465 3191 2499
rect 3433 2465 3467 2499
rect 3709 2465 3743 2499
rect 3985 2465 4019 2499
rect 4445 2465 4479 2499
rect 4629 2465 4663 2499
rect 5273 2465 5307 2499
rect 7205 2465 7239 2499
rect 7941 2465 7975 2499
rect 8208 2465 8242 2499
rect 9413 2465 9447 2499
rect 9680 2465 9714 2499
rect 11621 2465 11655 2499
rect 11877 2465 11911 2499
rect 13093 2465 13127 2499
rect 13349 2465 13383 2499
rect 14565 2465 14599 2499
rect 14821 2465 14855 2499
rect 16856 2465 16890 2499
rect 18153 2465 18187 2499
rect 18409 2465 18443 2499
rect 20177 2465 20211 2499
rect 22854 2465 22888 2499
rect 23121 2465 23155 2499
rect 24133 2465 24167 2499
rect 24225 2465 24259 2499
rect 25421 2465 25455 2499
rect 25513 2465 25547 2499
rect 25973 2465 26007 2499
rect 26065 2465 26099 2499
rect 26709 2465 26743 2499
rect 26801 2465 26835 2499
rect 27353 2465 27387 2499
rect 27445 2465 27479 2499
rect 3801 2397 3835 2431
rect 4077 2397 4111 2431
rect 16589 2397 16623 2431
rect 2697 2329 2731 2363
rect 2973 2329 3007 2363
rect 3249 2329 3283 2363
rect 25329 2329 25363 2363
rect 25881 2329 25915 2363
rect 3525 2261 3559 2295
rect 4353 2261 4387 2295
rect 4721 2261 4755 2295
rect 5181 2261 5215 2295
rect 7297 2261 7331 2295
rect 9321 2261 9355 2295
rect 21741 2261 21775 2295
rect 24317 2261 24351 2295
rect 25605 2261 25639 2295
rect 31033 2261 31067 2295
rect 2697 2057 2731 2091
rect 3341 2057 3375 2091
rect 6377 2057 6411 2091
rect 7205 2057 7239 2091
rect 7481 2057 7515 2091
rect 8125 2057 8159 2091
rect 12173 2057 12207 2091
rect 16129 2057 16163 2091
rect 17141 2057 17175 2091
rect 18061 2057 18095 2091
rect 19809 2057 19843 2091
rect 20085 2057 20119 2091
rect 21741 2057 21775 2091
rect 23949 2057 23983 2091
rect 24225 2057 24259 2091
rect 24501 2057 24535 2091
rect 25145 2057 25179 2091
rect 4997 1989 5031 2023
rect 6101 1921 6135 1955
rect 10793 1921 10827 1955
rect 15301 1921 15335 1955
rect 15853 1921 15887 1955
rect 20361 1921 20395 1955
rect 23581 1921 23615 1955
rect 2789 1853 2823 1887
rect 3249 1853 3283 1887
rect 4629 1853 4663 1887
rect 4721 1853 4755 1887
rect 5065 1853 5099 1887
rect 5173 1853 5207 1887
rect 5457 1853 5491 1887
rect 5917 1853 5951 1887
rect 6193 1853 6227 1887
rect 6285 1853 6319 1887
rect 6561 1853 6595 1887
rect 6837 1853 6871 1887
rect 7297 1853 7331 1887
rect 7389 1853 7423 1887
rect 7757 1853 7791 1887
rect 8033 1853 8067 1887
rect 8401 1853 8435 1887
rect 9505 1853 9539 1887
rect 9597 1853 9631 1887
rect 12449 1853 12483 1887
rect 12541 1853 12575 1887
rect 14565 1853 14599 1887
rect 15209 1853 15243 1887
rect 15485 1855 15519 1889
rect 15577 1853 15611 1887
rect 15761 1853 15795 1887
rect 16037 1853 16071 1887
rect 16313 1853 16347 1887
rect 16957 1853 16991 1887
rect 17057 1853 17091 1887
rect 17325 1853 17359 1887
rect 17417 1853 17451 1887
rect 17969 1853 18003 1887
rect 18245 1853 18279 1887
rect 19717 1853 19751 1887
rect 19993 1853 20027 1887
rect 22017 1853 22051 1887
rect 23489 1853 23523 1887
rect 23857 1853 23891 1887
rect 24317 1853 24351 1887
rect 24593 1853 24627 1887
rect 24685 1853 24719 1887
rect 26525 1853 26559 1887
rect 31033 1853 31067 1887
rect 5549 1785 5583 1819
rect 5825 1785 5859 1819
rect 6653 1785 6687 1819
rect 6929 1785 6963 1819
rect 7849 1785 7883 1819
rect 8493 1785 8527 1819
rect 11038 1785 11072 1819
rect 20606 1785 20640 1819
rect 24777 1785 24811 1819
rect 26258 1785 26292 1819
rect 5273 1717 5307 1751
rect 9413 1717 9447 1751
rect 9689 1717 9723 1751
rect 12357 1717 12391 1751
rect 12633 1717 12667 1751
rect 14473 1717 14507 1751
rect 16405 1717 16439 1751
rect 16865 1717 16899 1751
rect 18337 1717 18371 1751
rect 21925 1717 21959 1751
rect 7389 1513 7423 1547
rect 8217 1513 8251 1547
rect 9873 1513 9907 1547
rect 10149 1513 10183 1547
rect 12633 1513 12667 1547
rect 13093 1513 13127 1547
rect 13921 1513 13955 1547
rect 15853 1513 15887 1547
rect 16405 1513 16439 1547
rect 17325 1513 17359 1547
rect 17693 1513 17727 1547
rect 17969 1513 18003 1547
rect 18521 1513 18555 1547
rect 18797 1513 18831 1547
rect 19073 1513 19107 1547
rect 19349 1513 19383 1547
rect 20177 1513 20211 1547
rect 20729 1513 20763 1547
rect 22477 1513 22511 1547
rect 22753 1513 22787 1547
rect 23489 1513 23523 1547
rect 23765 1513 23799 1547
rect 25421 1513 25455 1547
rect 10425 1445 10459 1479
rect 10701 1445 10735 1479
rect 11069 1445 11103 1479
rect 13369 1445 13403 1479
rect 7481 1377 7515 1411
rect 7573 1377 7607 1411
rect 7849 1377 7883 1411
rect 7941 1377 7975 1411
rect 8125 1377 8159 1411
rect 8401 1377 8435 1411
rect 8677 1377 8711 1411
rect 9045 1377 9079 1411
rect 9137 1377 9171 1411
rect 9229 1377 9263 1411
rect 9689 1377 9723 1411
rect 9781 1377 9815 1411
rect 10241 1377 10275 1411
rect 10517 1377 10551 1411
rect 10793 1377 10827 1411
rect 10977 1377 11011 1411
rect 11253 1377 11287 1411
rect 11520 1377 11554 1411
rect 12725 1377 12759 1411
rect 13001 1377 13035 1411
rect 13277 1377 13311 1411
rect 13553 1377 13587 1411
rect 13645 1377 13679 1411
rect 14013 1377 14047 1411
rect 14289 1377 14323 1411
rect 14381 1377 14415 1411
rect 14657 1377 14691 1411
rect 14749 1377 14783 1411
rect 15301 1377 15335 1411
rect 15485 1377 15519 1411
rect 15577 1377 15611 1411
rect 15945 1377 15979 1411
rect 16221 1377 16255 1411
rect 17141 1377 17175 1411
rect 17233 1377 17267 1411
rect 17509 1377 17543 1411
rect 18061 1377 18095 1411
rect 18245 1377 18279 1411
rect 18705 1377 18739 1411
rect 19165 1377 19199 1411
rect 19257 1377 19291 1411
rect 19533 1377 19567 1411
rect 19809 1377 19843 1411
rect 20269 1377 20303 1411
rect 20361 1377 20395 1411
rect 20453 1377 20487 1411
rect 20637 1377 20671 1411
rect 20913 1377 20947 1411
rect 21465 1377 21499 1411
rect 21557 1377 21591 1411
rect 21833 1377 21867 1411
rect 22109 1377 22143 1411
rect 22385 1377 22419 1411
rect 22661 1377 22695 1411
rect 22937 1377 22971 1411
rect 23029 1377 23063 1411
rect 23581 1377 23615 1411
rect 24878 1377 24912 1411
rect 25145 1377 25179 1411
rect 25329 1377 25363 1411
rect 7665 1309 7699 1343
rect 8493 1309 8527 1343
rect 12817 1309 12851 1343
rect 21649 1309 21683 1343
rect 21925 1309 21959 1343
rect 8769 1241 8803 1275
rect 9321 1241 9355 1275
rect 9597 1241 9631 1275
rect 14473 1241 14507 1275
rect 15209 1241 15243 1275
rect 17049 1241 17083 1275
rect 19625 1241 19659 1275
rect 19901 1241 19935 1275
rect 14197 1173 14231 1207
rect 21005 1173 21039 1207
rect 21373 1173 21407 1207
rect 22201 1173 22235 1207
rect 8125 969 8159 1003
rect 8493 969 8527 1003
rect 9413 969 9447 1003
rect 9873 969 9907 1003
rect 12265 969 12299 1003
rect 13093 969 13127 1003
rect 14473 969 14507 1003
rect 15761 969 15795 1003
rect 17509 969 17543 1003
rect 20085 969 20119 1003
rect 20729 969 20763 1003
rect 21925 969 21959 1003
rect 23949 969 23983 1003
rect 24225 969 24259 1003
rect 24501 969 24535 1003
rect 14749 901 14783 935
rect 23489 901 23523 935
rect 18705 833 18739 867
rect 21373 833 21407 867
rect 21649 833 21683 867
rect 22109 833 22143 867
rect 8033 765 8067 799
rect 8585 765 8619 799
rect 9505 765 9539 799
rect 9965 765 9999 799
rect 11897 765 11931 799
rect 11989 765 12023 799
rect 12357 765 12391 799
rect 12633 765 12667 799
rect 13185 765 13219 799
rect 14565 765 14599 799
rect 14657 765 14691 799
rect 16129 765 16163 799
rect 17601 765 17635 799
rect 17877 765 17911 799
rect 18972 765 19006 799
rect 20821 765 20855 799
rect 21281 765 21315 799
rect 21741 765 21775 799
rect 21833 765 21867 799
rect 22376 765 22410 799
rect 24041 765 24075 799
rect 24133 765 24167 799
rect 24593 765 24627 799
rect 31033 765 31067 799
rect 12725 697 12759 731
rect 15669 697 15703 731
rect 16374 697 16408 731
<< metal1 >>
rect 552 19066 31531 19088
rect 552 19014 8102 19066
rect 8154 19014 8166 19066
rect 8218 19014 8230 19066
rect 8282 19014 8294 19066
rect 8346 19014 8358 19066
rect 8410 19014 15807 19066
rect 15859 19014 15871 19066
rect 15923 19014 15935 19066
rect 15987 19014 15999 19066
rect 16051 19014 16063 19066
rect 16115 19014 23512 19066
rect 23564 19014 23576 19066
rect 23628 19014 23640 19066
rect 23692 19014 23704 19066
rect 23756 19014 23768 19066
rect 23820 19014 31217 19066
rect 31269 19014 31281 19066
rect 31333 19014 31345 19066
rect 31397 19014 31409 19066
rect 31461 19014 31473 19066
rect 31525 19014 31531 19066
rect 552 18992 31531 19014
rect 10689 18887 10747 18893
rect 10689 18884 10701 18887
rect 10336 18856 10701 18884
rect 750 18776 756 18828
rect 808 18816 814 18828
rect 1397 18819 1455 18825
rect 1397 18816 1409 18819
rect 808 18788 1409 18816
rect 808 18776 814 18788
rect 1397 18785 1409 18788
rect 1443 18785 1455 18819
rect 1397 18779 1455 18785
rect 6454 18776 6460 18828
rect 6512 18816 6518 18828
rect 6549 18819 6607 18825
rect 6549 18816 6561 18819
rect 6512 18788 6561 18816
rect 6512 18776 6518 18788
rect 6549 18785 6561 18788
rect 6595 18785 6607 18819
rect 6549 18779 6607 18785
rect 7098 18776 7104 18828
rect 7156 18816 7162 18828
rect 7193 18819 7251 18825
rect 7193 18816 7205 18819
rect 7156 18788 7205 18816
rect 7156 18776 7162 18788
rect 7193 18785 7205 18788
rect 7239 18785 7251 18819
rect 7193 18779 7251 18785
rect 7742 18776 7748 18828
rect 7800 18816 7806 18828
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7800 18788 7849 18816
rect 7800 18776 7806 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 8573 18819 8631 18825
rect 8573 18816 8585 18819
rect 7837 18779 7895 18785
rect 7944 18788 8585 18816
rect 1118 18708 1124 18760
rect 1176 18708 1182 18760
rect 7944 18624 7972 18788
rect 8573 18785 8585 18788
rect 8619 18785 8631 18819
rect 8573 18779 8631 18785
rect 8588 18748 8616 18779
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 9548 18788 9689 18816
rect 9548 18776 9554 18788
rect 9677 18785 9689 18788
rect 9723 18816 9735 18819
rect 9861 18819 9919 18825
rect 9861 18816 9873 18819
rect 9723 18788 9873 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 9861 18785 9873 18788
rect 9907 18785 9919 18819
rect 9861 18779 9919 18785
rect 9953 18819 10011 18825
rect 9953 18785 9965 18819
rect 9999 18785 10011 18819
rect 9953 18779 10011 18785
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 8588 18720 9597 18748
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 9968 18748 9996 18779
rect 10134 18776 10140 18828
rect 10192 18816 10198 18828
rect 10229 18819 10287 18825
rect 10229 18816 10241 18819
rect 10192 18788 10241 18816
rect 10192 18776 10198 18788
rect 10229 18785 10241 18788
rect 10275 18785 10287 18819
rect 10229 18779 10287 18785
rect 10336 18748 10364 18856
rect 10689 18853 10701 18856
rect 10735 18853 10747 18887
rect 10689 18847 10747 18853
rect 20824 18856 22416 18884
rect 10502 18776 10508 18828
rect 10560 18776 10566 18828
rect 10597 18819 10655 18825
rect 10597 18785 10609 18819
rect 10643 18785 10655 18819
rect 10597 18779 10655 18785
rect 10612 18748 10640 18779
rect 9968 18720 10364 18748
rect 10428 18720 10640 18748
rect 10704 18748 10732 18847
rect 20824 18828 20852 18856
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 11422 18825 11428 18828
rect 11149 18819 11207 18825
rect 11149 18816 11161 18819
rect 10836 18788 11161 18816
rect 10836 18776 10842 18788
rect 11149 18785 11161 18788
rect 11195 18785 11207 18819
rect 11405 18819 11428 18825
rect 11405 18816 11417 18819
rect 11149 18779 11207 18785
rect 11256 18788 11417 18816
rect 11256 18748 11284 18788
rect 11405 18785 11417 18788
rect 11405 18779 11428 18785
rect 11422 18776 11428 18779
rect 11480 18776 11486 18828
rect 13900 18819 13958 18825
rect 13900 18785 13912 18819
rect 13946 18816 13958 18819
rect 14182 18816 14188 18828
rect 13946 18788 14188 18816
rect 13946 18785 13958 18788
rect 13900 18779 13958 18785
rect 14182 18776 14188 18788
rect 14240 18776 14246 18828
rect 16117 18819 16175 18825
rect 16117 18785 16129 18819
rect 16163 18816 16175 18819
rect 16206 18816 16212 18828
rect 16163 18788 16212 18816
rect 16163 18785 16175 18788
rect 16117 18779 16175 18785
rect 16206 18776 16212 18788
rect 16264 18776 16270 18828
rect 16384 18819 16442 18825
rect 16384 18785 16396 18819
rect 16430 18816 16442 18819
rect 16942 18816 16948 18828
rect 16430 18788 16948 18816
rect 16430 18785 16442 18788
rect 16384 18779 16442 18785
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 19236 18819 19294 18825
rect 19236 18785 19248 18819
rect 19282 18816 19294 18819
rect 20806 18816 20812 18828
rect 19282 18788 20812 18816
rect 19282 18785 19294 18788
rect 19236 18779 19294 18785
rect 20806 18776 20812 18788
rect 20864 18776 20870 18828
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18816 20959 18819
rect 20990 18816 20996 18828
rect 20947 18788 20996 18816
rect 20947 18785 20959 18788
rect 20901 18779 20959 18785
rect 20990 18776 20996 18788
rect 21048 18816 21054 18828
rect 21269 18819 21327 18825
rect 21269 18816 21281 18819
rect 21048 18788 21281 18816
rect 21048 18776 21054 18788
rect 21269 18785 21281 18788
rect 21315 18785 21327 18819
rect 21269 18779 21327 18785
rect 22005 18819 22063 18825
rect 22005 18785 22017 18819
rect 22051 18816 22063 18819
rect 22281 18819 22339 18825
rect 22281 18816 22293 18819
rect 22051 18788 22293 18816
rect 22051 18785 22063 18788
rect 22005 18779 22063 18785
rect 10704 18720 11284 18748
rect 9968 18680 9996 18720
rect 8956 18652 9996 18680
rect 8956 18624 8984 18652
rect 842 18572 848 18624
rect 900 18572 906 18624
rect 7926 18572 7932 18624
rect 7984 18572 7990 18624
rect 8478 18572 8484 18624
rect 8536 18572 8542 18624
rect 8938 18572 8944 18624
rect 8996 18572 9002 18624
rect 9858 18572 9864 18624
rect 9916 18612 9922 18624
rect 10428 18621 10456 18720
rect 13630 18708 13636 18760
rect 13688 18708 13694 18760
rect 17862 18708 17868 18760
rect 17920 18748 17926 18760
rect 18969 18751 19027 18757
rect 18969 18748 18981 18751
rect 17920 18720 18981 18748
rect 17920 18708 17926 18720
rect 18969 18717 18981 18720
rect 19015 18717 19027 18751
rect 18969 18711 19027 18717
rect 21361 18683 21419 18689
rect 21361 18680 21373 18683
rect 19996 18652 21373 18680
rect 19996 18624 20024 18652
rect 21361 18649 21373 18652
rect 21407 18680 21419 18683
rect 21913 18683 21971 18689
rect 21913 18680 21925 18683
rect 21407 18652 21925 18680
rect 21407 18649 21419 18652
rect 21361 18643 21419 18649
rect 21913 18649 21925 18652
rect 21959 18649 21971 18683
rect 21913 18643 21971 18649
rect 10137 18615 10195 18621
rect 10137 18612 10149 18615
rect 9916 18584 10149 18612
rect 9916 18572 9922 18584
rect 10137 18581 10149 18584
rect 10183 18612 10195 18615
rect 10413 18615 10471 18621
rect 10413 18612 10425 18615
rect 10183 18584 10425 18612
rect 10183 18581 10195 18584
rect 10137 18575 10195 18581
rect 10413 18581 10425 18584
rect 10459 18581 10471 18615
rect 10413 18575 10471 18581
rect 12526 18572 12532 18624
rect 12584 18572 12590 18624
rect 15010 18572 15016 18624
rect 15068 18572 15074 18624
rect 17034 18572 17040 18624
rect 17092 18612 17098 18624
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 17092 18584 17509 18612
rect 17092 18572 17098 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 19978 18572 19984 18624
rect 20036 18572 20042 18624
rect 20349 18615 20407 18621
rect 20349 18581 20361 18615
rect 20395 18612 20407 18615
rect 20714 18612 20720 18624
rect 20395 18584 20720 18612
rect 20395 18581 20407 18584
rect 20349 18575 20407 18581
rect 20714 18572 20720 18584
rect 20772 18572 20778 18624
rect 22112 18612 22140 18788
rect 22281 18785 22293 18788
rect 22327 18785 22339 18819
rect 22281 18779 22339 18785
rect 22189 18683 22247 18689
rect 22189 18649 22201 18683
rect 22235 18680 22247 18683
rect 22388 18680 22416 18856
rect 22833 18819 22891 18825
rect 22833 18785 22845 18819
rect 22879 18816 22891 18819
rect 23198 18816 23204 18828
rect 22879 18788 23204 18816
rect 22879 18785 22891 18788
rect 22833 18779 22891 18785
rect 23198 18776 23204 18788
rect 23256 18816 23262 18828
rect 24958 18819 25016 18825
rect 24958 18816 24970 18819
rect 23256 18788 24970 18816
rect 23256 18776 23262 18788
rect 24958 18785 24970 18788
rect 25004 18785 25016 18819
rect 24958 18779 25016 18785
rect 27706 18776 27712 18828
rect 27764 18816 27770 18828
rect 27801 18819 27859 18825
rect 27801 18816 27813 18819
rect 27764 18788 27813 18816
rect 27764 18776 27770 18788
rect 27801 18785 27813 18788
rect 27847 18785 27859 18819
rect 27801 18779 27859 18785
rect 28350 18776 28356 18828
rect 28408 18816 28414 18828
rect 28445 18819 28503 18825
rect 28445 18816 28457 18819
rect 28408 18788 28457 18816
rect 28408 18776 28414 18788
rect 28445 18785 28457 18788
rect 28491 18785 28503 18819
rect 28445 18779 28503 18785
rect 30745 18819 30803 18825
rect 30745 18785 30757 18819
rect 30791 18816 30803 18819
rect 31662 18816 31668 18828
rect 30791 18788 31668 18816
rect 30791 18785 30803 18788
rect 30745 18779 30803 18785
rect 31662 18776 31668 18788
rect 31720 18776 31726 18828
rect 25222 18708 25228 18760
rect 25280 18708 25286 18760
rect 22235 18652 23060 18680
rect 22235 18649 22247 18652
rect 22189 18643 22247 18649
rect 23032 18624 23060 18652
rect 22278 18612 22284 18624
rect 22112 18584 22284 18612
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 22738 18572 22744 18624
rect 22796 18572 22802 18624
rect 23014 18572 23020 18624
rect 23072 18572 23078 18624
rect 23845 18615 23903 18621
rect 23845 18581 23857 18615
rect 23891 18612 23903 18615
rect 24026 18612 24032 18624
rect 23891 18584 24032 18612
rect 23891 18581 23903 18584
rect 23845 18575 23903 18581
rect 24026 18572 24032 18584
rect 24084 18572 24090 18624
rect 31018 18572 31024 18624
rect 31076 18572 31082 18624
rect 552 18522 31372 18544
rect 552 18470 4250 18522
rect 4302 18470 4314 18522
rect 4366 18470 4378 18522
rect 4430 18470 4442 18522
rect 4494 18470 4506 18522
rect 4558 18470 11955 18522
rect 12007 18470 12019 18522
rect 12071 18470 12083 18522
rect 12135 18470 12147 18522
rect 12199 18470 12211 18522
rect 12263 18470 19660 18522
rect 19712 18470 19724 18522
rect 19776 18470 19788 18522
rect 19840 18470 19852 18522
rect 19904 18470 19916 18522
rect 19968 18470 27365 18522
rect 27417 18470 27429 18522
rect 27481 18470 27493 18522
rect 27545 18470 27557 18522
rect 27609 18470 27621 18522
rect 27673 18470 31372 18522
rect 552 18448 31372 18470
rect 9490 18368 9496 18420
rect 9548 18368 9554 18420
rect 10134 18408 10140 18420
rect 9600 18380 10140 18408
rect 8481 18343 8539 18349
rect 8481 18309 8493 18343
rect 8527 18340 8539 18343
rect 8570 18340 8576 18352
rect 8527 18312 8576 18340
rect 8527 18309 8539 18312
rect 8481 18303 8539 18309
rect 8570 18300 8576 18312
rect 8628 18300 8634 18352
rect 7009 18275 7067 18281
rect 7009 18241 7021 18275
rect 7055 18272 7067 18275
rect 7374 18272 7380 18284
rect 7055 18244 7380 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 7561 18275 7619 18281
rect 7561 18241 7573 18275
rect 7607 18272 7619 18275
rect 7742 18272 7748 18284
rect 7607 18244 7748 18272
rect 7607 18241 7619 18244
rect 7561 18235 7619 18241
rect 7742 18232 7748 18244
rect 7800 18272 7806 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7800 18244 7849 18272
rect 7800 18232 7806 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 842 18164 848 18216
rect 900 18164 906 18216
rect 7101 18207 7159 18213
rect 7101 18173 7113 18207
rect 7147 18173 7159 18207
rect 7101 18167 7159 18173
rect 7469 18207 7527 18213
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 7515 18176 7880 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 7116 18080 7144 18167
rect 7098 18028 7104 18080
rect 7156 18028 7162 18080
rect 7852 18068 7880 18176
rect 7926 18164 7932 18216
rect 7984 18164 7990 18216
rect 8205 18207 8263 18213
rect 8205 18173 8217 18207
rect 8251 18204 8263 18207
rect 8478 18204 8484 18216
rect 8251 18176 8484 18204
rect 8251 18173 8263 18176
rect 8205 18167 8263 18173
rect 8478 18164 8484 18176
rect 8536 18204 8542 18216
rect 8573 18207 8631 18213
rect 8573 18204 8585 18207
rect 8536 18176 8585 18204
rect 8536 18164 8542 18176
rect 8573 18173 8585 18176
rect 8619 18204 8631 18207
rect 8849 18207 8907 18213
rect 8849 18204 8861 18207
rect 8619 18176 8861 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 8849 18173 8861 18176
rect 8895 18173 8907 18207
rect 8849 18167 8907 18173
rect 8938 18164 8944 18216
rect 8996 18164 9002 18216
rect 9309 18207 9367 18213
rect 9309 18173 9321 18207
rect 9355 18204 9367 18207
rect 9508 18204 9536 18368
rect 9600 18213 9628 18380
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 10594 18368 10600 18420
rect 10652 18408 10658 18420
rect 12897 18411 12955 18417
rect 12897 18408 12909 18411
rect 10652 18380 12909 18408
rect 10652 18368 10658 18380
rect 11422 18300 11428 18352
rect 11480 18340 11486 18352
rect 11609 18343 11667 18349
rect 11609 18340 11621 18343
rect 11480 18312 11621 18340
rect 11480 18300 11486 18312
rect 11609 18309 11621 18312
rect 11655 18309 11667 18343
rect 11609 18303 11667 18309
rect 9766 18232 9772 18284
rect 9824 18272 9830 18284
rect 9953 18275 10011 18281
rect 9953 18272 9965 18275
rect 9824 18244 9965 18272
rect 9824 18232 9830 18244
rect 9953 18241 9965 18244
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 9355 18176 9536 18204
rect 9585 18207 9643 18213
rect 9355 18173 9367 18176
rect 9309 18167 9367 18173
rect 9585 18173 9597 18207
rect 9631 18173 9643 18207
rect 9585 18167 9643 18173
rect 9858 18164 9864 18216
rect 9916 18164 9922 18216
rect 11992 18213 12020 18380
rect 12897 18377 12909 18380
rect 12943 18408 12955 18411
rect 14182 18408 14188 18420
rect 12943 18380 14188 18408
rect 12943 18377 12955 18380
rect 12897 18371 12955 18377
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 20806 18368 20812 18420
rect 20864 18368 20870 18420
rect 20990 18368 20996 18420
rect 21048 18368 21054 18420
rect 22738 18368 22744 18420
rect 22796 18368 22802 18420
rect 23014 18368 23020 18420
rect 23072 18368 23078 18420
rect 13909 18343 13967 18349
rect 13909 18340 13921 18343
rect 12452 18312 13921 18340
rect 11701 18207 11759 18213
rect 11701 18173 11713 18207
rect 11747 18204 11759 18207
rect 11885 18207 11943 18213
rect 11885 18204 11897 18207
rect 11747 18176 11897 18204
rect 11747 18173 11759 18176
rect 11701 18167 11759 18173
rect 11885 18173 11897 18176
rect 11931 18173 11943 18207
rect 11885 18167 11943 18173
rect 11977 18207 12035 18213
rect 11977 18173 11989 18207
rect 12023 18173 12035 18207
rect 11977 18167 12035 18173
rect 7944 18136 7972 18164
rect 9769 18139 9827 18145
rect 9769 18136 9781 18139
rect 7944 18108 9781 18136
rect 9769 18105 9781 18108
rect 9815 18136 9827 18139
rect 10198 18139 10256 18145
rect 10198 18136 10210 18139
rect 9815 18108 10210 18136
rect 9815 18105 9827 18108
rect 9769 18099 9827 18105
rect 10198 18105 10210 18108
rect 10244 18105 10256 18139
rect 10198 18099 10256 18105
rect 10318 18096 10324 18148
rect 10376 18136 10382 18148
rect 11900 18136 11928 18167
rect 12250 18164 12256 18216
rect 12308 18164 12314 18216
rect 12345 18207 12403 18213
rect 12345 18173 12357 18207
rect 12391 18173 12403 18207
rect 12345 18167 12403 18173
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 10376 18108 11836 18136
rect 11900 18108 12173 18136
rect 10376 18096 10382 18108
rect 7926 18068 7932 18080
rect 7852 18040 7932 18068
rect 7926 18028 7932 18040
rect 7984 18068 7990 18080
rect 8113 18071 8171 18077
rect 8113 18068 8125 18071
rect 7984 18040 8125 18068
rect 7984 18028 7990 18040
rect 8113 18037 8125 18040
rect 8159 18068 8171 18071
rect 9214 18068 9220 18080
rect 8159 18040 9220 18068
rect 8159 18037 8171 18040
rect 8113 18031 8171 18037
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 11333 18071 11391 18077
rect 11333 18037 11345 18071
rect 11379 18068 11391 18071
rect 11606 18068 11612 18080
rect 11379 18040 11612 18068
rect 11379 18037 11391 18040
rect 11333 18031 11391 18037
rect 11606 18028 11612 18040
rect 11664 18028 11670 18080
rect 11808 18068 11836 18108
rect 12161 18105 12173 18108
rect 12207 18136 12219 18139
rect 12360 18136 12388 18167
rect 12207 18108 12388 18136
rect 12207 18105 12219 18108
rect 12161 18099 12219 18105
rect 12452 18077 12480 18312
rect 13909 18309 13921 18312
rect 13955 18309 13967 18343
rect 13909 18303 13967 18309
rect 13924 18272 13952 18303
rect 13998 18300 14004 18352
rect 14056 18340 14062 18352
rect 14056 18312 14596 18340
rect 14056 18300 14062 18312
rect 14568 18281 14596 18312
rect 14553 18275 14611 18281
rect 13924 18244 14228 18272
rect 12986 18164 12992 18216
rect 13044 18164 13050 18216
rect 13722 18164 13728 18216
rect 13780 18164 13786 18216
rect 13817 18207 13875 18213
rect 13817 18173 13829 18207
rect 13863 18204 13875 18207
rect 14093 18207 14151 18213
rect 14093 18204 14105 18207
rect 13863 18176 14105 18204
rect 13863 18173 13875 18176
rect 13817 18167 13875 18173
rect 14093 18173 14105 18176
rect 14139 18173 14151 18207
rect 14200 18204 14228 18244
rect 14553 18241 14565 18275
rect 14599 18241 14611 18275
rect 17129 18275 17187 18281
rect 17129 18272 17141 18275
rect 14553 18235 14611 18241
rect 16224 18244 17141 18272
rect 16224 18216 16252 18244
rect 17129 18241 17141 18244
rect 17175 18241 17187 18275
rect 19978 18272 19984 18284
rect 17129 18235 17187 18241
rect 19260 18244 19984 18272
rect 14809 18207 14867 18213
rect 14809 18204 14821 18207
rect 14200 18176 14821 18204
rect 14093 18167 14151 18173
rect 14809 18173 14821 18176
rect 14855 18173 14867 18207
rect 14809 18167 14867 18173
rect 13832 18136 13860 18167
rect 16206 18164 16212 18216
rect 16264 18164 16270 18216
rect 16761 18207 16819 18213
rect 16761 18173 16773 18207
rect 16807 18173 16819 18207
rect 16761 18167 16819 18173
rect 13648 18108 13860 18136
rect 16776 18136 16804 18167
rect 16942 18164 16948 18216
rect 17000 18204 17006 18216
rect 17037 18207 17095 18213
rect 17037 18204 17049 18207
rect 17000 18176 17049 18204
rect 17000 18164 17006 18176
rect 17037 18173 17049 18176
rect 17083 18204 17095 18207
rect 19260 18204 19288 18244
rect 19904 18213 19932 18244
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 20824 18272 20852 18368
rect 20180 18244 20852 18272
rect 20180 18213 20208 18244
rect 17083 18176 19288 18204
rect 19337 18207 19395 18213
rect 17083 18173 17095 18176
rect 17037 18167 17095 18173
rect 19337 18173 19349 18207
rect 19383 18204 19395 18207
rect 19613 18207 19671 18213
rect 19613 18204 19625 18207
rect 19383 18176 19625 18204
rect 19383 18173 19395 18176
rect 19337 18167 19395 18173
rect 19613 18173 19625 18176
rect 19659 18173 19671 18207
rect 19613 18167 19671 18173
rect 19889 18207 19947 18213
rect 19889 18173 19901 18207
rect 19935 18173 19947 18207
rect 19889 18167 19947 18173
rect 20165 18207 20223 18213
rect 20165 18173 20177 18207
rect 20211 18173 20223 18207
rect 20165 18167 20223 18173
rect 20717 18207 20775 18213
rect 20717 18173 20729 18207
rect 20763 18204 20775 18207
rect 21008 18204 21036 18368
rect 22756 18272 22784 18368
rect 22756 18244 23520 18272
rect 20763 18176 21036 18204
rect 21085 18207 21143 18213
rect 20763 18173 20775 18176
rect 20717 18167 20775 18173
rect 21085 18173 21097 18207
rect 21131 18204 21143 18207
rect 22373 18207 22431 18213
rect 22373 18204 22385 18207
rect 21131 18176 22385 18204
rect 21131 18173 21143 18176
rect 21085 18167 21143 18173
rect 17396 18139 17454 18145
rect 17396 18136 17408 18139
rect 16776 18108 17408 18136
rect 12437 18071 12495 18077
rect 12437 18068 12449 18071
rect 11808 18040 12449 18068
rect 12437 18037 12449 18040
rect 12483 18037 12495 18071
rect 12437 18031 12495 18037
rect 13354 18028 13360 18080
rect 13412 18068 13418 18080
rect 13648 18077 13676 18108
rect 17396 18105 17408 18108
rect 17442 18136 17454 18139
rect 18690 18136 18696 18148
rect 17442 18108 18696 18136
rect 17442 18105 17454 18108
rect 17396 18099 17454 18105
rect 18690 18096 18696 18108
rect 18748 18136 18754 18148
rect 19628 18136 19656 18167
rect 19797 18139 19855 18145
rect 19797 18136 19809 18139
rect 18748 18108 19564 18136
rect 19628 18108 19809 18136
rect 18748 18096 18754 18108
rect 13633 18071 13691 18077
rect 13633 18068 13645 18071
rect 13412 18040 13645 18068
rect 13412 18028 13418 18040
rect 13633 18037 13645 18040
rect 13679 18037 13691 18071
rect 13633 18031 13691 18037
rect 15933 18071 15991 18077
rect 15933 18037 15945 18071
rect 15979 18068 15991 18071
rect 16298 18068 16304 18080
rect 15979 18040 16304 18068
rect 15979 18037 15991 18040
rect 15933 18031 15991 18037
rect 16298 18028 16304 18040
rect 16356 18028 16362 18080
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 16669 18071 16727 18077
rect 16669 18068 16681 18071
rect 16632 18040 16681 18068
rect 16632 18028 16638 18040
rect 16669 18037 16681 18040
rect 16715 18068 16727 18071
rect 16942 18068 16948 18080
rect 16715 18040 16948 18068
rect 16715 18037 16727 18040
rect 16669 18031 16727 18037
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 18509 18071 18567 18077
rect 18509 18037 18521 18071
rect 18555 18068 18567 18071
rect 18782 18068 18788 18080
rect 18555 18040 18788 18068
rect 18555 18037 18567 18040
rect 18509 18031 18567 18037
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 19242 18028 19248 18080
rect 19300 18028 19306 18080
rect 19536 18077 19564 18108
rect 19797 18105 19809 18108
rect 19843 18136 19855 18139
rect 20073 18139 20131 18145
rect 20073 18136 20085 18139
rect 19843 18108 20085 18136
rect 19843 18105 19855 18108
rect 19797 18099 19855 18105
rect 20073 18105 20085 18108
rect 20119 18105 20131 18139
rect 20073 18099 20131 18105
rect 19521 18071 19579 18077
rect 19521 18037 19533 18071
rect 19567 18068 19579 18071
rect 20625 18071 20683 18077
rect 20625 18068 20637 18071
rect 19567 18040 20637 18068
rect 19567 18037 19579 18040
rect 19521 18031 19579 18037
rect 20625 18037 20637 18040
rect 20671 18037 20683 18071
rect 22112 18068 22140 18176
rect 22373 18173 22385 18176
rect 22419 18173 22431 18207
rect 22373 18167 22431 18173
rect 22830 18164 22836 18216
rect 22888 18164 22894 18216
rect 23124 18213 23152 18244
rect 23109 18207 23167 18213
rect 23109 18173 23121 18207
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 23198 18164 23204 18216
rect 23256 18204 23262 18216
rect 23492 18213 23520 18244
rect 23385 18207 23443 18213
rect 23385 18204 23397 18207
rect 23256 18176 23397 18204
rect 23256 18164 23262 18176
rect 23385 18173 23397 18176
rect 23431 18173 23443 18207
rect 23385 18167 23443 18173
rect 23477 18207 23535 18213
rect 23477 18173 23489 18207
rect 23523 18173 23535 18207
rect 23477 18167 23535 18173
rect 24029 18207 24087 18213
rect 24029 18173 24041 18207
rect 24075 18204 24087 18207
rect 24302 18204 24308 18216
rect 24075 18176 24308 18204
rect 24075 18173 24087 18176
rect 24029 18167 24087 18173
rect 22278 18096 22284 18148
rect 22336 18136 22342 18148
rect 23293 18139 23351 18145
rect 23293 18136 23305 18139
rect 22336 18108 23305 18136
rect 22336 18096 22342 18108
rect 23293 18105 23305 18108
rect 23339 18105 23351 18139
rect 23400 18136 23428 18167
rect 24302 18164 24308 18176
rect 24360 18204 24366 18216
rect 24397 18207 24455 18213
rect 24397 18204 24409 18207
rect 24360 18176 24409 18204
rect 24360 18164 24366 18176
rect 24397 18173 24409 18176
rect 24443 18173 24455 18207
rect 24397 18167 24455 18173
rect 24946 18164 24952 18216
rect 25004 18164 25010 18216
rect 24857 18139 24915 18145
rect 24857 18136 24869 18139
rect 23400 18108 24869 18136
rect 23293 18099 23351 18105
rect 22370 18068 22376 18080
rect 22112 18040 22376 18068
rect 20625 18031 20683 18037
rect 22370 18028 22376 18040
rect 22428 18068 22434 18080
rect 24320 18077 24348 18108
rect 24857 18105 24869 18108
rect 24903 18105 24915 18139
rect 24857 18099 24915 18105
rect 23569 18071 23627 18077
rect 23569 18068 23581 18071
rect 22428 18040 23581 18068
rect 22428 18028 22434 18040
rect 23569 18037 23581 18040
rect 23615 18068 23627 18071
rect 23937 18071 23995 18077
rect 23937 18068 23949 18071
rect 23615 18040 23949 18068
rect 23615 18037 23627 18040
rect 23569 18031 23627 18037
rect 23937 18037 23949 18040
rect 23983 18037 23995 18071
rect 23937 18031 23995 18037
rect 24305 18071 24363 18077
rect 24305 18037 24317 18071
rect 24351 18037 24363 18071
rect 24305 18031 24363 18037
rect 552 17978 31531 18000
rect 552 17926 8102 17978
rect 8154 17926 8166 17978
rect 8218 17926 8230 17978
rect 8282 17926 8294 17978
rect 8346 17926 8358 17978
rect 8410 17926 15807 17978
rect 15859 17926 15871 17978
rect 15923 17926 15935 17978
rect 15987 17926 15999 17978
rect 16051 17926 16063 17978
rect 16115 17926 23512 17978
rect 23564 17926 23576 17978
rect 23628 17926 23640 17978
rect 23692 17926 23704 17978
rect 23756 17926 23768 17978
rect 23820 17926 31217 17978
rect 31269 17926 31281 17978
rect 31333 17926 31345 17978
rect 31397 17926 31409 17978
rect 31461 17926 31473 17978
rect 31525 17926 31531 17978
rect 552 17904 31531 17926
rect 6733 17867 6791 17873
rect 6733 17833 6745 17867
rect 6779 17864 6791 17867
rect 7098 17864 7104 17876
rect 6779 17836 7104 17864
rect 6779 17833 6791 17836
rect 6733 17827 6791 17833
rect 6549 17731 6607 17737
rect 6549 17697 6561 17731
rect 6595 17728 6607 17731
rect 6748 17728 6776 17827
rect 7098 17824 7104 17836
rect 7156 17864 7162 17876
rect 7377 17867 7435 17873
rect 7377 17864 7389 17867
rect 7156 17836 7389 17864
rect 7156 17824 7162 17836
rect 7377 17833 7389 17836
rect 7423 17833 7435 17867
rect 7377 17827 7435 17833
rect 12250 17824 12256 17876
rect 12308 17824 12314 17876
rect 12805 17867 12863 17873
rect 12805 17833 12817 17867
rect 12851 17864 12863 17867
rect 12986 17864 12992 17876
rect 12851 17836 12992 17864
rect 12851 17833 12863 17836
rect 12805 17827 12863 17833
rect 8570 17805 8576 17808
rect 7653 17799 7711 17805
rect 7653 17796 7665 17799
rect 7116 17768 7665 17796
rect 7116 17737 7144 17768
rect 7653 17765 7665 17768
rect 7699 17796 7711 17799
rect 8542 17799 8576 17805
rect 8542 17796 8554 17799
rect 7699 17768 8554 17796
rect 7699 17765 7711 17768
rect 7653 17759 7711 17765
rect 8542 17765 8554 17768
rect 8542 17759 8576 17765
rect 8570 17756 8576 17759
rect 8628 17756 8634 17808
rect 6595 17700 6776 17728
rect 6825 17731 6883 17737
rect 6595 17697 6607 17700
rect 6549 17691 6607 17697
rect 6825 17697 6837 17731
rect 6871 17728 6883 17731
rect 7101 17731 7159 17737
rect 7101 17728 7113 17731
rect 6871 17700 7113 17728
rect 6871 17697 6883 17700
rect 6825 17691 6883 17697
rect 7101 17697 7113 17700
rect 7147 17697 7159 17731
rect 7101 17691 7159 17697
rect 7469 17731 7527 17737
rect 7469 17697 7481 17731
rect 7515 17697 7527 17731
rect 7469 17691 7527 17697
rect 7484 17660 7512 17691
rect 7742 17688 7748 17740
rect 7800 17728 7806 17740
rect 7837 17731 7895 17737
rect 7837 17728 7849 17731
rect 7800 17700 7849 17728
rect 7800 17688 7806 17700
rect 7837 17697 7849 17700
rect 7883 17697 7895 17731
rect 7837 17691 7895 17697
rect 7926 17688 7932 17740
rect 7984 17688 7990 17740
rect 7944 17660 7972 17688
rect 7484 17632 7972 17660
rect 8018 17620 8024 17672
rect 8076 17660 8082 17672
rect 8297 17663 8355 17669
rect 8297 17660 8309 17663
rect 8076 17632 8309 17660
rect 8076 17620 8082 17632
rect 8297 17629 8309 17632
rect 8343 17629 8355 17663
rect 12268 17660 12296 17824
rect 12342 17688 12348 17740
rect 12400 17688 12406 17740
rect 12621 17731 12679 17737
rect 12621 17697 12633 17731
rect 12667 17728 12679 17731
rect 12820 17728 12848 17827
rect 12986 17824 12992 17836
rect 13044 17864 13050 17876
rect 13081 17867 13139 17873
rect 13081 17864 13093 17867
rect 13044 17836 13093 17864
rect 13044 17824 13050 17836
rect 13081 17833 13093 17836
rect 13127 17833 13139 17867
rect 13081 17827 13139 17833
rect 13354 17824 13360 17876
rect 13412 17824 13418 17876
rect 13722 17824 13728 17876
rect 13780 17824 13786 17876
rect 16209 17867 16267 17873
rect 16209 17833 16221 17867
rect 16255 17864 16267 17867
rect 16255 17836 19104 17864
rect 16255 17833 16267 17836
rect 16209 17827 16267 17833
rect 13740 17796 13768 17824
rect 13878 17799 13936 17805
rect 13878 17796 13890 17799
rect 13740 17768 13890 17796
rect 12667 17700 12848 17728
rect 12667 17697 12679 17700
rect 12621 17691 12679 17697
rect 12894 17688 12900 17740
rect 12952 17688 12958 17740
rect 12986 17688 12992 17740
rect 13044 17728 13050 17740
rect 13173 17731 13231 17737
rect 13173 17728 13185 17731
rect 13044 17700 13185 17728
rect 13044 17688 13050 17700
rect 13173 17697 13185 17700
rect 13219 17728 13231 17731
rect 13265 17731 13323 17737
rect 13265 17728 13277 17731
rect 13219 17700 13277 17728
rect 13219 17697 13231 17700
rect 13173 17691 13231 17697
rect 13265 17697 13277 17700
rect 13311 17697 13323 17731
rect 13265 17691 13323 17697
rect 13630 17688 13636 17740
rect 13688 17688 13694 17740
rect 12529 17663 12587 17669
rect 12529 17660 12541 17663
rect 12268 17632 12541 17660
rect 8297 17623 8355 17629
rect 12529 17629 12541 17632
rect 12575 17660 12587 17663
rect 13740 17660 13768 17768
rect 13878 17765 13890 17768
rect 13924 17765 13936 17799
rect 13878 17759 13936 17765
rect 16482 17756 16488 17808
rect 16540 17756 16546 17808
rect 16206 17688 16212 17740
rect 16264 17688 16270 17740
rect 16301 17731 16359 17737
rect 16301 17697 16313 17731
rect 16347 17728 16359 17731
rect 16500 17728 16528 17756
rect 16347 17700 16528 17728
rect 16592 17728 16620 17836
rect 18690 17756 18696 17808
rect 18748 17756 18754 17808
rect 19076 17796 19104 17836
rect 24302 17824 24308 17876
rect 24360 17864 24366 17876
rect 24581 17867 24639 17873
rect 24581 17864 24593 17867
rect 24360 17836 24593 17864
rect 24360 17824 24366 17836
rect 24581 17833 24593 17836
rect 24627 17833 24639 17867
rect 24581 17827 24639 17833
rect 24946 17824 24952 17876
rect 25004 17864 25010 17876
rect 25501 17867 25559 17873
rect 25501 17864 25513 17867
rect 25004 17836 25513 17864
rect 25004 17824 25010 17836
rect 25501 17833 25513 17836
rect 25547 17864 25559 17867
rect 25547 17836 25912 17864
rect 25547 17833 25559 17836
rect 25501 17827 25559 17833
rect 19242 17796 19248 17808
rect 19076 17768 19248 17796
rect 16649 17731 16707 17737
rect 16649 17728 16661 17731
rect 16592 17700 16661 17728
rect 16347 17697 16359 17700
rect 16301 17691 16359 17697
rect 16649 17697 16661 17700
rect 16695 17697 16707 17731
rect 16649 17691 16707 17697
rect 16942 17688 16948 17740
rect 17000 17728 17006 17740
rect 17865 17731 17923 17737
rect 17865 17728 17877 17731
rect 17000 17700 17877 17728
rect 17000 17688 17006 17700
rect 17865 17697 17877 17700
rect 17911 17697 17923 17731
rect 17865 17691 17923 17697
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17728 18659 17731
rect 18708 17728 18736 17756
rect 19076 17737 19104 17768
rect 19242 17756 19248 17768
rect 19300 17796 19306 17808
rect 19300 17768 19472 17796
rect 19300 17756 19306 17768
rect 19444 17737 19472 17768
rect 22370 17756 22376 17808
rect 22428 17805 22434 17808
rect 22428 17796 22440 17805
rect 22428 17768 22473 17796
rect 22428 17759 22440 17768
rect 22428 17756 22434 17759
rect 22830 17756 22836 17808
rect 22888 17796 22894 17808
rect 23854 17799 23912 17805
rect 23854 17796 23866 17799
rect 22888 17768 23866 17796
rect 22888 17756 22894 17768
rect 23854 17765 23866 17768
rect 23900 17796 23912 17799
rect 25225 17799 25283 17805
rect 25225 17796 25237 17799
rect 23900 17768 24716 17796
rect 23900 17765 23912 17768
rect 23854 17759 23912 17765
rect 18647 17700 18736 17728
rect 19061 17731 19119 17737
rect 18647 17697 18659 17700
rect 18601 17691 18659 17697
rect 19061 17697 19073 17731
rect 19107 17697 19119 17731
rect 19061 17691 19119 17697
rect 19337 17731 19395 17737
rect 19337 17697 19349 17731
rect 19383 17697 19395 17731
rect 19337 17691 19395 17697
rect 19429 17731 19487 17737
rect 19429 17697 19441 17731
rect 19475 17697 19487 17731
rect 19429 17691 19487 17697
rect 19705 17731 19763 17737
rect 19705 17697 19717 17731
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 12575 17632 13768 17660
rect 16224 17660 16252 17688
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 16224 17632 16405 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 16393 17629 16405 17632
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17660 18751 17663
rect 18969 17663 19027 17669
rect 18969 17660 18981 17663
rect 18739 17632 18981 17660
rect 18739 17629 18751 17632
rect 18693 17623 18751 17629
rect 18969 17629 18981 17632
rect 19015 17660 19027 17663
rect 19352 17660 19380 17691
rect 19720 17660 19748 17691
rect 21910 17688 21916 17740
rect 21968 17728 21974 17740
rect 22649 17731 22707 17737
rect 22649 17728 22661 17731
rect 21968 17700 22661 17728
rect 21968 17688 21974 17700
rect 22649 17697 22661 17700
rect 22695 17697 22707 17731
rect 22649 17691 22707 17697
rect 24302 17688 24308 17740
rect 24360 17728 24366 17740
rect 24688 17737 24716 17768
rect 24826 17768 25237 17796
rect 24397 17731 24455 17737
rect 24397 17728 24409 17731
rect 24360 17700 24409 17728
rect 24360 17688 24366 17700
rect 24397 17697 24409 17700
rect 24443 17697 24455 17731
rect 24397 17691 24455 17697
rect 24673 17731 24731 17737
rect 24673 17697 24685 17731
rect 24719 17728 24731 17731
rect 24826 17728 24854 17768
rect 25225 17765 25237 17768
rect 25271 17796 25283 17799
rect 25777 17799 25835 17805
rect 25777 17796 25789 17799
rect 25271 17768 25789 17796
rect 25271 17765 25283 17768
rect 25225 17759 25283 17765
rect 25777 17765 25789 17768
rect 25823 17765 25835 17799
rect 25777 17759 25835 17765
rect 24719 17700 24854 17728
rect 24719 17697 24731 17700
rect 24673 17691 24731 17697
rect 25314 17688 25320 17740
rect 25372 17688 25378 17740
rect 25590 17688 25596 17740
rect 25648 17688 25654 17740
rect 25884 17737 25912 17836
rect 25869 17731 25927 17737
rect 25869 17697 25881 17731
rect 25915 17728 25927 17731
rect 26053 17731 26111 17737
rect 26053 17728 26065 17731
rect 25915 17700 26065 17728
rect 25915 17697 25927 17700
rect 25869 17691 25927 17697
rect 26053 17697 26065 17700
rect 26099 17697 26111 17731
rect 26053 17691 26111 17697
rect 26142 17688 26148 17740
rect 26200 17688 26206 17740
rect 19015 17632 19748 17660
rect 24121 17663 24179 17669
rect 19015 17629 19027 17632
rect 18969 17623 19027 17629
rect 24121 17629 24133 17663
rect 24167 17660 24179 17663
rect 25222 17660 25228 17672
rect 24167 17632 25228 17660
rect 24167 17629 24179 17632
rect 24121 17623 24179 17629
rect 17957 17595 18015 17601
rect 9692 17564 12434 17592
rect 6454 17484 6460 17536
rect 6512 17484 6518 17536
rect 7006 17484 7012 17536
rect 7064 17484 7070 17536
rect 7926 17484 7932 17536
rect 7984 17484 7990 17536
rect 9692 17533 9720 17564
rect 9677 17527 9735 17533
rect 9677 17493 9689 17527
rect 9723 17493 9735 17527
rect 12406 17524 12434 17564
rect 14568 17564 15700 17592
rect 14568 17524 14596 17564
rect 15672 17536 15700 17564
rect 17957 17561 17969 17595
rect 18003 17592 18015 17595
rect 18003 17564 19840 17592
rect 18003 17561 18015 17564
rect 17957 17555 18015 17561
rect 12406 17496 14596 17524
rect 9677 17487 9735 17493
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 15013 17527 15071 17533
rect 15013 17524 15025 17527
rect 14700 17496 15025 17524
rect 14700 17484 14706 17496
rect 15013 17493 15025 17496
rect 15059 17493 15071 17527
rect 15013 17487 15071 17493
rect 15654 17484 15660 17536
rect 15712 17484 15718 17536
rect 17770 17484 17776 17536
rect 17828 17484 17834 17536
rect 19242 17484 19248 17536
rect 19300 17484 19306 17536
rect 19518 17484 19524 17536
rect 19576 17484 19582 17536
rect 19812 17533 19840 17564
rect 19797 17527 19855 17533
rect 19797 17493 19809 17527
rect 19843 17524 19855 17527
rect 19978 17524 19984 17536
rect 19843 17496 19984 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 19978 17484 19984 17496
rect 20036 17484 20042 17536
rect 21266 17484 21272 17536
rect 21324 17484 21330 17536
rect 22741 17527 22799 17533
rect 22741 17493 22753 17527
rect 22787 17524 22799 17527
rect 23198 17524 23204 17536
rect 22787 17496 23204 17524
rect 22787 17493 22799 17496
rect 22741 17487 22799 17493
rect 23198 17484 23204 17496
rect 23256 17484 23262 17536
rect 23842 17484 23848 17536
rect 23900 17524 23906 17536
rect 24136 17524 24164 17623
rect 25222 17620 25228 17632
rect 25280 17620 25286 17672
rect 23900 17496 24164 17524
rect 23900 17484 23906 17496
rect 552 17434 31372 17456
rect 552 17382 4250 17434
rect 4302 17382 4314 17434
rect 4366 17382 4378 17434
rect 4430 17382 4442 17434
rect 4494 17382 4506 17434
rect 4558 17382 11955 17434
rect 12007 17382 12019 17434
rect 12071 17382 12083 17434
rect 12135 17382 12147 17434
rect 12199 17382 12211 17434
rect 12263 17382 19660 17434
rect 19712 17382 19724 17434
rect 19776 17382 19788 17434
rect 19840 17382 19852 17434
rect 19904 17382 19916 17434
rect 19968 17382 27365 17434
rect 27417 17382 27429 17434
rect 27481 17382 27493 17434
rect 27545 17382 27557 17434
rect 27609 17382 27621 17434
rect 27673 17382 31372 17434
rect 552 17360 31372 17382
rect 6454 17280 6460 17332
rect 6512 17320 6518 17332
rect 6733 17323 6791 17329
rect 6733 17320 6745 17323
rect 6512 17292 6745 17320
rect 6512 17280 6518 17292
rect 6733 17289 6745 17292
rect 6779 17289 6791 17323
rect 6733 17283 6791 17289
rect 7006 17280 7012 17332
rect 7064 17320 7070 17332
rect 7285 17323 7343 17329
rect 7285 17320 7297 17323
rect 7064 17292 7297 17320
rect 7064 17280 7070 17292
rect 5077 17255 5135 17261
rect 5077 17221 5089 17255
rect 5123 17252 5135 17255
rect 5994 17252 6000 17264
rect 5123 17224 6000 17252
rect 5123 17221 5135 17224
rect 5077 17215 5135 17221
rect 5994 17212 6000 17224
rect 6052 17212 6058 17264
rect 6472 17252 6500 17280
rect 6104 17224 6500 17252
rect 5626 17184 5632 17196
rect 5460 17156 5632 17184
rect 842 17076 848 17128
rect 900 17076 906 17128
rect 3697 17119 3755 17125
rect 3697 17085 3709 17119
rect 3743 17116 3755 17119
rect 5460 17116 5488 17156
rect 5626 17144 5632 17156
rect 5684 17144 5690 17196
rect 6104 17125 6132 17224
rect 7116 17125 7144 17292
rect 7285 17289 7297 17292
rect 7331 17289 7343 17323
rect 7285 17283 7343 17289
rect 11793 17323 11851 17329
rect 11793 17289 11805 17323
rect 11839 17320 11851 17323
rect 12069 17323 12127 17329
rect 12069 17320 12081 17323
rect 11839 17292 12081 17320
rect 11839 17289 11851 17292
rect 11793 17283 11851 17289
rect 12069 17289 12081 17292
rect 12115 17320 12127 17323
rect 12342 17320 12348 17332
rect 12115 17292 12348 17320
rect 12115 17289 12127 17292
rect 12069 17283 12127 17289
rect 3743 17088 5488 17116
rect 5537 17119 5595 17125
rect 3743 17085 3755 17088
rect 3697 17079 3755 17085
rect 5537 17085 5549 17119
rect 5583 17116 5595 17119
rect 5813 17119 5871 17125
rect 5813 17116 5825 17119
rect 5583 17088 5825 17116
rect 5583 17085 5595 17088
rect 5537 17079 5595 17085
rect 5813 17085 5825 17088
rect 5859 17116 5871 17119
rect 6089 17119 6147 17125
rect 5859 17088 6040 17116
rect 5859 17085 5871 17088
rect 5813 17079 5871 17085
rect 6012 17057 6040 17088
rect 6089 17085 6101 17119
rect 6135 17085 6147 17119
rect 6089 17079 6147 17085
rect 6365 17119 6423 17125
rect 6365 17085 6377 17119
rect 6411 17085 6423 17119
rect 6365 17079 6423 17085
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 7101 17119 7159 17125
rect 7101 17116 7113 17119
rect 6871 17088 7113 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 7101 17085 7113 17088
rect 7147 17085 7159 17119
rect 7101 17079 7159 17085
rect 3964 17051 4022 17057
rect 3964 17017 3976 17051
rect 4010 17048 4022 17051
rect 5997 17051 6055 17057
rect 4010 17020 5488 17048
rect 4010 17017 4022 17020
rect 3964 17011 4022 17017
rect 5460 16992 5488 17020
rect 5997 17017 6009 17051
rect 6043 17048 6055 17051
rect 6273 17051 6331 17057
rect 6273 17048 6285 17051
rect 6043 17020 6285 17048
rect 6043 17017 6055 17020
rect 5997 17011 6055 17017
rect 6273 17017 6285 17020
rect 6319 17017 6331 17051
rect 6380 17048 6408 17079
rect 7374 17076 7380 17128
rect 7432 17116 7438 17128
rect 7926 17116 7932 17128
rect 7432 17088 7932 17116
rect 7432 17076 7438 17088
rect 7926 17076 7932 17088
rect 7984 17076 7990 17128
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17116 9735 17119
rect 9766 17116 9772 17128
rect 9723 17088 9772 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 9766 17076 9772 17088
rect 9824 17116 9830 17128
rect 10778 17116 10784 17128
rect 9824 17088 10784 17116
rect 9824 17076 9830 17088
rect 10778 17076 10784 17088
rect 10836 17076 10842 17128
rect 7392 17048 7420 17076
rect 6380 17020 7420 17048
rect 6273 17011 6331 17017
rect 9214 17008 9220 17060
rect 9272 17048 9278 17060
rect 9922 17051 9980 17057
rect 9922 17048 9934 17051
rect 9272 17020 9934 17048
rect 9272 17008 9278 17020
rect 9922 17017 9934 17020
rect 9968 17017 9980 17051
rect 11808 17048 11836 17283
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 19429 17323 19487 17329
rect 19429 17289 19441 17323
rect 19475 17320 19487 17323
rect 19518 17320 19524 17332
rect 19475 17292 19524 17320
rect 19475 17289 19487 17292
rect 19429 17283 19487 17289
rect 19518 17280 19524 17292
rect 19576 17280 19582 17332
rect 21910 17320 21916 17332
rect 19628 17292 21916 17320
rect 12802 17252 12808 17264
rect 12406 17224 12808 17252
rect 12406 17184 12434 17224
rect 12636 17193 12664 17224
rect 12802 17212 12808 17224
rect 12860 17212 12866 17264
rect 16117 17255 16175 17261
rect 16117 17221 16129 17255
rect 16163 17252 16175 17255
rect 16850 17252 16856 17264
rect 16163 17224 16856 17252
rect 16163 17221 16175 17224
rect 16117 17215 16175 17221
rect 16850 17212 16856 17224
rect 16908 17212 16914 17264
rect 19628 17252 19656 17292
rect 19306 17224 19656 17252
rect 19705 17255 19763 17261
rect 11900 17156 12434 17184
rect 12621 17187 12679 17193
rect 11900 17128 11928 17156
rect 12621 17153 12633 17187
rect 12667 17184 12679 17187
rect 12667 17156 13232 17184
rect 12667 17153 12679 17156
rect 12621 17147 12679 17153
rect 11882 17076 11888 17128
rect 11940 17076 11946 17128
rect 12158 17076 12164 17128
rect 12216 17076 12222 17128
rect 12253 17119 12311 17125
rect 12253 17085 12265 17119
rect 12299 17116 12311 17119
rect 12434 17116 12440 17128
rect 12299 17088 12440 17116
rect 12299 17085 12311 17088
rect 12253 17079 12311 17085
rect 12434 17076 12440 17088
rect 12492 17116 12498 17128
rect 12529 17119 12587 17125
rect 12529 17116 12541 17119
rect 12492 17088 12541 17116
rect 12492 17076 12498 17088
rect 12529 17085 12541 17088
rect 12575 17085 12587 17119
rect 12529 17079 12587 17085
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17085 12863 17119
rect 13204 17116 13232 17156
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 13688 17156 14749 17184
rect 13688 17144 13694 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 17862 17144 17868 17196
rect 17920 17184 17926 17196
rect 19306 17184 19334 17224
rect 19705 17221 19717 17255
rect 19751 17252 19763 17255
rect 20257 17255 20315 17261
rect 20257 17252 20269 17255
rect 19751 17224 20269 17252
rect 19751 17221 19763 17224
rect 19705 17215 19763 17221
rect 20257 17221 20269 17224
rect 20303 17252 20315 17255
rect 20438 17252 20444 17264
rect 20303 17224 20444 17252
rect 20303 17221 20315 17224
rect 20257 17215 20315 17221
rect 20438 17212 20444 17224
rect 20496 17252 20502 17264
rect 20496 17224 20760 17252
rect 20496 17212 20502 17224
rect 17920 17156 19334 17184
rect 17920 17144 17926 17156
rect 19518 17144 19524 17196
rect 19576 17184 19582 17196
rect 19576 17156 20484 17184
rect 19576 17144 19582 17156
rect 14993 17119 15051 17125
rect 14993 17116 15005 17119
rect 13204 17088 15005 17116
rect 12805 17079 12863 17085
rect 14993 17085 15005 17088
rect 15039 17085 15051 17119
rect 14993 17079 15051 17085
rect 17609 17119 17667 17125
rect 17609 17085 17621 17119
rect 17655 17116 17667 17119
rect 19337 17119 19395 17125
rect 19337 17116 19349 17119
rect 17655 17088 19349 17116
rect 17655 17085 17667 17088
rect 17609 17079 17667 17085
rect 19337 17085 19349 17088
rect 19383 17116 19395 17119
rect 19613 17119 19671 17125
rect 19613 17116 19625 17119
rect 19383 17088 19625 17116
rect 19383 17085 19395 17088
rect 19337 17079 19395 17085
rect 19613 17085 19625 17088
rect 19659 17116 19671 17119
rect 19978 17116 19984 17128
rect 19659 17088 19984 17116
rect 19659 17085 19671 17088
rect 19613 17079 19671 17085
rect 12820 17048 12848 17079
rect 19978 17076 19984 17088
rect 20036 17076 20042 17128
rect 20088 17125 20116 17156
rect 20456 17125 20484 17156
rect 20732 17125 20760 17224
rect 21744 17193 21772 17292
rect 21910 17280 21916 17292
rect 21968 17280 21974 17332
rect 25041 17323 25099 17329
rect 25041 17289 25053 17323
rect 25087 17320 25099 17323
rect 25314 17320 25320 17332
rect 25087 17292 25320 17320
rect 25087 17289 25099 17292
rect 25041 17283 25099 17289
rect 25314 17280 25320 17292
rect 25372 17280 25378 17332
rect 25240 17224 26188 17252
rect 21729 17187 21787 17193
rect 21729 17153 21741 17187
rect 21775 17153 21787 17187
rect 21729 17147 21787 17153
rect 20073 17119 20131 17125
rect 20073 17085 20085 17119
rect 20119 17085 20131 17119
rect 20165 17119 20223 17125
rect 20165 17118 20177 17119
rect 20073 17079 20131 17085
rect 20164 17085 20177 17118
rect 20211 17085 20223 17119
rect 20164 17079 20223 17085
rect 20441 17119 20499 17125
rect 20441 17085 20453 17119
rect 20487 17085 20499 17119
rect 20441 17079 20499 17085
rect 20717 17119 20775 17125
rect 20717 17085 20729 17119
rect 20763 17085 20775 17119
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 20717 17079 20775 17085
rect 20824 17088 21189 17116
rect 20164 17048 20192 17079
rect 20824 17057 20852 17088
rect 21177 17085 21189 17088
rect 21223 17116 21235 17119
rect 21453 17119 21511 17125
rect 21453 17116 21465 17119
rect 21223 17088 21465 17116
rect 21223 17085 21235 17088
rect 21177 17079 21235 17085
rect 21453 17085 21465 17088
rect 21499 17085 21511 17119
rect 21453 17079 21511 17085
rect 25133 17119 25191 17125
rect 25133 17085 25145 17119
rect 25179 17116 25191 17119
rect 25240 17116 25268 17224
rect 25314 17144 25320 17196
rect 25372 17144 25378 17196
rect 25700 17156 26096 17184
rect 25179 17088 25268 17116
rect 25179 17085 25191 17088
rect 25133 17079 25191 17085
rect 11808 17020 12848 17048
rect 19996 17020 20192 17048
rect 20533 17051 20591 17057
rect 9922 17011 9980 17017
rect 5442 16940 5448 16992
rect 5500 16940 5506 16992
rect 5718 16940 5724 16992
rect 5776 16980 5782 16992
rect 7009 16983 7067 16989
rect 7009 16980 7021 16983
rect 5776 16952 7021 16980
rect 5776 16940 5782 16952
rect 7009 16949 7021 16952
rect 7055 16980 7067 16983
rect 8478 16980 8484 16992
rect 7055 16952 8484 16980
rect 7055 16949 7067 16952
rect 7009 16943 7067 16949
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 11057 16983 11115 16989
rect 11057 16949 11069 16983
rect 11103 16980 11115 16983
rect 11698 16980 11704 16992
rect 11103 16952 11704 16980
rect 11103 16949 11115 16952
rect 11057 16943 11115 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 12345 16983 12403 16989
rect 12345 16949 12357 16983
rect 12391 16980 12403 16983
rect 12894 16980 12900 16992
rect 12391 16952 12900 16980
rect 12391 16949 12403 16952
rect 12345 16943 12403 16949
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 16485 16983 16543 16989
rect 16485 16949 16497 16983
rect 16531 16980 16543 16983
rect 17402 16980 17408 16992
rect 16531 16952 17408 16980
rect 16531 16949 16543 16952
rect 16485 16943 16543 16949
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 19242 16940 19248 16992
rect 19300 16980 19306 16992
rect 19996 16989 20024 17020
rect 20533 17017 20545 17051
rect 20579 17048 20591 17051
rect 20809 17051 20867 17057
rect 20809 17048 20821 17051
rect 20579 17020 20821 17048
rect 20579 17017 20591 17020
rect 20533 17011 20591 17017
rect 20809 17017 20821 17020
rect 20855 17017 20867 17051
rect 21468 17048 21496 17079
rect 21974 17051 22032 17057
rect 21974 17048 21986 17051
rect 21468 17020 21986 17048
rect 20809 17011 20867 17017
rect 21974 17017 21986 17020
rect 22020 17017 22032 17051
rect 21974 17011 22032 17017
rect 24302 17008 24308 17060
rect 24360 17008 24366 17060
rect 25332 17048 25360 17144
rect 25700 17128 25728 17156
rect 25406 17076 25412 17128
rect 25464 17076 25470 17128
rect 25682 17076 25688 17128
rect 25740 17076 25746 17128
rect 26068 17125 26096 17156
rect 25777 17119 25835 17125
rect 25777 17085 25789 17119
rect 25823 17085 25835 17119
rect 25777 17079 25835 17085
rect 26053 17119 26111 17125
rect 26053 17085 26065 17119
rect 26099 17085 26111 17119
rect 26053 17079 26111 17085
rect 25792 17048 25820 17079
rect 26160 17060 26188 17224
rect 27062 17076 27068 17128
rect 27120 17116 27126 17128
rect 27709 17119 27767 17125
rect 27709 17116 27721 17119
rect 27120 17088 27721 17116
rect 27120 17076 27126 17088
rect 27709 17085 27721 17088
rect 27755 17116 27767 17119
rect 27755 17088 30052 17116
rect 27755 17085 27767 17088
rect 27709 17079 27767 17085
rect 25332 17020 25820 17048
rect 26142 17008 26148 17060
rect 26200 17048 26206 17060
rect 27430 17048 27436 17060
rect 27488 17057 27494 17060
rect 26200 17020 27436 17048
rect 26200 17008 26206 17020
rect 27430 17008 27436 17020
rect 27488 17048 27500 17057
rect 27488 17020 27533 17048
rect 27488 17011 27500 17020
rect 27488 17008 27494 17011
rect 19981 16983 20039 16989
rect 19981 16980 19993 16983
rect 19300 16952 19993 16980
rect 19300 16940 19306 16952
rect 19981 16949 19993 16952
rect 20027 16949 20039 16983
rect 19981 16943 20039 16949
rect 21082 16940 21088 16992
rect 21140 16940 21146 16992
rect 21542 16940 21548 16992
rect 21600 16940 21606 16992
rect 23106 16940 23112 16992
rect 23164 16940 23170 16992
rect 24320 16980 24348 17008
rect 30024 16992 30052 17088
rect 25590 16980 25596 16992
rect 24320 16952 25596 16980
rect 25590 16940 25596 16952
rect 25648 16980 25654 16992
rect 25869 16983 25927 16989
rect 25869 16980 25881 16983
rect 25648 16952 25881 16980
rect 25648 16940 25654 16952
rect 25869 16949 25881 16952
rect 25915 16949 25927 16983
rect 25869 16943 25927 16949
rect 26326 16940 26332 16992
rect 26384 16940 26390 16992
rect 30006 16940 30012 16992
rect 30064 16940 30070 16992
rect 552 16890 31531 16912
rect 552 16838 8102 16890
rect 8154 16838 8166 16890
rect 8218 16838 8230 16890
rect 8282 16838 8294 16890
rect 8346 16838 8358 16890
rect 8410 16838 15807 16890
rect 15859 16838 15871 16890
rect 15923 16838 15935 16890
rect 15987 16838 15999 16890
rect 16051 16838 16063 16890
rect 16115 16838 23512 16890
rect 23564 16838 23576 16890
rect 23628 16838 23640 16890
rect 23692 16838 23704 16890
rect 23756 16838 23768 16890
rect 23820 16838 31217 16890
rect 31269 16838 31281 16890
rect 31333 16838 31345 16890
rect 31397 16838 31409 16890
rect 31461 16838 31473 16890
rect 31525 16838 31531 16890
rect 552 16816 31531 16838
rect 5261 16779 5319 16785
rect 5261 16745 5273 16779
rect 5307 16776 5319 16779
rect 5442 16776 5448 16788
rect 5307 16748 5448 16776
rect 5307 16745 5319 16748
rect 5261 16739 5319 16745
rect 5276 16708 5304 16739
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 6546 16776 6552 16788
rect 6289 16748 6552 16776
rect 5537 16711 5595 16717
rect 5537 16708 5549 16711
rect 3804 16680 5304 16708
rect 5368 16680 5549 16708
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 2406 16640 2412 16652
rect 2087 16612 2412 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 2406 16600 2412 16612
rect 2464 16600 2470 16652
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 3804 16649 3832 16680
rect 5368 16649 5396 16680
rect 5537 16677 5549 16680
rect 5583 16708 5595 16711
rect 5583 16680 6040 16708
rect 5583 16677 5595 16680
rect 5537 16671 5595 16677
rect 3697 16643 3755 16649
rect 3292 16612 3648 16640
rect 3292 16600 3298 16612
rect 3620 16572 3648 16612
rect 3697 16609 3709 16643
rect 3743 16640 3755 16643
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3743 16612 3801 16640
rect 3743 16609 3755 16612
rect 3697 16603 3755 16609
rect 3789 16609 3801 16612
rect 3835 16609 3847 16643
rect 3789 16603 3847 16609
rect 3881 16643 3939 16649
rect 3881 16609 3893 16643
rect 3927 16640 3939 16643
rect 4249 16643 4307 16649
rect 4249 16640 4261 16643
rect 3927 16612 4261 16640
rect 3927 16609 3939 16612
rect 3881 16603 3939 16609
rect 4249 16609 4261 16612
rect 4295 16640 4307 16643
rect 4525 16643 4583 16649
rect 4525 16640 4537 16643
rect 4295 16612 4537 16640
rect 4295 16609 4307 16612
rect 4249 16603 4307 16609
rect 4525 16609 4537 16612
rect 4571 16640 4583 16643
rect 4801 16643 4859 16649
rect 4801 16640 4813 16643
rect 4571 16612 4813 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 4801 16609 4813 16612
rect 4847 16609 4859 16643
rect 4801 16603 4859 16609
rect 4893 16643 4951 16649
rect 4893 16609 4905 16643
rect 4939 16640 4951 16643
rect 5353 16643 5411 16649
rect 4939 16612 5304 16640
rect 4939 16609 4951 16612
rect 4893 16603 4951 16609
rect 5276 16572 5304 16612
rect 5353 16609 5365 16643
rect 5399 16609 5411 16643
rect 5629 16643 5687 16649
rect 5629 16640 5641 16643
rect 5353 16603 5411 16609
rect 5460 16612 5641 16640
rect 5460 16572 5488 16612
rect 5629 16609 5641 16612
rect 5675 16640 5687 16643
rect 5718 16640 5724 16652
rect 5675 16612 5724 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 5718 16600 5724 16612
rect 5776 16600 5782 16652
rect 6012 16649 6040 16680
rect 6289 16649 6317 16748
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 8018 16736 8024 16788
rect 8076 16736 8082 16788
rect 11793 16779 11851 16785
rect 11793 16745 11805 16779
rect 11839 16776 11851 16779
rect 11882 16776 11888 16788
rect 11839 16748 11888 16776
rect 11839 16745 11851 16748
rect 11793 16739 11851 16745
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12161 16779 12219 16785
rect 12161 16745 12173 16779
rect 12207 16776 12219 16779
rect 12434 16776 12440 16788
rect 12207 16748 12440 16776
rect 12207 16745 12219 16748
rect 12161 16739 12219 16745
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 12894 16736 12900 16788
rect 12952 16736 12958 16788
rect 20073 16779 20131 16785
rect 20073 16745 20085 16779
rect 20119 16776 20131 16779
rect 21082 16776 21088 16788
rect 20119 16748 21088 16776
rect 20119 16745 20131 16748
rect 20073 16739 20131 16745
rect 6454 16708 6460 16720
rect 6380 16680 6460 16708
rect 6380 16649 6408 16680
rect 6454 16668 6460 16680
rect 6512 16708 6518 16720
rect 8036 16708 8064 16736
rect 8386 16708 8392 16720
rect 6512 16680 8392 16708
rect 6512 16668 6518 16680
rect 8036 16649 8064 16680
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 12912 16708 12940 16736
rect 13418 16711 13476 16717
rect 13418 16708 13430 16711
rect 11440 16680 11744 16708
rect 12912 16680 13430 16708
rect 11440 16652 11468 16680
rect 5997 16643 6055 16649
rect 5997 16609 6009 16643
rect 6043 16640 6055 16643
rect 6181 16643 6239 16649
rect 6181 16640 6193 16643
rect 6043 16612 6193 16640
rect 6043 16609 6055 16612
rect 5997 16603 6055 16609
rect 6181 16609 6193 16612
rect 6227 16609 6239 16643
rect 6181 16603 6239 16609
rect 6273 16643 6331 16649
rect 6273 16609 6285 16643
rect 6319 16609 6331 16643
rect 6273 16603 6331 16609
rect 6365 16643 6423 16649
rect 6365 16609 6377 16643
rect 6411 16609 6423 16643
rect 6621 16643 6679 16649
rect 6621 16640 6633 16643
rect 6365 16603 6423 16609
rect 6472 16612 6633 16640
rect 3620 16544 4476 16572
rect 5276 16544 5488 16572
rect 6289 16572 6317 16603
rect 6472 16572 6500 16612
rect 6621 16609 6633 16612
rect 6667 16609 6679 16643
rect 6621 16603 6679 16609
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 8110 16600 8116 16652
rect 8168 16640 8174 16652
rect 8277 16643 8335 16649
rect 8277 16640 8289 16643
rect 8168 16612 8289 16640
rect 8168 16600 8174 16612
rect 8277 16609 8289 16612
rect 8323 16609 8335 16643
rect 8277 16603 8335 16609
rect 10134 16600 10140 16652
rect 10192 16600 10198 16652
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16640 11299 16643
rect 11422 16640 11428 16652
rect 11287 16612 11428 16640
rect 11287 16609 11299 16612
rect 11241 16603 11299 16609
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 11716 16649 11744 16680
rect 13418 16677 13430 16680
rect 13464 16677 13476 16711
rect 13418 16671 13476 16677
rect 13630 16668 13636 16720
rect 13688 16668 13694 16720
rect 18040 16711 18098 16717
rect 18040 16677 18052 16711
rect 18086 16708 18098 16711
rect 19242 16708 19248 16720
rect 18086 16680 19248 16708
rect 18086 16677 18098 16680
rect 18040 16671 18098 16677
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16609 11575 16643
rect 11517 16603 11575 16609
rect 11701 16643 11759 16649
rect 11701 16609 11713 16643
rect 11747 16609 11759 16643
rect 11701 16603 11759 16609
rect 6289 16544 6500 16572
rect 1946 16396 1952 16448
rect 2004 16396 2010 16448
rect 3329 16439 3387 16445
rect 3329 16405 3341 16439
rect 3375 16436 3387 16439
rect 3510 16436 3516 16448
rect 3375 16408 3516 16436
rect 3375 16405 3387 16408
rect 3329 16399 3387 16405
rect 3510 16396 3516 16408
rect 3568 16436 3574 16448
rect 3605 16439 3663 16445
rect 3605 16436 3617 16439
rect 3568 16408 3617 16436
rect 3568 16396 3574 16408
rect 3605 16405 3617 16408
rect 3651 16405 3663 16439
rect 3605 16399 3663 16405
rect 4154 16396 4160 16448
rect 4212 16396 4218 16448
rect 4448 16445 4476 16544
rect 11532 16504 11560 16603
rect 11790 16600 11796 16652
rect 11848 16640 11854 16652
rect 12069 16643 12127 16649
rect 12069 16640 12081 16643
rect 11848 16612 12081 16640
rect 11848 16600 11854 16612
rect 12069 16609 12081 16612
rect 12115 16609 12127 16643
rect 12069 16603 12127 16609
rect 12342 16600 12348 16652
rect 12400 16600 12406 16652
rect 13648 16640 13676 16668
rect 13188 16612 13676 16640
rect 17773 16643 17831 16649
rect 12618 16532 12624 16584
rect 12676 16572 12682 16584
rect 13188 16581 13216 16612
rect 17773 16609 17785 16643
rect 17819 16640 17831 16643
rect 17862 16640 17868 16652
rect 17819 16612 17868 16640
rect 17819 16609 17831 16612
rect 17773 16603 17831 16609
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 19260 16640 19288 16668
rect 19889 16643 19947 16649
rect 19260 16612 19748 16640
rect 13173 16575 13231 16581
rect 13173 16572 13185 16575
rect 12676 16544 13185 16572
rect 12676 16532 12682 16544
rect 13173 16541 13185 16544
rect 13219 16541 13231 16575
rect 19720 16572 19748 16612
rect 19889 16609 19901 16643
rect 19935 16640 19947 16643
rect 20088 16640 20116 16739
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 25682 16736 25688 16788
rect 25740 16776 25746 16788
rect 25961 16779 26019 16785
rect 25961 16776 25973 16779
rect 25740 16748 25973 16776
rect 25740 16736 25746 16748
rect 25961 16745 25973 16748
rect 26007 16745 26019 16779
rect 27154 16776 27160 16788
rect 25961 16739 26019 16745
rect 26252 16748 27160 16776
rect 20438 16668 20444 16720
rect 20496 16668 20502 16720
rect 19935 16612 20116 16640
rect 20165 16643 20223 16649
rect 19935 16609 19947 16612
rect 19889 16603 19947 16609
rect 20165 16609 20177 16643
rect 20211 16609 20223 16643
rect 20456 16639 20484 16668
rect 20165 16603 20223 16609
rect 20441 16633 20499 16639
rect 20180 16572 20208 16603
rect 20441 16599 20453 16633
rect 20487 16599 20499 16633
rect 20714 16600 20720 16652
rect 20772 16600 20778 16652
rect 21100 16640 21128 16736
rect 25424 16680 26004 16708
rect 25424 16652 25452 16680
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 21100 16612 21281 16640
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 21542 16600 21548 16652
rect 21600 16640 21606 16652
rect 21729 16643 21787 16649
rect 21729 16640 21741 16643
rect 21600 16612 21741 16640
rect 21600 16600 21606 16612
rect 21729 16609 21741 16612
rect 21775 16640 21787 16643
rect 22005 16643 22063 16649
rect 22005 16640 22017 16643
rect 21775 16612 22017 16640
rect 21775 16609 21787 16612
rect 21729 16603 21787 16609
rect 22005 16609 22017 16612
rect 22051 16640 22063 16643
rect 22189 16643 22247 16649
rect 22189 16640 22201 16643
rect 22051 16612 22201 16640
rect 22051 16609 22063 16612
rect 22005 16603 22063 16609
rect 22189 16609 22201 16612
rect 22235 16609 22247 16643
rect 22189 16603 22247 16609
rect 22281 16643 22339 16649
rect 22281 16609 22293 16643
rect 22327 16640 22339 16643
rect 22370 16640 22376 16652
rect 22327 16612 22376 16640
rect 22327 16609 22339 16612
rect 22281 16603 22339 16609
rect 20441 16593 20499 16599
rect 22296 16572 22324 16603
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 23569 16643 23627 16649
rect 23569 16609 23581 16643
rect 23615 16640 23627 16643
rect 23658 16640 23664 16652
rect 23615 16612 23664 16640
rect 23615 16609 23627 16612
rect 23569 16603 23627 16609
rect 23658 16600 23664 16612
rect 23716 16600 23722 16652
rect 23836 16643 23894 16649
rect 23836 16609 23848 16643
rect 23882 16640 23894 16643
rect 24302 16640 24308 16652
rect 23882 16612 24308 16640
rect 23882 16609 23894 16612
rect 23836 16603 23894 16609
rect 24302 16600 24308 16612
rect 24360 16600 24366 16652
rect 25406 16600 25412 16652
rect 25464 16600 25470 16652
rect 25777 16643 25835 16649
rect 25777 16609 25789 16643
rect 25823 16609 25835 16643
rect 25976 16638 26004 16680
rect 26053 16643 26111 16649
rect 26053 16638 26065 16643
rect 25976 16610 26065 16638
rect 25777 16603 25835 16609
rect 26053 16609 26065 16610
rect 26099 16638 26111 16643
rect 26252 16638 26280 16748
rect 27154 16736 27160 16748
rect 27212 16736 27218 16788
rect 27985 16711 28043 16717
rect 27985 16708 27997 16711
rect 26804 16680 27997 16708
rect 26804 16649 26832 16680
rect 27985 16677 27997 16680
rect 28031 16677 28043 16711
rect 27985 16671 28043 16677
rect 26099 16610 26280 16638
rect 26789 16643 26847 16649
rect 26099 16609 26111 16610
rect 26053 16603 26111 16609
rect 26789 16609 26801 16643
rect 26835 16609 26847 16643
rect 27249 16643 27307 16649
rect 27249 16640 27261 16643
rect 26789 16603 26847 16609
rect 26896 16612 27261 16640
rect 19720 16544 20208 16572
rect 20999 16544 22324 16572
rect 25792 16572 25820 16603
rect 26418 16572 26424 16584
rect 25792 16544 26424 16572
rect 13173 16535 13231 16541
rect 11790 16504 11796 16516
rect 11532 16476 11796 16504
rect 11790 16464 11796 16476
rect 11848 16464 11854 16516
rect 19426 16504 19432 16516
rect 19076 16476 19432 16504
rect 4433 16439 4491 16445
rect 4433 16405 4445 16439
rect 4479 16436 4491 16439
rect 5905 16439 5963 16445
rect 5905 16436 5917 16439
rect 4479 16408 5917 16436
rect 4479 16405 4491 16408
rect 4433 16399 4491 16405
rect 5905 16405 5917 16408
rect 5951 16436 5963 16439
rect 6546 16436 6552 16448
rect 5951 16408 6552 16436
rect 5951 16405 5963 16408
rect 5905 16399 5963 16405
rect 6546 16396 6552 16408
rect 6604 16396 6610 16448
rect 7742 16396 7748 16448
rect 7800 16396 7806 16448
rect 9398 16396 9404 16448
rect 9456 16396 9462 16448
rect 10226 16396 10232 16448
rect 10284 16396 10290 16448
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 11149 16439 11207 16445
rect 11149 16436 11161 16439
rect 11112 16408 11161 16436
rect 11112 16396 11118 16408
rect 11149 16405 11161 16408
rect 11195 16405 11207 16439
rect 11149 16399 11207 16405
rect 11422 16396 11428 16448
rect 11480 16396 11486 16448
rect 14550 16396 14556 16448
rect 14608 16396 14614 16448
rect 18138 16396 18144 16448
rect 18196 16436 18202 16448
rect 19076 16436 19104 16476
rect 19426 16464 19432 16476
rect 19484 16504 19490 16516
rect 19797 16507 19855 16513
rect 19484 16476 19725 16504
rect 19484 16464 19490 16476
rect 18196 16408 19104 16436
rect 18196 16396 18202 16408
rect 19150 16396 19156 16448
rect 19208 16396 19214 16448
rect 19697 16436 19725 16476
rect 19797 16473 19809 16507
rect 19843 16504 19855 16507
rect 19978 16504 19984 16516
rect 19843 16476 19984 16504
rect 19843 16473 19855 16476
rect 19797 16467 19855 16473
rect 19978 16464 19984 16476
rect 20036 16504 20042 16516
rect 20349 16507 20407 16513
rect 20349 16504 20361 16507
rect 20036 16476 20361 16504
rect 20036 16464 20042 16476
rect 20349 16473 20361 16476
rect 20395 16504 20407 16507
rect 20999 16504 21027 16544
rect 26418 16532 26424 16544
rect 26476 16572 26482 16584
rect 26804 16572 26832 16603
rect 26476 16544 26832 16572
rect 26476 16532 26482 16544
rect 20395 16476 21027 16504
rect 21361 16507 21419 16513
rect 20395 16473 20407 16476
rect 20349 16467 20407 16473
rect 21361 16473 21373 16507
rect 21407 16504 21419 16507
rect 21407 16476 21956 16504
rect 21407 16473 21419 16476
rect 21361 16467 21419 16473
rect 20809 16439 20867 16445
rect 20809 16436 20821 16439
rect 19697 16408 20821 16436
rect 20809 16405 20821 16408
rect 20855 16436 20867 16439
rect 21450 16436 21456 16448
rect 20855 16408 21456 16436
rect 20855 16405 20867 16408
rect 20809 16399 20867 16405
rect 21450 16396 21456 16408
rect 21508 16436 21514 16448
rect 21928 16445 21956 16476
rect 26896 16448 26924 16612
rect 27249 16609 27261 16612
rect 27295 16640 27307 16643
rect 27341 16643 27399 16649
rect 27341 16640 27353 16643
rect 27295 16612 27353 16640
rect 27295 16609 27307 16612
rect 27249 16603 27307 16609
rect 27341 16609 27353 16612
rect 27387 16609 27399 16643
rect 27341 16603 27399 16609
rect 27430 16600 27436 16652
rect 27488 16600 27494 16652
rect 27801 16643 27859 16649
rect 27801 16609 27813 16643
rect 27847 16640 27859 16643
rect 28077 16643 28135 16649
rect 28077 16640 28089 16643
rect 27847 16612 28089 16640
rect 27847 16609 27859 16612
rect 27801 16603 27859 16609
rect 28077 16609 28089 16612
rect 28123 16640 28135 16643
rect 28718 16640 28724 16652
rect 28123 16612 28724 16640
rect 28123 16609 28135 16612
rect 28077 16603 28135 16609
rect 28718 16600 28724 16612
rect 28776 16600 28782 16652
rect 29178 16600 29184 16652
rect 29236 16640 29242 16652
rect 29742 16643 29800 16649
rect 29742 16640 29754 16643
rect 29236 16612 29754 16640
rect 29236 16600 29242 16612
rect 29742 16609 29754 16612
rect 29788 16609 29800 16643
rect 29742 16603 29800 16609
rect 27154 16532 27160 16584
rect 27212 16572 27218 16584
rect 27709 16575 27767 16581
rect 27709 16572 27721 16575
rect 27212 16544 27721 16572
rect 27212 16532 27218 16544
rect 27709 16541 27721 16544
rect 27755 16541 27767 16575
rect 27709 16535 27767 16541
rect 30006 16532 30012 16584
rect 30064 16532 30070 16584
rect 21637 16439 21695 16445
rect 21637 16436 21649 16439
rect 21508 16408 21649 16436
rect 21508 16396 21514 16408
rect 21637 16405 21649 16408
rect 21683 16405 21695 16439
rect 21637 16399 21695 16405
rect 21913 16439 21971 16445
rect 21913 16405 21925 16439
rect 21959 16436 21971 16439
rect 22002 16436 22008 16448
rect 21959 16408 22008 16436
rect 21959 16405 21971 16408
rect 21913 16399 21971 16405
rect 22002 16396 22008 16408
rect 22060 16396 22066 16448
rect 24946 16396 24952 16448
rect 25004 16396 25010 16448
rect 26878 16396 26884 16448
rect 26936 16396 26942 16448
rect 28258 16396 28264 16448
rect 28316 16436 28322 16448
rect 28629 16439 28687 16445
rect 28629 16436 28641 16439
rect 28316 16408 28641 16436
rect 28316 16396 28322 16408
rect 28629 16405 28641 16408
rect 28675 16405 28687 16439
rect 28629 16399 28687 16405
rect 552 16346 31372 16368
rect 552 16294 4250 16346
rect 4302 16294 4314 16346
rect 4366 16294 4378 16346
rect 4430 16294 4442 16346
rect 4494 16294 4506 16346
rect 4558 16294 11955 16346
rect 12007 16294 12019 16346
rect 12071 16294 12083 16346
rect 12135 16294 12147 16346
rect 12199 16294 12211 16346
rect 12263 16294 19660 16346
rect 19712 16294 19724 16346
rect 19776 16294 19788 16346
rect 19840 16294 19852 16346
rect 19904 16294 19916 16346
rect 19968 16294 27365 16346
rect 27417 16294 27429 16346
rect 27481 16294 27493 16346
rect 27545 16294 27557 16346
rect 27609 16294 27621 16346
rect 27673 16294 31372 16346
rect 552 16272 31372 16294
rect 1857 16235 1915 16241
rect 1857 16201 1869 16235
rect 1903 16232 1915 16235
rect 1946 16232 1952 16244
rect 1903 16204 1952 16232
rect 1903 16201 1915 16204
rect 1857 16195 1915 16201
rect 1673 16031 1731 16037
rect 1673 15997 1685 16031
rect 1719 16028 1731 16031
rect 1872 16028 1900 16195
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 11054 16192 11060 16244
rect 11112 16192 11118 16244
rect 11422 16192 11428 16244
rect 11480 16192 11486 16244
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 14826 16232 14832 16244
rect 11664 16204 14832 16232
rect 11664 16192 11670 16204
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 19337 16235 19395 16241
rect 19337 16232 19349 16235
rect 19076 16204 19349 16232
rect 2406 16124 2412 16176
rect 2464 16164 2470 16176
rect 9769 16167 9827 16173
rect 2464 16136 3464 16164
rect 2464 16124 2470 16136
rect 2056 16068 3372 16096
rect 2056 16037 2084 16068
rect 1719 16000 1900 16028
rect 1949 16031 2007 16037
rect 1719 15997 1731 16000
rect 1673 15991 1731 15997
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1995 16000 2053 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 2501 16031 2559 16037
rect 2501 16028 2513 16031
rect 2179 16000 2513 16028
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 2501 15997 2513 16000
rect 2547 16028 2559 16031
rect 2777 16031 2835 16037
rect 2777 16028 2789 16031
rect 2547 16000 2789 16028
rect 2547 15997 2559 16000
rect 2501 15991 2559 15997
rect 2777 15997 2789 16000
rect 2823 16028 2835 16031
rect 2961 16031 3019 16037
rect 2961 16028 2973 16031
rect 2823 16000 2973 16028
rect 2823 15997 2835 16000
rect 2777 15991 2835 15997
rect 2961 15997 2973 16000
rect 3007 15997 3019 16031
rect 2961 15991 3019 15997
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 16028 3111 16031
rect 3234 16028 3240 16040
rect 3099 16000 3240 16028
rect 3099 15997 3111 16000
rect 3053 15991 3111 15997
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 1627 15932 2728 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 2700 15904 2728 15932
rect 1486 15852 1492 15904
rect 1544 15892 1550 15904
rect 2406 15892 2412 15904
rect 1544 15864 2412 15892
rect 1544 15852 1550 15864
rect 2406 15852 2412 15864
rect 2464 15852 2470 15904
rect 2682 15852 2688 15904
rect 2740 15852 2746 15904
rect 3344 15892 3372 16068
rect 3436 15969 3464 16136
rect 9769 16133 9781 16167
rect 9815 16164 9827 16167
rect 10870 16164 10876 16176
rect 9815 16136 10876 16164
rect 9815 16133 9827 16136
rect 9769 16127 9827 16133
rect 10870 16124 10876 16136
rect 10928 16124 10934 16176
rect 11072 16164 11100 16192
rect 11072 16136 11744 16164
rect 8386 16056 8392 16108
rect 8444 16056 8450 16108
rect 10134 16096 10140 16108
rect 9876 16068 10140 16096
rect 3510 15988 3516 16040
rect 3568 16028 3574 16040
rect 3605 16031 3663 16037
rect 3605 16028 3617 16031
rect 3568 16000 3617 16028
rect 3568 15988 3574 16000
rect 3605 15997 3617 16000
rect 3651 15997 3663 16031
rect 3605 15991 3663 15997
rect 4985 16031 5043 16037
rect 4985 15997 4997 16031
rect 5031 16028 5043 16031
rect 5626 16028 5632 16040
rect 5031 16000 5632 16028
rect 5031 15997 5043 16000
rect 4985 15991 5043 15997
rect 5626 15988 5632 16000
rect 5684 16028 5690 16040
rect 6454 16028 6460 16040
rect 5684 16000 6460 16028
rect 5684 15988 5690 16000
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 8478 15988 8484 16040
rect 8536 16028 8542 16040
rect 9876 16037 9904 16068
rect 10134 16056 10140 16068
rect 10192 16056 10198 16108
rect 10226 16056 10232 16108
rect 10284 16096 10290 16108
rect 10284 16068 11560 16096
rect 10284 16056 10290 16068
rect 8645 16031 8703 16037
rect 8645 16028 8657 16031
rect 8536 16000 8657 16028
rect 8536 15988 8542 16000
rect 8645 15997 8657 16000
rect 8691 15997 8703 16031
rect 8645 15991 8703 15997
rect 9861 16031 9919 16037
rect 9861 15997 9873 16031
rect 9907 15997 9919 16031
rect 9861 15991 9919 15997
rect 10321 16031 10379 16037
rect 10321 15997 10333 16031
rect 10367 16028 10379 16031
rect 10597 16031 10655 16037
rect 10367 16000 10548 16028
rect 10367 15997 10379 16000
rect 10321 15991 10379 15997
rect 10520 15969 10548 16000
rect 10597 15997 10609 16031
rect 10643 16028 10655 16031
rect 10686 16028 10692 16040
rect 10643 16000 10692 16028
rect 10643 15997 10655 16000
rect 10597 15991 10655 15997
rect 10686 15988 10692 16000
rect 10744 15988 10750 16040
rect 10888 16037 10916 16068
rect 11532 16037 11560 16068
rect 10873 16031 10931 16037
rect 10873 15997 10885 16031
rect 10919 15997 10931 16031
rect 10873 15991 10931 15997
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 11517 16031 11575 16037
rect 11517 15997 11529 16031
rect 11563 15997 11575 16031
rect 11517 15991 11575 15997
rect 3421 15963 3479 15969
rect 3421 15929 3433 15963
rect 3467 15960 3479 15963
rect 5230 15963 5288 15969
rect 5230 15960 5242 15963
rect 3467 15932 5242 15960
rect 3467 15929 3479 15932
rect 3421 15923 3479 15929
rect 5230 15929 5242 15932
rect 5276 15929 5288 15963
rect 5230 15923 5288 15929
rect 10505 15963 10563 15969
rect 10505 15929 10517 15963
rect 10551 15960 10563 15963
rect 10781 15963 10839 15969
rect 10781 15960 10793 15963
rect 10551 15932 10793 15960
rect 10551 15929 10563 15932
rect 10505 15923 10563 15929
rect 10781 15929 10793 15932
rect 10827 15960 10839 15963
rect 10980 15960 11008 15991
rect 10827 15932 11008 15960
rect 11716 15960 11744 16136
rect 17497 16099 17555 16105
rect 17497 16065 17509 16099
rect 17543 16096 17555 16099
rect 17862 16096 17868 16108
rect 17543 16068 17868 16096
rect 17543 16065 17555 16068
rect 17497 16059 17555 16065
rect 17862 16056 17868 16068
rect 17920 16056 17926 16108
rect 19076 16096 19104 16204
rect 19337 16201 19349 16204
rect 19383 16232 19395 16235
rect 19613 16235 19671 16241
rect 19613 16232 19625 16235
rect 19383 16204 19625 16232
rect 19383 16201 19395 16204
rect 19337 16195 19395 16201
rect 19613 16201 19625 16204
rect 19659 16201 19671 16235
rect 19613 16195 19671 16201
rect 20530 16192 20536 16244
rect 20588 16232 20594 16244
rect 20588 16204 21312 16232
rect 20588 16192 20594 16204
rect 19978 16124 19984 16176
rect 20036 16124 20042 16176
rect 20073 16167 20131 16173
rect 20073 16133 20085 16167
rect 20119 16164 20131 16167
rect 20349 16167 20407 16173
rect 20349 16164 20361 16167
rect 20119 16136 20361 16164
rect 20119 16133 20131 16136
rect 20073 16127 20131 16133
rect 20349 16133 20361 16136
rect 20395 16164 20407 16167
rect 20714 16164 20720 16176
rect 20395 16136 20720 16164
rect 20395 16133 20407 16136
rect 20349 16127 20407 16133
rect 20714 16124 20720 16136
rect 20772 16164 20778 16176
rect 20772 16136 20860 16164
rect 20772 16124 20778 16136
rect 18892 16068 19104 16096
rect 11882 15988 11888 16040
rect 11940 16028 11946 16040
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 11940 16000 11989 16028
rect 11940 15988 11946 16000
rect 11977 15997 11989 16000
rect 12023 16028 12035 16031
rect 12618 16028 12624 16040
rect 12023 16000 12624 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12618 15988 12624 16000
rect 12676 16028 12682 16040
rect 14645 16031 14703 16037
rect 14645 16028 14657 16031
rect 12676 16000 14657 16028
rect 12676 15988 12682 16000
rect 14645 15997 14657 16000
rect 14691 15997 14703 16031
rect 14645 15991 14703 15997
rect 17241 16031 17299 16037
rect 17241 15997 17253 16031
rect 17287 16028 17299 16031
rect 18138 16028 18144 16040
rect 17287 16000 18144 16028
rect 17287 15997 17299 16000
rect 17241 15991 17299 15997
rect 18138 15988 18144 16000
rect 18196 15988 18202 16040
rect 18892 16037 18920 16068
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 18340 16000 18889 16028
rect 12222 15963 12280 15969
rect 12222 15960 12234 15963
rect 11716 15932 12234 15960
rect 10827 15929 10839 15932
rect 10781 15923 10839 15929
rect 12222 15929 12234 15932
rect 12268 15960 12280 15963
rect 12342 15960 12348 15972
rect 12268 15932 12348 15960
rect 12268 15929 12280 15932
rect 12222 15923 12280 15929
rect 12342 15920 12348 15932
rect 12400 15920 12406 15972
rect 14912 15963 14970 15969
rect 14912 15929 14924 15963
rect 14958 15960 14970 15963
rect 15470 15960 15476 15972
rect 14958 15932 15476 15960
rect 14958 15929 14970 15932
rect 14912 15923 14970 15929
rect 15470 15920 15476 15932
rect 15528 15920 15534 15972
rect 18340 15904 18368 16000
rect 18877 15997 18889 16000
rect 18923 15997 18935 16031
rect 18877 15991 18935 15997
rect 19153 16031 19211 16037
rect 19153 15997 19165 16031
rect 19199 15997 19211 16031
rect 19153 15991 19211 15997
rect 3697 15895 3755 15901
rect 3697 15892 3709 15895
rect 3344 15864 3709 15892
rect 3697 15861 3709 15864
rect 3743 15892 3755 15895
rect 4154 15892 4160 15904
rect 3743 15864 4160 15892
rect 3743 15861 3755 15864
rect 3697 15855 3755 15861
rect 4154 15852 4160 15864
rect 4212 15852 4218 15904
rect 6362 15852 6368 15904
rect 6420 15852 6426 15904
rect 9953 15895 10011 15901
rect 9953 15861 9965 15895
rect 9999 15892 10011 15895
rect 10229 15895 10287 15901
rect 10229 15892 10241 15895
rect 9999 15864 10241 15892
rect 9999 15861 10011 15864
rect 9953 15855 10011 15861
rect 10229 15861 10241 15864
rect 10275 15892 10287 15895
rect 11790 15892 11796 15904
rect 10275 15864 11796 15892
rect 10275 15861 10287 15864
rect 10229 15855 10287 15861
rect 11790 15852 11796 15864
rect 11848 15852 11854 15904
rect 13357 15895 13415 15901
rect 13357 15861 13369 15895
rect 13403 15892 13415 15895
rect 13446 15892 13452 15904
rect 13403 15864 13452 15892
rect 13403 15861 13415 15864
rect 13357 15855 13415 15861
rect 13446 15852 13452 15864
rect 13504 15852 13510 15904
rect 16022 15852 16028 15904
rect 16080 15852 16086 15904
rect 16117 15895 16175 15901
rect 16117 15861 16129 15895
rect 16163 15892 16175 15895
rect 16482 15892 16488 15904
rect 16163 15864 16488 15892
rect 16163 15861 16175 15864
rect 16117 15855 16175 15861
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 18322 15852 18328 15904
rect 18380 15852 18386 15904
rect 18506 15852 18512 15904
rect 18564 15892 18570 15904
rect 18785 15895 18843 15901
rect 18785 15892 18797 15895
rect 18564 15864 18797 15892
rect 18564 15852 18570 15864
rect 18785 15861 18797 15864
rect 18831 15861 18843 15895
rect 18785 15855 18843 15861
rect 19058 15852 19064 15904
rect 19116 15852 19122 15904
rect 19168 15892 19196 15991
rect 19426 15988 19432 16040
rect 19484 16037 19490 16040
rect 19996 16037 20024 16124
rect 19484 16028 19495 16037
rect 19713 16031 19771 16037
rect 19484 16000 19529 16028
rect 19484 15991 19495 16000
rect 19713 15997 19725 16031
rect 19759 15997 19771 16031
rect 19713 15991 19771 15997
rect 19981 16031 20039 16037
rect 19981 15997 19993 16031
rect 20027 15997 20039 16031
rect 19981 15991 20039 15997
rect 20441 16031 20499 16037
rect 20441 15997 20453 16031
rect 20487 16028 20499 16031
rect 20530 16028 20536 16040
rect 20487 16000 20536 16028
rect 20487 15997 20499 16000
rect 20441 15991 20499 15997
rect 19484 15988 19490 15991
rect 19728 15960 19756 15991
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 20832 16037 20860 16136
rect 21284 16096 21312 16204
rect 26878 16192 26884 16244
rect 26936 16192 26942 16244
rect 27617 16235 27675 16241
rect 27617 16201 27629 16235
rect 27663 16232 27675 16235
rect 28718 16232 28724 16244
rect 27663 16204 28724 16232
rect 27663 16201 27675 16204
rect 27617 16195 27675 16201
rect 28718 16192 28724 16204
rect 28776 16192 28782 16244
rect 29089 16235 29147 16241
rect 29089 16201 29101 16235
rect 29135 16232 29147 16235
rect 29178 16232 29184 16244
rect 29135 16204 29184 16232
rect 29135 16201 29147 16204
rect 29089 16195 29147 16201
rect 23477 16167 23535 16173
rect 23477 16133 23489 16167
rect 23523 16164 23535 16167
rect 23934 16164 23940 16176
rect 23523 16136 23940 16164
rect 23523 16133 23535 16136
rect 23477 16127 23535 16133
rect 23934 16124 23940 16136
rect 23992 16124 23998 16176
rect 29104 16164 29132 16195
rect 29178 16192 29184 16204
rect 29236 16192 29242 16244
rect 28828 16136 29132 16164
rect 22002 16096 22008 16108
rect 21284 16068 22008 16096
rect 21284 16037 21312 16068
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 26697 16099 26755 16105
rect 26697 16065 26709 16099
rect 26743 16096 26755 16099
rect 27062 16096 27068 16108
rect 26743 16068 27068 16096
rect 26743 16065 26755 16068
rect 26697 16059 26755 16065
rect 20717 16031 20775 16037
rect 20717 15997 20729 16031
rect 20763 15997 20775 16031
rect 20717 15991 20775 15997
rect 20809 16031 20867 16037
rect 20809 15997 20821 16031
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 21269 16031 21327 16037
rect 21269 15997 21281 16031
rect 21315 15997 21327 16031
rect 21269 15991 21327 15997
rect 20732 15960 20760 15991
rect 21450 15988 21456 16040
rect 21508 16028 21514 16040
rect 21545 16031 21603 16037
rect 21545 16028 21557 16031
rect 21508 16000 21557 16028
rect 21508 15988 21514 16000
rect 21545 15997 21557 16000
rect 21591 15997 21603 16031
rect 21545 15991 21603 15997
rect 21910 15988 21916 16040
rect 21968 16028 21974 16040
rect 22370 16037 22376 16040
rect 22097 16031 22155 16037
rect 22097 16028 22109 16031
rect 21968 16000 22109 16028
rect 21968 15988 21974 16000
rect 22097 15997 22109 16000
rect 22143 15997 22155 16031
rect 22097 15991 22155 15997
rect 22364 15991 22376 16037
rect 22370 15988 22376 15991
rect 22428 15988 22434 16040
rect 23658 15988 23664 16040
rect 23716 16028 23722 16040
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 23716 16000 25237 16028
rect 23716 15988 23722 16000
rect 25225 15997 25237 16000
rect 25271 16028 25283 16031
rect 26712 16028 26740 16059
rect 27062 16056 27068 16068
rect 27120 16056 27126 16108
rect 25271 16000 26740 16028
rect 26973 16031 27031 16037
rect 25271 15997 25283 16000
rect 25225 15991 25283 15997
rect 26973 15997 26985 16031
rect 27019 16028 27031 16031
rect 27522 16028 27528 16040
rect 27019 16000 27528 16028
rect 27019 15997 27031 16000
rect 26973 15991 27031 15997
rect 27522 15988 27528 16000
rect 27580 15988 27586 16040
rect 28828 16037 28856 16136
rect 29365 16099 29423 16105
rect 29365 16096 29377 16099
rect 28966 16068 29377 16096
rect 27985 16031 28043 16037
rect 27985 15997 27997 16031
rect 28031 16028 28043 16031
rect 28261 16031 28319 16037
rect 28261 16028 28273 16031
rect 28031 16000 28273 16028
rect 28031 15997 28043 16000
rect 27985 15991 28043 15997
rect 28261 15997 28273 16000
rect 28307 16028 28319 16031
rect 28537 16031 28595 16037
rect 28307 16000 28488 16028
rect 28307 15997 28319 16000
rect 28261 15991 28319 15997
rect 20990 15960 20996 15972
rect 19728 15932 20024 15960
rect 20732 15932 20996 15960
rect 19996 15904 20024 15932
rect 20990 15920 20996 15932
rect 21048 15960 21054 15972
rect 24980 15963 25038 15969
rect 21048 15932 21220 15960
rect 21048 15920 21054 15932
rect 19242 15892 19248 15904
rect 19168 15864 19248 15892
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 19978 15852 19984 15904
rect 20036 15892 20042 15904
rect 21192 15901 21220 15932
rect 24980 15929 24992 15963
rect 25026 15960 25038 15963
rect 25406 15960 25412 15972
rect 25026 15932 25412 15960
rect 25026 15929 25038 15932
rect 24980 15923 25038 15929
rect 25406 15920 25412 15932
rect 25464 15920 25470 15972
rect 26418 15920 26424 15972
rect 26476 15969 26482 15972
rect 26476 15960 26488 15969
rect 27540 15960 27568 15988
rect 28169 15963 28227 15969
rect 28169 15960 28181 15963
rect 26476 15932 27200 15960
rect 27540 15932 28181 15960
rect 26476 15923 26488 15932
rect 26476 15920 26482 15923
rect 20625 15895 20683 15901
rect 20625 15892 20637 15895
rect 20036 15864 20637 15892
rect 20036 15852 20042 15864
rect 20625 15861 20637 15864
rect 20671 15892 20683 15895
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20671 15864 20913 15892
rect 20671 15861 20683 15864
rect 20625 15855 20683 15861
rect 20901 15861 20913 15864
rect 20947 15861 20959 15895
rect 20901 15855 20959 15861
rect 21177 15895 21235 15901
rect 21177 15861 21189 15895
rect 21223 15892 21235 15895
rect 21453 15895 21511 15901
rect 21453 15892 21465 15895
rect 21223 15864 21465 15892
rect 21223 15861 21235 15864
rect 21177 15855 21235 15861
rect 21453 15861 21465 15864
rect 21499 15861 21511 15895
rect 21453 15855 21511 15861
rect 23842 15852 23848 15904
rect 23900 15852 23906 15904
rect 24762 15852 24768 15904
rect 24820 15892 24826 15904
rect 25317 15895 25375 15901
rect 25317 15892 25329 15895
rect 24820 15864 25329 15892
rect 24820 15852 24826 15864
rect 25317 15861 25329 15864
rect 25363 15861 25375 15895
rect 27172 15892 27200 15932
rect 28169 15929 28181 15932
rect 28215 15929 28227 15963
rect 28169 15923 28227 15929
rect 28460 15904 28488 16000
rect 28537 15997 28549 16031
rect 28583 16028 28595 16031
rect 28813 16031 28871 16037
rect 28813 16028 28825 16031
rect 28583 16000 28825 16028
rect 28583 15997 28595 16000
rect 28537 15991 28595 15997
rect 28813 15997 28825 16000
rect 28859 15997 28871 16031
rect 28813 15991 28871 15997
rect 28966 15972 28994 16068
rect 29365 16065 29377 16068
rect 29411 16065 29423 16099
rect 29365 16059 29423 16065
rect 29181 16031 29239 16037
rect 29181 15997 29193 16031
rect 29227 16028 29239 16031
rect 29457 16031 29515 16037
rect 29457 16028 29469 16031
rect 29227 16000 29469 16028
rect 29227 15997 29239 16000
rect 29181 15991 29239 15997
rect 28966 15960 29000 15972
rect 28644 15932 29000 15960
rect 28644 15904 28672 15932
rect 28994 15920 29000 15932
rect 29052 15920 29058 15972
rect 29288 15904 29316 16000
rect 29457 15997 29469 16000
rect 29503 15997 29515 16031
rect 29457 15991 29515 15997
rect 27893 15895 27951 15901
rect 27893 15892 27905 15895
rect 27172 15864 27905 15892
rect 25317 15855 25375 15861
rect 27893 15861 27905 15864
rect 27939 15861 27951 15895
rect 27893 15855 27951 15861
rect 28442 15852 28448 15904
rect 28500 15852 28506 15904
rect 28626 15852 28632 15904
rect 28684 15852 28690 15904
rect 29270 15852 29276 15904
rect 29328 15852 29334 15904
rect 552 15802 31531 15824
rect 552 15750 8102 15802
rect 8154 15750 8166 15802
rect 8218 15750 8230 15802
rect 8282 15750 8294 15802
rect 8346 15750 8358 15802
rect 8410 15750 15807 15802
rect 15859 15750 15871 15802
rect 15923 15750 15935 15802
rect 15987 15750 15999 15802
rect 16051 15750 16063 15802
rect 16115 15750 23512 15802
rect 23564 15750 23576 15802
rect 23628 15750 23640 15802
rect 23692 15750 23704 15802
rect 23756 15750 23768 15802
rect 23820 15750 31217 15802
rect 31269 15750 31281 15802
rect 31333 15750 31345 15802
rect 31397 15750 31409 15802
rect 31461 15750 31473 15802
rect 31525 15750 31531 15802
rect 552 15728 31531 15750
rect 1946 15648 1952 15700
rect 2004 15648 2010 15700
rect 2682 15648 2688 15700
rect 2740 15648 2746 15700
rect 9217 15691 9275 15697
rect 9217 15657 9229 15691
rect 9263 15688 9275 15691
rect 10045 15691 10103 15697
rect 10045 15688 10057 15691
rect 9263 15660 10057 15688
rect 9263 15657 9275 15660
rect 9217 15651 9275 15657
rect 10045 15657 10057 15660
rect 10091 15688 10103 15691
rect 10134 15688 10140 15700
rect 10091 15660 10140 15688
rect 10091 15657 10103 15660
rect 10045 15651 10103 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 10226 15648 10232 15700
rect 10284 15688 10290 15700
rect 10597 15691 10655 15697
rect 10597 15688 10609 15691
rect 10284 15660 10609 15688
rect 10284 15648 10290 15660
rect 10597 15657 10609 15660
rect 10643 15657 10655 15691
rect 10597 15651 10655 15657
rect 1305 15555 1363 15561
rect 1305 15521 1317 15555
rect 1351 15552 1363 15555
rect 1486 15552 1492 15564
rect 1351 15524 1492 15552
rect 1351 15521 1363 15524
rect 1305 15515 1363 15521
rect 1486 15512 1492 15524
rect 1544 15512 1550 15564
rect 1964 15561 1992 15648
rect 2700 15620 2728 15648
rect 2930 15623 2988 15629
rect 2930 15620 2942 15623
rect 2148 15592 2942 15620
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15552 1639 15555
rect 1857 15555 1915 15561
rect 1857 15552 1869 15555
rect 1627 15524 1869 15552
rect 1627 15521 1639 15524
rect 1581 15515 1639 15521
rect 1857 15521 1869 15524
rect 1903 15521 1915 15555
rect 1857 15515 1915 15521
rect 1949 15555 2007 15561
rect 1949 15521 1961 15555
rect 1995 15521 2007 15555
rect 1949 15515 2007 15521
rect 1872 15484 1900 15515
rect 2148 15484 2176 15592
rect 2930 15589 2942 15592
rect 2976 15589 2988 15623
rect 2930 15583 2988 15589
rect 4172 15592 6500 15620
rect 4172 15561 4200 15592
rect 6472 15564 6500 15592
rect 6546 15580 6552 15632
rect 6604 15620 6610 15632
rect 6702 15623 6760 15629
rect 6702 15620 6714 15623
rect 6604 15592 6714 15620
rect 6604 15580 6610 15592
rect 6702 15589 6714 15592
rect 6748 15589 6760 15623
rect 6702 15583 6760 15589
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15521 2283 15555
rect 2225 15515 2283 15521
rect 4157 15555 4215 15561
rect 4157 15521 4169 15555
rect 4203 15521 4215 15555
rect 4157 15515 4215 15521
rect 1872 15456 2176 15484
rect 2130 15416 2136 15428
rect 1504 15388 2136 15416
rect 1504 15357 1532 15388
rect 2130 15376 2136 15388
rect 2188 15416 2194 15428
rect 2240 15416 2268 15515
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 4413 15555 4471 15561
rect 4413 15552 4425 15555
rect 4304 15524 4425 15552
rect 4304 15512 4310 15524
rect 4413 15521 4425 15524
rect 4459 15521 4471 15555
rect 4413 15515 4471 15521
rect 6454 15512 6460 15564
rect 6512 15512 6518 15564
rect 9309 15555 9367 15561
rect 9309 15521 9321 15555
rect 9355 15521 9367 15555
rect 9309 15515 9367 15521
rect 2682 15444 2688 15496
rect 2740 15444 2746 15496
rect 9324 15484 9352 15515
rect 9490 15512 9496 15564
rect 9548 15552 9554 15564
rect 9585 15555 9643 15561
rect 9585 15552 9597 15555
rect 9548 15524 9597 15552
rect 9548 15512 9554 15524
rect 9585 15521 9597 15524
rect 9631 15521 9643 15555
rect 9585 15515 9643 15521
rect 9600 15484 9628 15515
rect 9674 15512 9680 15564
rect 9732 15512 9738 15564
rect 10134 15512 10140 15564
rect 10192 15552 10198 15564
rect 10413 15555 10471 15561
rect 10413 15552 10425 15555
rect 10192 15524 10425 15552
rect 10192 15512 10198 15524
rect 10413 15521 10425 15524
rect 10459 15521 10471 15555
rect 10413 15515 10471 15521
rect 10505 15555 10563 15561
rect 10505 15521 10517 15555
rect 10551 15521 10563 15555
rect 10505 15515 10563 15521
rect 10321 15487 10379 15493
rect 10321 15484 10333 15487
rect 9324 15456 9536 15484
rect 9600 15456 10333 15484
rect 2188 15388 2268 15416
rect 2188 15376 2194 15388
rect 1213 15351 1271 15357
rect 1213 15317 1225 15351
rect 1259 15348 1271 15351
rect 1489 15351 1547 15357
rect 1489 15348 1501 15351
rect 1259 15320 1501 15348
rect 1259 15317 1271 15320
rect 1213 15311 1271 15317
rect 1489 15317 1501 15320
rect 1535 15317 1547 15351
rect 1489 15311 1547 15317
rect 1762 15308 1768 15360
rect 1820 15308 1826 15360
rect 2041 15351 2099 15357
rect 2041 15317 2053 15351
rect 2087 15348 2099 15351
rect 2314 15348 2320 15360
rect 2087 15320 2320 15348
rect 2087 15317 2099 15320
rect 2041 15311 2099 15317
rect 2314 15308 2320 15320
rect 2372 15308 2378 15360
rect 4062 15308 4068 15360
rect 4120 15308 4126 15360
rect 5537 15351 5595 15357
rect 5537 15317 5549 15351
rect 5583 15348 5595 15351
rect 5810 15348 5816 15360
rect 5583 15320 5816 15348
rect 5583 15317 5595 15320
rect 5537 15311 5595 15317
rect 5810 15308 5816 15320
rect 5868 15308 5874 15360
rect 7374 15308 7380 15360
rect 7432 15348 7438 15360
rect 9508 15357 9536 15456
rect 10321 15453 10333 15456
rect 10367 15484 10379 15487
rect 10520 15484 10548 15515
rect 10367 15456 10548 15484
rect 10612 15484 10640 15651
rect 11790 15648 11796 15700
rect 11848 15688 11854 15700
rect 11848 15660 12434 15688
rect 11848 15648 11854 15660
rect 10778 15580 10784 15632
rect 10836 15620 10842 15632
rect 11882 15620 11888 15632
rect 10836 15592 11888 15620
rect 10836 15580 10842 15592
rect 10686 15512 10692 15564
rect 10744 15552 10750 15564
rect 11238 15552 11244 15564
rect 10744 15524 11244 15552
rect 10744 15512 10750 15524
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11532 15561 11560 15592
rect 11882 15580 11888 15592
rect 11940 15580 11946 15632
rect 11517 15555 11575 15561
rect 11517 15521 11529 15555
rect 11563 15521 11575 15555
rect 11773 15555 11831 15561
rect 11773 15552 11785 15555
rect 11517 15515 11575 15521
rect 11624 15524 11785 15552
rect 11624 15484 11652 15524
rect 11773 15521 11785 15524
rect 11819 15521 11831 15555
rect 12406 15552 12434 15660
rect 12618 15648 12624 15700
rect 12676 15648 12682 15700
rect 15470 15648 15476 15700
rect 15528 15648 15534 15700
rect 19058 15648 19064 15700
rect 19116 15648 19122 15700
rect 19242 15648 19248 15700
rect 19300 15688 19306 15700
rect 19978 15688 19984 15700
rect 19300 15660 19984 15688
rect 19300 15648 19306 15660
rect 12636 15620 12664 15648
rect 15488 15620 15516 15648
rect 18506 15620 18512 15632
rect 12636 15592 13676 15620
rect 13648 15561 13676 15592
rect 15488 15592 18512 15620
rect 13633 15555 13691 15561
rect 12406 15524 13216 15552
rect 11773 15515 11831 15521
rect 10612 15456 11652 15484
rect 13188 15484 13216 15524
rect 13633 15521 13645 15555
rect 13679 15521 13691 15555
rect 13889 15555 13947 15561
rect 13889 15552 13901 15555
rect 13633 15515 13691 15521
rect 13740 15524 13901 15552
rect 13740 15484 13768 15524
rect 13889 15521 13901 15524
rect 13935 15521 13947 15555
rect 13889 15515 13947 15521
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15521 15347 15555
rect 15488 15552 15516 15592
rect 17420 15561 17448 15592
rect 18506 15580 18512 15592
rect 18564 15580 18570 15632
rect 15565 15555 15623 15561
rect 15565 15552 15577 15555
rect 15488 15524 15577 15552
rect 15289 15515 15347 15521
rect 15565 15521 15577 15524
rect 15611 15521 15623 15555
rect 15565 15515 15623 15521
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15552 16911 15555
rect 17129 15555 17187 15561
rect 17129 15552 17141 15555
rect 16899 15524 17141 15552
rect 16899 15521 16911 15524
rect 16853 15515 16911 15521
rect 17129 15521 17141 15524
rect 17175 15521 17187 15555
rect 17129 15515 17187 15521
rect 17405 15555 17463 15561
rect 17405 15521 17417 15555
rect 17451 15521 17463 15555
rect 17405 15515 17463 15521
rect 17681 15555 17739 15561
rect 17681 15521 17693 15555
rect 17727 15552 17739 15555
rect 17727 15524 18276 15552
rect 17727 15521 17739 15524
rect 17681 15515 17739 15521
rect 13188 15456 13768 15484
rect 15304 15484 15332 15515
rect 15838 15484 15844 15496
rect 15304 15456 15844 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 17144 15484 17172 15515
rect 18248 15493 18276 15524
rect 18322 15512 18328 15564
rect 18380 15512 18386 15564
rect 18601 15555 18659 15561
rect 18601 15521 18613 15555
rect 18647 15552 18659 15555
rect 18877 15555 18935 15561
rect 18877 15552 18889 15555
rect 18647 15524 18889 15552
rect 18647 15521 18659 15524
rect 18601 15515 18659 15521
rect 18877 15521 18889 15524
rect 18923 15552 18935 15555
rect 19076 15552 19104 15648
rect 19619 15629 19647 15660
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 20990 15648 20996 15700
rect 21048 15648 21054 15700
rect 23842 15648 23848 15700
rect 23900 15648 23906 15700
rect 28169 15691 28227 15697
rect 28169 15688 28181 15691
rect 27724 15660 28181 15688
rect 19604 15623 19662 15629
rect 19604 15589 19616 15623
rect 19650 15589 19662 15623
rect 19604 15583 19662 15589
rect 21008 15561 21036 15648
rect 22002 15580 22008 15632
rect 22060 15620 22066 15632
rect 22158 15623 22216 15629
rect 22158 15620 22170 15623
rect 22060 15592 22170 15620
rect 22060 15580 22066 15592
rect 22158 15589 22170 15592
rect 22204 15589 22216 15623
rect 23860 15620 23888 15648
rect 23860 15592 24624 15620
rect 22158 15583 22216 15589
rect 18923 15524 19104 15552
rect 19153 15555 19211 15561
rect 18923 15521 18935 15524
rect 18877 15515 18935 15521
rect 19153 15521 19165 15555
rect 19199 15552 19211 15555
rect 20993 15555 21051 15561
rect 19199 15524 20944 15552
rect 19199 15521 19211 15524
rect 19153 15515 19211 15521
rect 17313 15487 17371 15493
rect 17313 15484 17325 15487
rect 17144 15456 17325 15484
rect 17313 15453 17325 15456
rect 17359 15484 17371 15487
rect 17589 15487 17647 15493
rect 17589 15484 17601 15487
rect 17359 15456 17601 15484
rect 17359 15453 17371 15456
rect 17313 15447 17371 15453
rect 17589 15453 17601 15456
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 18233 15487 18291 15493
rect 18233 15453 18245 15487
rect 18279 15484 18291 15487
rect 19168 15484 19196 15515
rect 18279 15456 19196 15484
rect 18279 15453 18291 15456
rect 18233 15447 18291 15453
rect 19334 15444 19340 15496
rect 19392 15444 19398 15496
rect 9769 15419 9827 15425
rect 9769 15416 9781 15419
rect 9646 15388 9781 15416
rect 7837 15351 7895 15357
rect 7837 15348 7849 15351
rect 7432 15320 7849 15348
rect 7432 15308 7438 15320
rect 7837 15317 7849 15320
rect 7883 15317 7895 15351
rect 7837 15311 7895 15317
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 9646 15348 9674 15388
rect 9769 15385 9781 15388
rect 9815 15416 9827 15419
rect 10686 15416 10692 15428
rect 9815 15388 10692 15416
rect 9815 15385 9827 15388
rect 9769 15379 9827 15385
rect 10686 15376 10692 15388
rect 10744 15376 10750 15428
rect 14918 15376 14924 15428
rect 14976 15416 14982 15428
rect 14976 15388 15240 15416
rect 14976 15376 14982 15388
rect 9539 15320 9674 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 12894 15308 12900 15360
rect 12952 15308 12958 15360
rect 15013 15351 15071 15357
rect 15013 15317 15025 15351
rect 15059 15348 15071 15351
rect 15102 15348 15108 15360
rect 15059 15320 15108 15348
rect 15059 15317 15071 15320
rect 15013 15311 15071 15317
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 15212 15357 15240 15388
rect 15562 15376 15568 15428
rect 15620 15416 15626 15428
rect 15620 15388 17080 15416
rect 15620 15376 15626 15388
rect 15197 15351 15255 15357
rect 15197 15317 15209 15351
rect 15243 15348 15255 15351
rect 15378 15348 15384 15360
rect 15243 15320 15384 15348
rect 15243 15317 15255 15320
rect 15197 15311 15255 15317
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 15470 15308 15476 15360
rect 15528 15308 15534 15360
rect 16758 15308 16764 15360
rect 16816 15308 16822 15360
rect 17052 15357 17080 15388
rect 20916 15360 20944 15524
rect 20993 15521 21005 15555
rect 21039 15521 21051 15555
rect 20993 15515 21051 15521
rect 21910 15512 21916 15564
rect 21968 15512 21974 15564
rect 24302 15561 24308 15564
rect 24300 15552 24308 15561
rect 24263 15524 24308 15552
rect 24300 15515 24308 15524
rect 24302 15512 24308 15515
rect 24360 15512 24366 15564
rect 24394 15512 24400 15564
rect 24452 15512 24458 15564
rect 24596 15561 24624 15592
rect 27522 15580 27528 15632
rect 27580 15629 27586 15632
rect 27580 15620 27592 15629
rect 27724 15620 27752 15660
rect 28169 15657 28181 15660
rect 28215 15657 28227 15691
rect 28169 15651 28227 15657
rect 28442 15648 28448 15700
rect 28500 15648 28506 15700
rect 28994 15648 29000 15700
rect 29052 15648 29058 15700
rect 30006 15648 30012 15700
rect 30064 15648 30070 15700
rect 27580 15592 27752 15620
rect 29012 15620 29040 15648
rect 30024 15620 30052 15648
rect 29012 15592 29500 15620
rect 27580 15583 27592 15592
rect 27580 15580 27586 15583
rect 24489 15555 24547 15561
rect 24489 15521 24501 15555
rect 24535 15521 24547 15555
rect 24596 15555 24675 15561
rect 24596 15524 24629 15555
rect 24489 15515 24547 15521
rect 24617 15521 24629 15524
rect 24663 15521 24675 15555
rect 24617 15515 24675 15521
rect 24765 15555 24823 15561
rect 24765 15521 24777 15555
rect 24811 15521 24823 15555
rect 24765 15515 24823 15521
rect 24210 15444 24216 15496
rect 24268 15484 24274 15496
rect 24504 15484 24532 15515
rect 24268 15456 24532 15484
rect 24268 15444 24274 15456
rect 24780 15416 24808 15515
rect 25958 15512 25964 15564
rect 26016 15552 26022 15564
rect 27062 15552 27068 15564
rect 26016 15524 27068 15552
rect 26016 15512 26022 15524
rect 27062 15512 27068 15524
rect 27120 15552 27126 15564
rect 28261 15555 28319 15561
rect 27120 15524 27752 15552
rect 27120 15512 27126 15524
rect 27724 15484 27752 15524
rect 28261 15521 28273 15555
rect 28307 15521 28319 15555
rect 28261 15515 28319 15521
rect 28537 15555 28595 15561
rect 28537 15521 28549 15555
rect 28583 15552 28595 15555
rect 28626 15552 28632 15564
rect 28583 15524 28632 15552
rect 28583 15521 28595 15524
rect 28537 15515 28595 15521
rect 27801 15487 27859 15493
rect 27801 15484 27813 15487
rect 27724 15456 27813 15484
rect 27801 15453 27813 15456
rect 27847 15453 27859 15487
rect 28276 15484 28304 15515
rect 28626 15512 28632 15524
rect 28684 15512 28690 15564
rect 29012 15552 29040 15592
rect 29089 15555 29147 15561
rect 29089 15552 29101 15555
rect 28813 15545 28871 15551
rect 28813 15511 28825 15545
rect 28859 15511 28871 15545
rect 29012 15524 29101 15552
rect 29089 15521 29101 15524
rect 29135 15521 29147 15555
rect 29089 15515 29147 15521
rect 29189 15553 29247 15559
rect 29189 15519 29201 15553
rect 29235 15550 29247 15553
rect 29288 15550 29408 15552
rect 29235 15524 29408 15550
rect 29235 15522 29316 15524
rect 29235 15519 29247 15522
rect 29189 15513 29247 15519
rect 28813 15505 28871 15511
rect 28721 15487 28779 15493
rect 28721 15484 28733 15487
rect 28276 15456 28733 15484
rect 27801 15447 27859 15453
rect 28721 15453 28733 15456
rect 28767 15453 28779 15487
rect 28721 15447 28779 15453
rect 23221 15388 24808 15416
rect 17037 15351 17095 15357
rect 17037 15317 17049 15351
rect 17083 15348 17095 15351
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 17083 15320 18797 15348
rect 17083 15317 17095 15320
rect 17037 15311 17095 15317
rect 18785 15317 18797 15320
rect 18831 15348 18843 15351
rect 19058 15348 19064 15360
rect 18831 15320 19064 15348
rect 18831 15317 18843 15320
rect 18785 15311 18843 15317
rect 19058 15308 19064 15320
rect 19116 15308 19122 15360
rect 20714 15308 20720 15360
rect 20772 15308 20778 15360
rect 20898 15308 20904 15360
rect 20956 15308 20962 15360
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 23221 15348 23249 15388
rect 21048 15320 23249 15348
rect 23293 15351 23351 15357
rect 21048 15308 21054 15320
rect 23293 15317 23305 15351
rect 23339 15348 23351 15351
rect 23934 15348 23940 15360
rect 23339 15320 23940 15348
rect 23339 15317 23351 15320
rect 23293 15311 23351 15317
rect 23934 15308 23940 15320
rect 23992 15308 23998 15360
rect 24118 15308 24124 15360
rect 24176 15308 24182 15360
rect 26234 15308 26240 15360
rect 26292 15348 26298 15360
rect 26421 15351 26479 15357
rect 26421 15348 26433 15351
rect 26292 15320 26433 15348
rect 26292 15308 26298 15320
rect 26421 15317 26433 15320
rect 26467 15317 26479 15351
rect 28736 15348 28764 15447
rect 28828 15428 28856 15505
rect 28810 15376 28816 15428
rect 28868 15376 28874 15428
rect 29178 15376 29184 15428
rect 29236 15416 29242 15428
rect 29273 15419 29331 15425
rect 29273 15416 29285 15419
rect 29236 15388 29285 15416
rect 29236 15376 29242 15388
rect 29273 15385 29285 15388
rect 29319 15385 29331 15419
rect 29273 15379 29331 15385
rect 28997 15351 29055 15357
rect 28997 15348 29009 15351
rect 28736 15320 29009 15348
rect 26421 15311 26479 15317
rect 28997 15317 29009 15320
rect 29043 15348 29055 15351
rect 29380 15348 29408 15524
rect 29472 15484 29500 15592
rect 29564 15592 30052 15620
rect 29564 15564 29592 15592
rect 29546 15512 29552 15564
rect 29604 15512 29610 15564
rect 29805 15555 29863 15561
rect 29805 15552 29817 15555
rect 29647 15524 29817 15552
rect 29647 15484 29675 15524
rect 29805 15521 29817 15524
rect 29851 15521 29863 15555
rect 29805 15515 29863 15521
rect 29472 15456 29675 15484
rect 29043 15320 29408 15348
rect 29043 15317 29055 15320
rect 28997 15311 29055 15317
rect 30926 15308 30932 15360
rect 30984 15308 30990 15360
rect 552 15258 31372 15280
rect 552 15206 4250 15258
rect 4302 15206 4314 15258
rect 4366 15206 4378 15258
rect 4430 15206 4442 15258
rect 4494 15206 4506 15258
rect 4558 15206 11955 15258
rect 12007 15206 12019 15258
rect 12071 15206 12083 15258
rect 12135 15206 12147 15258
rect 12199 15206 12211 15258
rect 12263 15206 19660 15258
rect 19712 15206 19724 15258
rect 19776 15206 19788 15258
rect 19840 15206 19852 15258
rect 19904 15206 19916 15258
rect 19968 15206 27365 15258
rect 27417 15206 27429 15258
rect 27481 15206 27493 15258
rect 27545 15206 27557 15258
rect 27609 15206 27621 15258
rect 27673 15206 31372 15258
rect 552 15184 31372 15206
rect 1762 15104 1768 15156
rect 1820 15144 1826 15156
rect 1949 15147 2007 15153
rect 1949 15144 1961 15147
rect 1820 15116 1961 15144
rect 1820 15104 1826 15116
rect 1949 15113 1961 15116
rect 1995 15113 2007 15147
rect 1949 15107 2007 15113
rect 9309 15147 9367 15153
rect 9309 15113 9321 15147
rect 9355 15144 9367 15147
rect 9490 15144 9496 15156
rect 9355 15116 9496 15144
rect 9355 15113 9367 15116
rect 9309 15107 9367 15113
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 13722 15144 13728 15156
rect 11900 15116 13728 15144
rect 1780 14949 1808 15104
rect 8202 15036 8208 15088
rect 8260 15036 8266 15088
rect 11425 15079 11483 15085
rect 11425 15045 11437 15079
rect 11471 15076 11483 15079
rect 11900 15076 11928 15116
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 14737 15147 14795 15153
rect 14737 15144 14749 15147
rect 14200 15116 14749 15144
rect 11471 15048 11928 15076
rect 11471 15045 11483 15048
rect 11425 15039 11483 15045
rect 2056 14980 2360 15008
rect 2056 14949 2084 14980
rect 2332 14952 2360 14980
rect 2682 14968 2688 15020
rect 2740 15008 2746 15020
rect 2740 14980 4660 15008
rect 2740 14968 2746 14980
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14909 1823 14943
rect 1765 14903 1823 14909
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 2130 14900 2136 14952
rect 2188 14900 2194 14952
rect 2314 14900 2320 14952
rect 2372 14900 2378 14952
rect 4632 14949 4660 14980
rect 6454 14968 6460 15020
rect 6512 15008 6518 15020
rect 6825 15011 6883 15017
rect 6825 15008 6837 15011
rect 6512 14980 6837 15008
rect 6512 14968 6518 14980
rect 6825 14977 6837 14980
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 9692 14980 9996 15008
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14940 4675 14943
rect 6472 14940 6500 14968
rect 9692 14949 9720 14980
rect 9968 14952 9996 14980
rect 13078 14968 13084 15020
rect 13136 15008 13142 15020
rect 14200 15008 14228 15116
rect 14737 15113 14749 15116
rect 14783 15144 14795 15147
rect 14783 15116 15240 15144
rect 14783 15113 14795 15116
rect 14737 15107 14795 15113
rect 15212 15076 15240 15116
rect 15378 15104 15384 15156
rect 15436 15144 15442 15156
rect 15565 15147 15623 15153
rect 15565 15144 15577 15147
rect 15436 15116 15577 15144
rect 15436 15104 15442 15116
rect 15565 15113 15577 15116
rect 15611 15113 15623 15147
rect 15565 15107 15623 15113
rect 18782 15104 18788 15156
rect 18840 15104 18846 15156
rect 19245 15147 19303 15153
rect 19245 15113 19257 15147
rect 19291 15144 19303 15147
rect 20990 15144 20996 15156
rect 19291 15116 20996 15144
rect 19291 15113 19303 15116
rect 19245 15107 19303 15113
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 24394 15104 24400 15156
rect 24452 15144 24458 15156
rect 25225 15147 25283 15153
rect 25225 15144 25237 15147
rect 24452 15116 25237 15144
rect 24452 15104 24458 15116
rect 25225 15113 25237 15116
rect 25271 15113 25283 15147
rect 25225 15107 25283 15113
rect 28718 15104 28724 15156
rect 28776 15104 28782 15156
rect 29270 15144 29276 15156
rect 29012 15116 29276 15144
rect 15286 15076 15292 15088
rect 15212 15048 15292 15076
rect 15286 15036 15292 15048
rect 15344 15036 15350 15088
rect 18800 15076 18828 15104
rect 18800 15048 19012 15076
rect 15013 15011 15071 15017
rect 13136 14980 14228 15008
rect 14292 14980 14872 15008
rect 13136 14968 13142 14980
rect 4663 14912 6500 14940
rect 9401 14943 9459 14949
rect 4663 14909 4675 14912
rect 4617 14903 4675 14909
rect 9401 14909 9413 14943
rect 9447 14940 9459 14943
rect 9677 14943 9735 14949
rect 9677 14940 9689 14943
rect 9447 14912 9689 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 9677 14909 9689 14912
rect 9723 14909 9735 14943
rect 9677 14903 9735 14909
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14909 9827 14943
rect 9769 14903 9827 14909
rect 4706 14832 4712 14884
rect 4764 14872 4770 14884
rect 4862 14875 4920 14881
rect 4862 14872 4874 14875
rect 4764 14844 4874 14872
rect 4764 14832 4770 14844
rect 4862 14841 4874 14844
rect 4908 14841 4920 14875
rect 4862 14835 4920 14841
rect 6086 14832 6092 14884
rect 6144 14872 6150 14884
rect 7070 14875 7128 14881
rect 7070 14872 7082 14875
rect 6144 14844 7082 14872
rect 6144 14832 6150 14844
rect 7070 14841 7082 14844
rect 7116 14841 7128 14875
rect 9784 14872 9812 14903
rect 9950 14900 9956 14952
rect 10008 14900 10014 14952
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14940 10103 14943
rect 10778 14940 10784 14952
rect 10091 14912 10784 14940
rect 10091 14909 10103 14912
rect 10045 14903 10103 14909
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 11882 14940 11888 14952
rect 11112 14912 11888 14940
rect 11112 14900 11118 14912
rect 11882 14900 11888 14912
rect 11940 14940 11946 14952
rect 14292 14949 14320 14980
rect 14844 14949 14872 14980
rect 15013 14977 15025 15011
rect 15059 15008 15071 15011
rect 15470 15008 15476 15020
rect 15059 14980 15476 15008
rect 15059 14977 15071 14980
rect 15013 14971 15071 14977
rect 15470 14968 15476 14980
rect 15528 15008 15534 15020
rect 15528 14980 15792 15008
rect 15528 14968 15534 14980
rect 11977 14943 12035 14949
rect 11977 14940 11989 14943
rect 11940 14912 11989 14940
rect 11940 14900 11946 14912
rect 11977 14909 11989 14912
rect 12023 14909 12035 14943
rect 11977 14903 12035 14909
rect 12244 14943 12302 14949
rect 12244 14909 12256 14943
rect 12290 14940 12302 14943
rect 14277 14943 14335 14949
rect 12290 14912 14228 14940
rect 12290 14909 12302 14912
rect 12244 14903 12302 14909
rect 7070 14835 7128 14841
rect 9692 14844 9812 14872
rect 9861 14875 9919 14881
rect 9692 14816 9720 14844
rect 9861 14841 9873 14875
rect 9907 14872 9919 14875
rect 10134 14872 10140 14884
rect 9907 14844 10140 14872
rect 9907 14841 9919 14844
rect 9861 14835 9919 14841
rect 10134 14832 10140 14844
rect 10192 14872 10198 14884
rect 10312 14875 10370 14881
rect 10312 14872 10324 14875
rect 10192 14844 10324 14872
rect 10192 14832 10198 14844
rect 10312 14841 10324 14844
rect 10358 14872 10370 14875
rect 10502 14872 10508 14884
rect 10358 14844 10508 14872
rect 10358 14841 10370 14844
rect 10312 14835 10370 14841
rect 10502 14832 10508 14844
rect 10560 14832 10566 14884
rect 14200 14816 14228 14912
rect 14277 14909 14289 14943
rect 14323 14909 14335 14943
rect 14277 14903 14335 14909
rect 14553 14943 14611 14949
rect 14553 14909 14565 14943
rect 14599 14940 14611 14943
rect 14829 14943 14887 14949
rect 14599 14912 14796 14940
rect 14599 14909 14611 14912
rect 14553 14903 14611 14909
rect 1673 14807 1731 14813
rect 1673 14773 1685 14807
rect 1719 14804 1731 14807
rect 2222 14804 2228 14816
rect 1719 14776 2228 14804
rect 1719 14773 1731 14776
rect 1673 14767 1731 14773
rect 2222 14764 2228 14776
rect 2280 14764 2286 14816
rect 5994 14764 6000 14816
rect 6052 14764 6058 14816
rect 9585 14807 9643 14813
rect 9585 14773 9597 14807
rect 9631 14804 9643 14807
rect 9674 14804 9680 14816
rect 9631 14776 9680 14804
rect 9631 14773 9643 14776
rect 9585 14767 9643 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 13357 14807 13415 14813
rect 13357 14773 13369 14807
rect 13403 14804 13415 14807
rect 13630 14804 13636 14816
rect 13403 14776 13636 14804
rect 13403 14773 13415 14776
rect 13357 14767 13415 14773
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 14182 14764 14188 14816
rect 14240 14764 14246 14816
rect 14458 14764 14464 14816
rect 14516 14764 14522 14816
rect 14768 14804 14796 14912
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 14918 14940 14924 14952
rect 14875 14912 14924 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 14918 14900 14924 14912
rect 14976 14900 14982 14952
rect 15105 14943 15163 14949
rect 15105 14909 15117 14943
rect 15151 14909 15163 14943
rect 15105 14903 15163 14909
rect 15381 14943 15439 14949
rect 15381 14909 15393 14943
rect 15427 14940 15439 14943
rect 15488 14940 15516 14968
rect 15764 14949 15792 14980
rect 16206 14968 16212 15020
rect 16264 14968 16270 15020
rect 17880 14980 18920 15008
rect 17880 14952 17908 14980
rect 15427 14912 15516 14940
rect 15657 14943 15715 14949
rect 15427 14909 15439 14912
rect 15381 14903 15439 14909
rect 15657 14909 15669 14943
rect 15703 14909 15715 14943
rect 15657 14903 15715 14909
rect 15749 14943 15807 14949
rect 15749 14909 15761 14943
rect 15795 14909 15807 14943
rect 15749 14903 15807 14909
rect 15120 14872 15148 14903
rect 15562 14872 15568 14884
rect 15120 14844 15568 14872
rect 15562 14832 15568 14844
rect 15620 14872 15626 14884
rect 15672 14872 15700 14903
rect 15838 14900 15844 14952
rect 15896 14940 15902 14952
rect 16476 14943 16534 14949
rect 16476 14940 16488 14943
rect 15896 14912 16488 14940
rect 15896 14900 15902 14912
rect 16476 14909 16488 14912
rect 16522 14940 16534 14943
rect 16758 14940 16764 14952
rect 16522 14912 16764 14940
rect 16522 14909 16534 14912
rect 16476 14903 16534 14909
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 17678 14900 17684 14952
rect 17736 14900 17742 14952
rect 17862 14900 17868 14952
rect 17920 14900 17926 14952
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 15620 14844 15700 14872
rect 15620 14832 15626 14844
rect 15856 14804 15884 14900
rect 17957 14875 18015 14881
rect 17957 14841 17969 14875
rect 18003 14841 18015 14875
rect 18064 14872 18092 14903
rect 18690 14900 18696 14952
rect 18748 14900 18754 14952
rect 18892 14949 18920 14980
rect 18984 14949 19012 15048
rect 19058 15036 19064 15088
rect 19116 15076 19122 15088
rect 19794 15076 19800 15088
rect 19116 15048 19800 15076
rect 19116 15036 19122 15048
rect 19794 15036 19800 15048
rect 19852 15036 19858 15088
rect 22738 15036 22744 15088
rect 22796 15076 22802 15088
rect 24489 15079 24547 15085
rect 24489 15076 24501 15079
rect 22796 15048 24501 15076
rect 22796 15036 22802 15048
rect 24489 15045 24501 15048
rect 24535 15045 24547 15079
rect 24489 15039 24547 15045
rect 28445 15079 28503 15085
rect 28445 15045 28457 15079
rect 28491 15076 28503 15079
rect 29012 15076 29040 15116
rect 29270 15104 29276 15116
rect 29328 15144 29334 15156
rect 29917 15147 29975 15153
rect 29917 15144 29929 15147
rect 29328 15116 29929 15144
rect 29328 15104 29334 15116
rect 29917 15113 29929 15116
rect 29963 15113 29975 15147
rect 29917 15107 29975 15113
rect 28491 15048 29040 15076
rect 29089 15079 29147 15085
rect 28491 15045 28503 15048
rect 28445 15039 28503 15045
rect 29089 15045 29101 15079
rect 29135 15076 29147 15079
rect 29638 15076 29644 15088
rect 29135 15048 29644 15076
rect 29135 15045 29147 15048
rect 29089 15039 29147 15045
rect 20530 15008 20536 15020
rect 19352 14980 20536 15008
rect 19352 14952 19380 14980
rect 20530 14968 20536 14980
rect 20588 15008 20594 15020
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20588 14980 20729 15008
rect 20588 14968 20594 14980
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 23290 14968 23296 15020
rect 23348 15008 23354 15020
rect 28718 15008 28724 15020
rect 23348 14980 24164 15008
rect 23348 14968 23354 14980
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14909 19027 14943
rect 18969 14903 19027 14909
rect 19058 14900 19064 14952
rect 19116 14940 19122 14952
rect 19116 14912 19288 14940
rect 19116 14900 19122 14912
rect 19260 14872 19288 14912
rect 19334 14900 19340 14952
rect 19392 14900 19398 14952
rect 20990 14949 20996 14952
rect 20984 14903 20996 14949
rect 20990 14900 20996 14903
rect 21048 14900 21054 14952
rect 23845 14943 23903 14949
rect 23845 14909 23857 14943
rect 23891 14909 23903 14943
rect 23845 14903 23903 14909
rect 21174 14872 21180 14884
rect 18064 14844 18828 14872
rect 19260 14844 21180 14872
rect 17957 14835 18015 14841
rect 14768 14776 15884 14804
rect 17589 14807 17647 14813
rect 17589 14773 17601 14807
rect 17635 14804 17647 14807
rect 17972 14804 18000 14835
rect 17635 14776 18000 14804
rect 17635 14773 17647 14776
rect 17589 14767 17647 14773
rect 18230 14764 18236 14816
rect 18288 14764 18294 14816
rect 18800 14804 18828 14844
rect 21174 14832 21180 14844
rect 21232 14832 21238 14884
rect 21358 14804 21364 14816
rect 18800 14776 21364 14804
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 22094 14764 22100 14816
rect 22152 14764 22158 14816
rect 23860 14804 23888 14903
rect 23934 14900 23940 14952
rect 23992 14940 23998 14952
rect 24136 14949 24164 14980
rect 28552 14980 28724 15008
rect 24121 14943 24179 14949
rect 23992 14912 24037 14940
rect 23992 14900 23998 14912
rect 24121 14909 24133 14943
rect 24167 14909 24179 14943
rect 24121 14903 24179 14909
rect 24302 14900 24308 14952
rect 24360 14949 24366 14952
rect 24360 14943 24409 14949
rect 24360 14909 24363 14943
rect 24397 14940 24409 14943
rect 24578 14940 24584 14952
rect 24397 14912 24584 14940
rect 24397 14909 24409 14912
rect 24360 14903 24409 14909
rect 24360 14900 24366 14903
rect 24578 14900 24584 14912
rect 24636 14900 24642 14952
rect 25958 14900 25964 14952
rect 26016 14940 26022 14952
rect 28552 14949 28580 14980
rect 28718 14968 28724 14980
rect 28776 15008 28782 15020
rect 29104 15008 29132 15039
rect 29638 15036 29644 15048
rect 29696 15036 29702 15088
rect 28776 14980 29132 15008
rect 29472 14980 29868 15008
rect 28776 14968 28782 14980
rect 29472 14952 29500 14980
rect 26605 14943 26663 14949
rect 26605 14940 26617 14943
rect 26016 14912 26617 14940
rect 26016 14900 26022 14912
rect 26605 14909 26617 14912
rect 26651 14909 26663 14943
rect 26605 14903 26663 14909
rect 28537 14943 28595 14949
rect 28537 14909 28549 14943
rect 28583 14909 28595 14943
rect 28537 14903 28595 14909
rect 28813 14943 28871 14949
rect 28813 14909 28825 14943
rect 28859 14909 28871 14943
rect 28813 14903 28871 14909
rect 24213 14875 24271 14881
rect 24213 14841 24225 14875
rect 24259 14872 24271 14875
rect 26234 14872 26240 14884
rect 24259 14844 26240 14872
rect 24259 14841 24271 14844
rect 24213 14835 24271 14841
rect 26234 14832 26240 14844
rect 26292 14832 26298 14884
rect 26360 14875 26418 14881
rect 26360 14841 26372 14875
rect 26406 14872 26418 14875
rect 26786 14872 26792 14884
rect 26406 14844 26792 14872
rect 26406 14841 26418 14844
rect 26360 14835 26418 14841
rect 26786 14832 26792 14844
rect 26844 14832 26850 14884
rect 28828 14872 28856 14903
rect 29178 14900 29184 14952
rect 29236 14900 29242 14952
rect 29454 14900 29460 14952
rect 29512 14900 29518 14952
rect 29840 14949 29868 14980
rect 29549 14943 29607 14949
rect 29549 14909 29561 14943
rect 29595 14909 29607 14943
rect 29549 14903 29607 14909
rect 29825 14943 29883 14949
rect 29825 14909 29837 14943
rect 29871 14909 29883 14943
rect 29825 14903 29883 14909
rect 29564 14872 29592 14903
rect 28828 14844 29592 14872
rect 29380 14816 29408 14844
rect 24302 14804 24308 14816
rect 23860 14776 24308 14804
rect 24302 14764 24308 14776
rect 24360 14764 24366 14816
rect 29362 14764 29368 14816
rect 29420 14764 29426 14816
rect 29638 14764 29644 14816
rect 29696 14764 29702 14816
rect 552 14714 31531 14736
rect 552 14662 8102 14714
rect 8154 14662 8166 14714
rect 8218 14662 8230 14714
rect 8282 14662 8294 14714
rect 8346 14662 8358 14714
rect 8410 14662 15807 14714
rect 15859 14662 15871 14714
rect 15923 14662 15935 14714
rect 15987 14662 15999 14714
rect 16051 14662 16063 14714
rect 16115 14662 23512 14714
rect 23564 14662 23576 14714
rect 23628 14662 23640 14714
rect 23692 14662 23704 14714
rect 23756 14662 23768 14714
rect 23820 14662 31217 14714
rect 31269 14662 31281 14714
rect 31333 14662 31345 14714
rect 31397 14662 31409 14714
rect 31461 14662 31473 14714
rect 31525 14662 31531 14714
rect 552 14640 31531 14662
rect 1762 14560 1768 14612
rect 1820 14560 1826 14612
rect 2222 14560 2228 14612
rect 2280 14560 2286 14612
rect 4157 14603 4215 14609
rect 4157 14569 4169 14603
rect 4203 14600 4215 14603
rect 5350 14600 5356 14612
rect 4203 14572 5356 14600
rect 4203 14569 4215 14572
rect 4157 14563 4215 14569
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 7929 14603 7987 14609
rect 7929 14569 7941 14603
rect 7975 14569 7987 14603
rect 7929 14563 7987 14569
rect 9401 14603 9459 14609
rect 9401 14569 9413 14603
rect 9447 14600 9459 14603
rect 9674 14600 9680 14612
rect 9447 14572 9680 14600
rect 9447 14569 9459 14572
rect 9401 14563 9459 14569
rect 1780 14532 1808 14560
rect 1412 14504 1808 14532
rect 1412 14473 1440 14504
rect 2240 14473 2268 14560
rect 2314 14492 2320 14544
rect 2372 14532 2378 14544
rect 3022 14535 3080 14541
rect 3022 14532 3034 14535
rect 2372 14504 3034 14532
rect 2372 14492 2378 14504
rect 2516 14473 2544 14504
rect 3022 14501 3034 14504
rect 3068 14501 3080 14535
rect 4706 14532 4712 14544
rect 3022 14495 3080 14501
rect 4632 14504 4712 14532
rect 4632 14473 4660 14504
rect 4706 14492 4712 14504
rect 4764 14492 4770 14544
rect 7944 14532 7972 14563
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 10502 14560 10508 14612
rect 10560 14560 10566 14612
rect 14182 14600 14188 14612
rect 13832 14572 14188 14600
rect 13725 14535 13783 14541
rect 13725 14532 13737 14535
rect 7944 14504 13737 14532
rect 13725 14501 13737 14504
rect 13771 14501 13783 14535
rect 13725 14495 13783 14501
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14433 1455 14467
rect 1397 14427 1455 14433
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14464 1731 14467
rect 1949 14467 2007 14473
rect 1949 14464 1961 14467
rect 1719 14436 1961 14464
rect 1719 14433 1731 14436
rect 1673 14427 1731 14433
rect 1949 14433 1961 14436
rect 1995 14433 2007 14467
rect 1949 14427 2007 14433
rect 2225 14467 2283 14473
rect 2225 14433 2237 14467
rect 2271 14433 2283 14467
rect 2225 14427 2283 14433
rect 2501 14467 2559 14473
rect 2501 14433 2513 14467
rect 2547 14433 2559 14467
rect 2501 14427 2559 14433
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14433 4675 14467
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 4617 14427 4675 14433
rect 4908 14436 5089 14464
rect 1578 14356 1584 14408
rect 1636 14356 1642 14408
rect 1305 14331 1363 14337
rect 1305 14297 1317 14331
rect 1351 14328 1363 14331
rect 1394 14328 1400 14340
rect 1351 14300 1400 14328
rect 1351 14297 1363 14300
rect 1305 14291 1363 14297
rect 1394 14288 1400 14300
rect 1452 14328 1458 14340
rect 1964 14328 1992 14427
rect 2682 14356 2688 14408
rect 2740 14396 2746 14408
rect 2777 14399 2835 14405
rect 2777 14396 2789 14399
rect 2740 14368 2789 14396
rect 2740 14356 2746 14368
rect 2777 14365 2789 14368
rect 2823 14365 2835 14399
rect 2777 14359 2835 14365
rect 2133 14331 2191 14337
rect 2133 14328 2145 14331
rect 1452 14300 1624 14328
rect 1964 14300 2145 14328
rect 1452 14288 1458 14300
rect 1596 14260 1624 14300
rect 2133 14297 2145 14300
rect 2179 14328 2191 14331
rect 2409 14331 2467 14337
rect 2409 14328 2421 14331
rect 2179 14300 2421 14328
rect 2179 14297 2191 14300
rect 2133 14291 2191 14297
rect 2409 14297 2421 14300
rect 2455 14297 2467 14331
rect 2409 14291 2467 14297
rect 4908 14272 4936 14436
rect 5077 14433 5089 14436
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 5813 14467 5871 14473
rect 5813 14433 5825 14467
rect 5859 14433 5871 14467
rect 5813 14427 5871 14433
rect 5828 14396 5856 14427
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 6181 14467 6239 14473
rect 6181 14464 6193 14467
rect 5960 14436 6193 14464
rect 5960 14424 5966 14436
rect 6181 14433 6193 14436
rect 6227 14433 6239 14467
rect 6181 14427 6239 14433
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 6549 14467 6607 14473
rect 6549 14464 6561 14467
rect 6512 14436 6561 14464
rect 6512 14424 6518 14436
rect 6549 14433 6561 14436
rect 6595 14433 6607 14467
rect 6805 14467 6863 14473
rect 6805 14464 6817 14467
rect 6549 14427 6607 14433
rect 6656 14436 6817 14464
rect 6270 14396 6276 14408
rect 5000 14368 6276 14396
rect 5000 14272 5028 14368
rect 6270 14356 6276 14368
rect 6328 14396 6334 14408
rect 6656 14396 6684 14436
rect 6805 14433 6817 14436
rect 6851 14433 6863 14467
rect 6805 14427 6863 14433
rect 9493 14467 9551 14473
rect 9493 14433 9505 14467
rect 9539 14433 9551 14467
rect 9493 14427 9551 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 9766 14464 9772 14476
rect 9631 14436 9772 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 6328 14368 6684 14396
rect 9508 14396 9536 14427
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 9876 14436 10057 14464
rect 9876 14408 9904 14436
rect 10045 14433 10057 14436
rect 10091 14433 10103 14467
rect 10045 14427 10103 14433
rect 10321 14467 10379 14473
rect 10321 14433 10333 14467
rect 10367 14464 10379 14467
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 10367 14436 10425 14464
rect 10367 14433 10379 14436
rect 10321 14427 10379 14433
rect 10413 14433 10425 14436
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 11054 14464 11060 14476
rect 11011 14436 11060 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 9858 14396 9864 14408
rect 9508 14368 9864 14396
rect 6328 14356 6334 14368
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 10336 14396 10364 14427
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 11238 14473 11244 14476
rect 11232 14427 11244 14473
rect 11238 14424 11244 14427
rect 11296 14424 11302 14476
rect 12621 14467 12679 14473
rect 12621 14464 12633 14467
rect 12452 14436 12633 14464
rect 12452 14408 12480 14436
rect 12621 14433 12633 14436
rect 12667 14433 12679 14467
rect 12621 14427 12679 14433
rect 13078 14424 13084 14476
rect 13136 14424 13142 14476
rect 13173 14467 13231 14473
rect 13173 14433 13185 14467
rect 13219 14464 13231 14467
rect 13609 14467 13667 14473
rect 13609 14464 13621 14467
rect 13219 14436 13621 14464
rect 13219 14433 13231 14436
rect 13173 14427 13231 14433
rect 13609 14433 13621 14436
rect 13655 14464 13667 14467
rect 13832 14464 13860 14572
rect 14182 14560 14188 14572
rect 14240 14600 14246 14612
rect 15381 14603 15439 14609
rect 15381 14600 15393 14603
rect 14240 14572 15393 14600
rect 14240 14560 14246 14572
rect 15381 14569 15393 14572
rect 15427 14569 15439 14603
rect 15381 14563 15439 14569
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 20438 14600 20444 14612
rect 18288 14572 20444 14600
rect 18288 14560 18294 14572
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 20901 14603 20959 14609
rect 20901 14569 20913 14603
rect 20947 14569 20959 14603
rect 21910 14600 21916 14612
rect 20901 14563 20959 14569
rect 21468 14572 21916 14600
rect 13998 14541 14004 14544
rect 13941 14535 14004 14541
rect 13941 14501 13953 14535
rect 13987 14501 14004 14535
rect 13941 14495 14004 14501
rect 13998 14492 14004 14495
rect 14056 14532 14062 14544
rect 15010 14532 15016 14544
rect 14056 14504 15016 14532
rect 14056 14492 14062 14504
rect 15010 14492 15016 14504
rect 15068 14492 15074 14544
rect 19334 14532 19340 14544
rect 15120 14504 15332 14532
rect 13655 14436 13860 14464
rect 14185 14467 14243 14473
rect 13655 14433 13667 14436
rect 13609 14427 13667 14433
rect 14185 14433 14197 14467
rect 14231 14433 14243 14467
rect 14185 14427 14243 14433
rect 9968 14368 10364 14396
rect 9968 14337 9996 14368
rect 12434 14356 12440 14408
rect 12492 14356 12498 14408
rect 12989 14399 13047 14405
rect 12989 14365 13001 14399
rect 13035 14396 13047 14399
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 13035 14368 13277 14396
rect 13035 14365 13047 14368
rect 12989 14359 13047 14365
rect 13265 14365 13277 14368
rect 13311 14396 13323 14399
rect 13354 14396 13360 14408
rect 13311 14368 13360 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 13354 14356 13360 14368
rect 13412 14396 13418 14408
rect 14200 14396 14228 14427
rect 14458 14424 14464 14476
rect 14516 14464 14522 14476
rect 15120 14473 15148 14504
rect 14737 14467 14795 14473
rect 14737 14464 14749 14467
rect 14516 14436 14749 14464
rect 14516 14424 14522 14436
rect 14737 14433 14749 14436
rect 14783 14464 14795 14467
rect 15105 14467 15163 14473
rect 15105 14464 15117 14467
rect 14783 14436 15117 14464
rect 14783 14433 14795 14436
rect 14737 14427 14795 14433
rect 15105 14433 15117 14436
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 15194 14424 15200 14476
rect 15252 14424 15258 14476
rect 15304 14473 15332 14504
rect 16592 14504 19340 14532
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 16206 14424 16212 14476
rect 16264 14464 16270 14476
rect 16592 14473 16620 14504
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 16577 14467 16635 14473
rect 16577 14464 16589 14467
rect 16264 14436 16589 14464
rect 16264 14424 16270 14436
rect 16577 14433 16589 14436
rect 16623 14433 16635 14467
rect 16833 14467 16891 14473
rect 16833 14464 16845 14467
rect 16577 14427 16635 14433
rect 16684 14436 16845 14464
rect 13412 14368 14228 14396
rect 15212 14396 15240 14424
rect 16684 14396 16712 14436
rect 16833 14433 16845 14436
rect 16879 14433 16891 14467
rect 19352 14464 19380 14492
rect 19794 14473 19800 14476
rect 19528 14467 19586 14473
rect 19352 14462 19472 14464
rect 19528 14462 19540 14467
rect 19352 14436 19540 14462
rect 19444 14434 19540 14436
rect 16833 14427 16891 14433
rect 19528 14433 19540 14434
rect 19574 14433 19586 14467
rect 19528 14427 19586 14433
rect 19777 14467 19800 14473
rect 19777 14433 19789 14467
rect 19777 14427 19800 14433
rect 19794 14424 19800 14427
rect 19852 14424 19858 14476
rect 15212 14368 16712 14396
rect 13412 14356 13418 14368
rect 17862 14356 17868 14408
rect 17920 14396 17926 14408
rect 19058 14396 19064 14408
rect 17920 14368 19064 14396
rect 17920 14356 17926 14368
rect 19058 14356 19064 14368
rect 19116 14356 19122 14408
rect 20916 14396 20944 14563
rect 21468 14541 21496 14572
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 22960 14572 23796 14600
rect 21453 14535 21511 14541
rect 21453 14501 21465 14535
rect 21499 14501 21511 14535
rect 22189 14535 22247 14541
rect 22189 14532 22201 14535
rect 21453 14495 21511 14501
rect 21652 14504 22201 14532
rect 21652 14476 21680 14504
rect 22189 14501 22201 14504
rect 22235 14501 22247 14535
rect 22189 14495 22247 14501
rect 22327 14535 22385 14541
rect 22327 14501 22339 14535
rect 22373 14532 22385 14535
rect 22373 14501 22407 14532
rect 22960 14507 22988 14572
rect 22327 14495 22407 14501
rect 21634 14424 21640 14476
rect 21692 14424 21698 14476
rect 22379 14396 22407 14495
rect 22511 14501 22569 14507
rect 22511 14467 22523 14501
rect 22557 14498 22569 14501
rect 22960 14501 23029 14507
rect 22557 14476 22591 14498
rect 22960 14476 22983 14501
rect 22557 14467 22560 14476
rect 22511 14461 22560 14467
rect 22554 14424 22560 14461
rect 22612 14424 22618 14476
rect 22922 14424 22928 14476
rect 22980 14467 22983 14476
rect 23017 14467 23029 14501
rect 23198 14492 23204 14544
rect 23256 14492 23262 14544
rect 23431 14501 23489 14507
rect 22980 14461 23029 14467
rect 23431 14467 23443 14501
rect 23477 14498 23489 14501
rect 23477 14467 23499 14498
rect 23658 14492 23664 14544
rect 23716 14492 23722 14544
rect 23768 14532 23796 14572
rect 26786 14560 26792 14612
rect 26844 14600 26850 14612
rect 27433 14603 27491 14609
rect 27433 14600 27445 14603
rect 26844 14572 27445 14600
rect 26844 14560 26850 14572
rect 27433 14569 27445 14572
rect 27479 14600 27491 14603
rect 28813 14603 28871 14609
rect 27479 14572 28488 14600
rect 27479 14569 27491 14572
rect 27433 14563 27491 14569
rect 24825 14535 24883 14541
rect 24825 14532 24837 14535
rect 23768 14504 24837 14532
rect 24825 14501 24837 14504
rect 24871 14501 24883 14535
rect 24825 14495 24883 14501
rect 24946 14492 24952 14544
rect 25004 14532 25010 14544
rect 25041 14535 25099 14541
rect 25041 14532 25053 14535
rect 25004 14504 25053 14532
rect 25004 14492 25010 14504
rect 25041 14501 25053 14504
rect 25087 14501 25099 14535
rect 25041 14495 25099 14501
rect 27709 14535 27767 14541
rect 27709 14501 27721 14535
rect 27755 14532 27767 14535
rect 28261 14535 28319 14541
rect 28261 14532 28273 14535
rect 27755 14504 28273 14532
rect 27755 14501 27767 14504
rect 27709 14495 27767 14501
rect 28261 14501 28273 14504
rect 28307 14501 28319 14535
rect 28261 14495 28319 14501
rect 28460 14532 28488 14572
rect 28813 14569 28825 14603
rect 28859 14600 28871 14603
rect 29178 14600 29184 14612
rect 28859 14572 29184 14600
rect 28859 14569 28871 14572
rect 28813 14563 28871 14569
rect 29178 14560 29184 14572
rect 29236 14600 29242 14612
rect 29365 14603 29423 14609
rect 29365 14600 29377 14603
rect 29236 14572 29377 14600
rect 29236 14560 29242 14572
rect 29365 14569 29377 14572
rect 29411 14569 29423 14603
rect 30929 14603 30987 14609
rect 30929 14600 30941 14603
rect 29365 14563 29423 14569
rect 29472 14572 30941 14600
rect 28460 14504 28764 14532
rect 23431 14464 23499 14467
rect 23431 14461 23520 14464
rect 22980 14436 22988 14461
rect 23471 14436 23520 14461
rect 22980 14424 22986 14436
rect 23492 14408 23520 14436
rect 23934 14424 23940 14476
rect 23992 14424 23998 14476
rect 24026 14424 24032 14476
rect 24084 14464 24090 14476
rect 24084 14436 24129 14464
rect 24084 14424 24090 14436
rect 24210 14424 24216 14476
rect 24268 14424 24274 14476
rect 24305 14467 24363 14473
rect 24305 14433 24317 14467
rect 24351 14433 24363 14467
rect 24305 14427 24363 14433
rect 24443 14467 24501 14473
rect 24443 14433 24455 14467
rect 24489 14464 24501 14467
rect 24578 14464 24584 14476
rect 24489 14436 24584 14464
rect 24489 14433 24501 14436
rect 24443 14427 24501 14433
rect 23474 14396 23480 14408
rect 20916 14368 22407 14396
rect 23124 14368 23480 14396
rect 9677 14331 9735 14337
rect 9677 14297 9689 14331
rect 9723 14328 9735 14331
rect 9953 14331 10011 14337
rect 9953 14328 9965 14331
rect 9723 14300 9965 14328
rect 9723 14297 9735 14300
rect 9677 14291 9735 14297
rect 9953 14297 9965 14300
rect 9999 14297 10011 14331
rect 12529 14331 12587 14337
rect 12529 14328 12541 14331
rect 9953 14291 10011 14297
rect 11900 14300 12541 14328
rect 1857 14263 1915 14269
rect 1857 14260 1869 14263
rect 1596 14232 1869 14260
rect 1857 14229 1869 14232
rect 1903 14229 1915 14263
rect 1857 14223 1915 14229
rect 4709 14263 4767 14269
rect 4709 14229 4721 14263
rect 4755 14260 4767 14263
rect 4890 14260 4896 14272
rect 4755 14232 4896 14260
rect 4755 14229 4767 14232
rect 4709 14223 4767 14229
rect 4890 14220 4896 14232
rect 4948 14220 4954 14272
rect 4982 14220 4988 14272
rect 5040 14220 5046 14272
rect 6086 14220 6092 14272
rect 6144 14260 6150 14272
rect 6273 14263 6331 14269
rect 6273 14260 6285 14263
rect 6144 14232 6285 14260
rect 6144 14220 6150 14232
rect 6273 14229 6285 14232
rect 6319 14229 6331 14263
rect 6273 14223 6331 14229
rect 10134 14220 10140 14272
rect 10192 14260 10198 14272
rect 10229 14263 10287 14269
rect 10229 14260 10241 14263
rect 10192 14232 10241 14260
rect 10192 14220 10198 14232
rect 10229 14229 10241 14232
rect 10275 14229 10287 14263
rect 10229 14223 10287 14229
rect 11698 14220 11704 14272
rect 11756 14260 11762 14272
rect 11900 14260 11928 14300
rect 12529 14297 12541 14300
rect 12575 14328 12587 14331
rect 13541 14331 13599 14337
rect 13541 14328 13553 14331
rect 12575 14300 13553 14328
rect 12575 14297 12587 14300
rect 12529 14291 12587 14297
rect 13541 14297 13553 14300
rect 13587 14297 13599 14331
rect 15470 14328 15476 14340
rect 13541 14291 13599 14297
rect 13924 14300 15476 14328
rect 11756 14232 11928 14260
rect 11756 14220 11762 14232
rect 12342 14220 12348 14272
rect 12400 14220 12406 14272
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 13924 14269 13952 14300
rect 15470 14288 15476 14300
rect 15528 14288 15534 14340
rect 19426 14328 19432 14340
rect 17512 14300 19432 14328
rect 13909 14263 13967 14269
rect 13909 14260 13921 14263
rect 13320 14232 13921 14260
rect 13320 14220 13326 14232
rect 13909 14229 13921 14232
rect 13955 14229 13967 14263
rect 13909 14223 13967 14229
rect 14093 14263 14151 14269
rect 14093 14229 14105 14263
rect 14139 14260 14151 14263
rect 14182 14260 14188 14272
rect 14139 14232 14188 14260
rect 14139 14229 14151 14232
rect 14093 14223 14151 14229
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 14829 14263 14887 14269
rect 14829 14260 14841 14263
rect 14332 14232 14841 14260
rect 14332 14220 14338 14232
rect 14829 14229 14841 14232
rect 14875 14229 14887 14263
rect 14829 14223 14887 14229
rect 15286 14220 15292 14272
rect 15344 14260 15350 14272
rect 17512 14260 17540 14300
rect 19426 14288 19432 14300
rect 19484 14288 19490 14340
rect 15344 14232 17540 14260
rect 15344 14220 15350 14232
rect 17954 14220 17960 14272
rect 18012 14220 18018 14272
rect 18874 14220 18880 14272
rect 18932 14260 18938 14272
rect 21082 14260 21088 14272
rect 18932 14232 21088 14260
rect 18932 14220 18938 14232
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 22278 14220 22284 14272
rect 22336 14260 22342 14272
rect 22465 14263 22523 14269
rect 22465 14260 22477 14263
rect 22336 14232 22477 14260
rect 22336 14220 22342 14232
rect 22465 14229 22477 14232
rect 22511 14229 22523 14263
rect 22465 14223 22523 14229
rect 22646 14220 22652 14272
rect 22704 14220 22710 14272
rect 22830 14220 22836 14272
rect 22888 14220 22894 14272
rect 23017 14263 23075 14269
rect 23017 14229 23029 14263
rect 23063 14260 23075 14263
rect 23124 14260 23152 14368
rect 23474 14356 23480 14368
rect 23532 14356 23538 14408
rect 24320 14396 24348 14427
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 26421 14467 26479 14473
rect 26421 14433 26433 14467
rect 26467 14433 26479 14467
rect 26421 14427 26479 14433
rect 26513 14467 26571 14473
rect 26513 14433 26525 14467
rect 26559 14464 26571 14467
rect 26786 14464 26792 14476
rect 26559 14436 26792 14464
rect 26559 14433 26571 14436
rect 26513 14427 26571 14433
rect 26436 14396 26464 14427
rect 26786 14424 26792 14436
rect 26844 14464 26850 14476
rect 26881 14467 26939 14473
rect 26881 14464 26893 14467
rect 26844 14436 26893 14464
rect 26844 14424 26850 14436
rect 26881 14433 26893 14436
rect 26927 14433 26939 14467
rect 26881 14427 26939 14433
rect 27525 14467 27583 14473
rect 27525 14433 27537 14467
rect 27571 14433 27583 14467
rect 27525 14427 27583 14433
rect 27617 14467 27675 14473
rect 27617 14433 27629 14467
rect 27663 14464 27675 14467
rect 27798 14464 27804 14476
rect 27663 14436 27804 14464
rect 27663 14433 27675 14436
rect 27617 14427 27675 14433
rect 26602 14396 26608 14408
rect 24320 14368 24440 14396
rect 26436 14368 26608 14396
rect 24412 14328 24440 14368
rect 26602 14356 26608 14368
rect 26660 14356 26666 14408
rect 27540 14396 27568 14427
rect 27798 14424 27804 14436
rect 27856 14424 27862 14476
rect 27893 14467 27951 14473
rect 27893 14433 27905 14467
rect 27939 14433 27951 14467
rect 27893 14427 27951 14433
rect 27706 14396 27712 14408
rect 27540 14368 27712 14396
rect 27706 14356 27712 14368
rect 27764 14396 27770 14408
rect 27908 14396 27936 14427
rect 27764 14368 27936 14396
rect 28276 14396 28304 14495
rect 28353 14467 28411 14473
rect 28353 14433 28365 14467
rect 28399 14462 28411 14467
rect 28460 14462 28488 14504
rect 28736 14473 28764 14504
rect 28902 14492 28908 14544
rect 28960 14532 28966 14544
rect 29472 14532 29500 14572
rect 30929 14569 30941 14572
rect 30975 14569 30987 14603
rect 30929 14563 30987 14569
rect 28960 14504 29500 14532
rect 28960 14492 28966 14504
rect 29546 14492 29552 14544
rect 29604 14492 29610 14544
rect 29638 14492 29644 14544
rect 29696 14532 29702 14544
rect 29794 14535 29852 14541
rect 29794 14532 29806 14535
rect 29696 14504 29806 14532
rect 29696 14492 29702 14504
rect 29794 14501 29806 14504
rect 29840 14501 29852 14535
rect 29794 14495 29852 14501
rect 28399 14434 28488 14462
rect 28629 14467 28687 14473
rect 28399 14433 28411 14434
rect 28353 14427 28411 14433
rect 28629 14433 28641 14467
rect 28675 14433 28687 14467
rect 28629 14427 28687 14433
rect 28721 14467 28779 14473
rect 28721 14433 28733 14467
rect 28767 14433 28779 14467
rect 28721 14427 28779 14433
rect 28997 14467 29055 14473
rect 28997 14433 29009 14467
rect 29043 14433 29055 14467
rect 28997 14427 29055 14433
rect 29457 14467 29515 14473
rect 29457 14433 29469 14467
rect 29503 14433 29515 14467
rect 29457 14427 29515 14433
rect 28644 14396 28672 14427
rect 29012 14396 29040 14427
rect 28276 14368 29040 14396
rect 27764 14356 27770 14368
rect 28074 14328 28080 14340
rect 24412 14300 28080 14328
rect 28074 14288 28080 14300
rect 28132 14288 28138 14340
rect 29270 14328 29276 14340
rect 28552 14300 29276 14328
rect 23063 14232 23152 14260
rect 23063 14229 23075 14232
rect 23017 14223 23075 14229
rect 23290 14220 23296 14272
rect 23348 14220 23354 14272
rect 23477 14263 23535 14269
rect 23477 14229 23489 14263
rect 23523 14260 23535 14263
rect 23934 14260 23940 14272
rect 23523 14232 23940 14260
rect 23523 14229 23535 14232
rect 23477 14223 23535 14229
rect 23934 14220 23940 14232
rect 23992 14220 23998 14272
rect 24026 14220 24032 14272
rect 24084 14260 24090 14272
rect 24581 14263 24639 14269
rect 24581 14260 24593 14263
rect 24084 14232 24593 14260
rect 24084 14220 24090 14232
rect 24581 14229 24593 14232
rect 24627 14229 24639 14263
rect 24581 14223 24639 14229
rect 24670 14220 24676 14272
rect 24728 14220 24734 14272
rect 24854 14220 24860 14272
rect 24912 14220 24918 14272
rect 28552 14269 28580 14300
rect 29270 14288 29276 14300
rect 29328 14328 29334 14340
rect 29472 14328 29500 14427
rect 29564 14405 29592 14492
rect 29549 14399 29607 14405
rect 29549 14365 29561 14399
rect 29595 14365 29607 14399
rect 29549 14359 29607 14365
rect 29328 14300 29500 14328
rect 29328 14288 29334 14300
rect 27985 14263 28043 14269
rect 27985 14229 27997 14263
rect 28031 14260 28043 14263
rect 28537 14263 28595 14269
rect 28537 14260 28549 14263
rect 28031 14232 28549 14260
rect 28031 14229 28043 14232
rect 27985 14223 28043 14229
rect 28537 14229 28549 14232
rect 28583 14229 28595 14263
rect 28537 14223 28595 14229
rect 29089 14263 29147 14269
rect 29089 14229 29101 14263
rect 29135 14260 29147 14263
rect 29454 14260 29460 14272
rect 29135 14232 29460 14260
rect 29135 14229 29147 14232
rect 29089 14223 29147 14229
rect 29454 14220 29460 14232
rect 29512 14220 29518 14272
rect 552 14170 31372 14192
rect 552 14118 4250 14170
rect 4302 14118 4314 14170
rect 4366 14118 4378 14170
rect 4430 14118 4442 14170
rect 4494 14118 4506 14170
rect 4558 14118 11955 14170
rect 12007 14118 12019 14170
rect 12071 14118 12083 14170
rect 12135 14118 12147 14170
rect 12199 14118 12211 14170
rect 12263 14118 19660 14170
rect 19712 14118 19724 14170
rect 19776 14118 19788 14170
rect 19840 14118 19852 14170
rect 19904 14118 19916 14170
rect 19968 14118 27365 14170
rect 27417 14118 27429 14170
rect 27481 14118 27493 14170
rect 27545 14118 27557 14170
rect 27609 14118 27621 14170
rect 27673 14118 31372 14170
rect 552 14096 31372 14118
rect 1489 14059 1547 14065
rect 1489 14025 1501 14059
rect 1535 14056 1547 14059
rect 1578 14056 1584 14068
rect 1535 14028 1584 14056
rect 1535 14025 1547 14028
rect 1489 14019 1547 14025
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 2682 14056 2688 14068
rect 1688 14028 2688 14056
rect 1210 13880 1216 13932
rect 1268 13920 1274 13932
rect 1688 13929 1716 14028
rect 2682 14016 2688 14028
rect 2740 14016 2746 14068
rect 4341 14059 4399 14065
rect 4341 14025 4353 14059
rect 4387 14056 4399 14059
rect 4982 14056 4988 14068
rect 4387 14028 4988 14056
rect 4387 14025 4399 14028
rect 4341 14019 4399 14025
rect 4982 14016 4988 14028
rect 5040 14016 5046 14068
rect 5902 14016 5908 14068
rect 5960 14016 5966 14068
rect 6457 14059 6515 14065
rect 6457 14025 6469 14059
rect 6503 14056 6515 14059
rect 6733 14059 6791 14065
rect 6733 14056 6745 14059
rect 6503 14028 6745 14056
rect 6503 14025 6515 14028
rect 6457 14019 6515 14025
rect 6733 14025 6745 14028
rect 6779 14056 6791 14059
rect 6914 14056 6920 14068
rect 6779 14028 6920 14056
rect 6779 14025 6791 14028
rect 6733 14019 6791 14025
rect 6914 14016 6920 14028
rect 6972 14056 6978 14068
rect 7834 14056 7840 14068
rect 6972 14028 7840 14056
rect 6972 14016 6978 14028
rect 7834 14016 7840 14028
rect 7892 14016 7898 14068
rect 12897 14059 12955 14065
rect 9784 14028 11928 14056
rect 3053 13991 3111 13997
rect 3053 13957 3065 13991
rect 3099 13988 3111 13991
rect 3970 13988 3976 14000
rect 3099 13960 3976 13988
rect 3099 13957 3111 13960
rect 3053 13951 3111 13957
rect 3970 13948 3976 13960
rect 4028 13948 4034 14000
rect 1673 13923 1731 13929
rect 1268 13892 1440 13920
rect 1268 13880 1274 13892
rect 1412 13861 1440 13892
rect 1673 13889 1685 13923
rect 1719 13889 1731 13923
rect 5353 13923 5411 13929
rect 1673 13883 1731 13889
rect 4816 13892 5304 13920
rect 4157 13865 4215 13871
rect 1305 13855 1363 13861
rect 1305 13821 1317 13855
rect 1351 13821 1363 13855
rect 1305 13815 1363 13821
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13821 1455 13855
rect 1940 13855 1998 13861
rect 1940 13852 1952 13855
rect 1397 13815 1455 13821
rect 1504 13824 1952 13852
rect 1320 13784 1348 13815
rect 1504 13784 1532 13824
rect 1940 13821 1952 13824
rect 1986 13852 1998 13855
rect 2222 13852 2228 13864
rect 1986 13824 2228 13852
rect 1986 13821 1998 13824
rect 1940 13815 1998 13821
rect 2222 13812 2228 13824
rect 2280 13812 2286 13864
rect 4157 13831 4169 13865
rect 4203 13831 4215 13865
rect 4816 13861 4844 13892
rect 4157 13825 4215 13831
rect 4249 13855 4307 13861
rect 4172 13796 4200 13825
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 4525 13855 4583 13861
rect 4525 13852 4537 13855
rect 4295 13824 4537 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 4525 13821 4537 13824
rect 4571 13821 4583 13855
rect 4525 13815 4583 13821
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 4801 13855 4859 13861
rect 4801 13852 4813 13855
rect 4663 13824 4813 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 4801 13821 4813 13824
rect 4847 13821 4859 13855
rect 4801 13815 4859 13821
rect 1320 13756 1532 13784
rect 4154 13744 4160 13796
rect 4212 13744 4218 13796
rect 4065 13719 4123 13725
rect 4065 13685 4077 13719
rect 4111 13716 4123 13719
rect 4540 13716 4568 13815
rect 4890 13812 4896 13864
rect 4948 13852 4954 13864
rect 5276 13861 5304 13892
rect 5353 13889 5365 13923
rect 5399 13920 5411 13923
rect 5920 13920 5948 14016
rect 6086 13948 6092 14000
rect 6144 13988 6150 14000
rect 9784 13997 9812 14028
rect 7929 13991 7987 13997
rect 7929 13988 7941 13991
rect 6144 13960 7941 13988
rect 6144 13948 6150 13960
rect 5399 13892 5948 13920
rect 5399 13889 5411 13892
rect 5353 13883 5411 13889
rect 5261 13855 5319 13861
rect 4948 13824 5212 13852
rect 4948 13812 4954 13824
rect 5184 13784 5212 13824
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 5442 13852 5448 13864
rect 5307 13824 5448 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 5644 13861 5672 13892
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 7558 13920 7564 13932
rect 6328 13892 6408 13920
rect 6328 13880 6334 13892
rect 6380 13861 6408 13892
rect 6748 13892 7564 13920
rect 5629 13855 5687 13861
rect 5629 13821 5641 13855
rect 5675 13821 5687 13855
rect 5905 13855 5963 13861
rect 5905 13852 5917 13855
rect 5629 13815 5687 13821
rect 5736 13824 5917 13852
rect 5736 13784 5764 13824
rect 5905 13821 5917 13824
rect 5951 13821 5963 13855
rect 5905 13815 5963 13821
rect 6365 13855 6423 13861
rect 6365 13821 6377 13855
rect 6411 13821 6423 13855
rect 6365 13815 6423 13821
rect 6748 13846 6776 13892
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 7852 13920 7880 13960
rect 7929 13957 7941 13960
rect 7975 13957 7987 13991
rect 7929 13951 7987 13957
rect 9769 13991 9827 13997
rect 9769 13957 9781 13991
rect 9815 13957 9827 13991
rect 9769 13951 9827 13957
rect 7760 13892 7880 13920
rect 6817 13849 6875 13855
rect 6817 13846 6829 13849
rect 6748 13818 6829 13846
rect 5184 13756 5764 13784
rect 5166 13716 5172 13728
rect 4111 13688 5172 13716
rect 4111 13685 4123 13688
rect 4065 13679 4123 13685
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 5721 13719 5779 13725
rect 5721 13685 5733 13719
rect 5767 13716 5779 13719
rect 5997 13719 6055 13725
rect 5997 13716 6009 13719
rect 5767 13688 6009 13716
rect 5767 13685 5779 13688
rect 5721 13679 5779 13685
rect 5997 13685 6009 13688
rect 6043 13716 6055 13719
rect 6748 13716 6776 13818
rect 6817 13815 6829 13818
rect 6863 13815 6875 13849
rect 6817 13809 6875 13815
rect 6914 13812 6920 13864
rect 6972 13812 6978 13864
rect 7469 13855 7527 13861
rect 7469 13821 7481 13855
rect 7515 13852 7527 13855
rect 7650 13852 7656 13864
rect 7515 13824 7656 13852
rect 7515 13821 7527 13824
rect 7469 13815 7527 13821
rect 7650 13812 7656 13824
rect 7708 13812 7714 13864
rect 7760 13861 7788 13892
rect 8018 13880 8024 13932
rect 8076 13920 8082 13932
rect 8386 13920 8392 13932
rect 8076 13892 8392 13920
rect 8076 13880 8082 13892
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 7834 13812 7840 13864
rect 7892 13812 7898 13864
rect 9861 13855 9919 13861
rect 9861 13821 9873 13855
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 11609 13855 11667 13861
rect 11609 13821 11621 13855
rect 11655 13852 11667 13855
rect 11698 13852 11704 13864
rect 11655 13824 11704 13852
rect 11655 13821 11667 13824
rect 11609 13815 11667 13821
rect 8478 13744 8484 13796
rect 8536 13784 8542 13796
rect 8634 13787 8692 13793
rect 8634 13784 8646 13787
rect 8536 13756 8646 13784
rect 8536 13744 8542 13756
rect 8634 13753 8646 13756
rect 8680 13753 8692 13787
rect 8634 13747 8692 13753
rect 6043 13688 6776 13716
rect 7009 13719 7067 13725
rect 6043 13685 6055 13688
rect 5997 13679 6055 13685
rect 7009 13685 7021 13719
rect 7055 13716 7067 13719
rect 7377 13719 7435 13725
rect 7377 13716 7389 13719
rect 7055 13688 7389 13716
rect 7055 13685 7067 13688
rect 7009 13679 7067 13685
rect 7377 13685 7389 13688
rect 7423 13716 7435 13719
rect 7466 13716 7472 13728
rect 7423 13688 7472 13716
rect 7423 13685 7435 13688
rect 7377 13679 7435 13685
rect 7466 13676 7472 13688
rect 7524 13676 7530 13728
rect 9876 13716 9904 13815
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 10134 13793 10140 13796
rect 10128 13784 10140 13793
rect 10095 13756 10140 13784
rect 10128 13747 10140 13756
rect 10134 13744 10140 13747
rect 10192 13744 10198 13796
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 10836 13756 11805 13784
rect 10836 13744 10842 13756
rect 11793 13753 11805 13756
rect 11839 13753 11851 13787
rect 11793 13747 11851 13753
rect 10042 13716 10048 13728
rect 9876 13688 10048 13716
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 11238 13676 11244 13728
rect 11296 13676 11302 13728
rect 11514 13676 11520 13728
rect 11572 13676 11578 13728
rect 11900 13716 11928 14028
rect 12897 14025 12909 14059
rect 12943 14056 12955 14059
rect 13262 14056 13268 14068
rect 12943 14028 13268 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 13814 14016 13820 14068
rect 13872 14016 13878 14068
rect 14277 14059 14335 14065
rect 14277 14025 14289 14059
rect 14323 14056 14335 14059
rect 14323 14028 14780 14056
rect 14323 14025 14335 14028
rect 14277 14019 14335 14025
rect 14752 13988 14780 14028
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 15749 14059 15807 14065
rect 15749 14056 15761 14059
rect 15528 14028 15761 14056
rect 15528 14016 15534 14028
rect 15749 14025 15761 14028
rect 15795 14025 15807 14059
rect 15749 14019 15807 14025
rect 16393 14059 16451 14065
rect 16393 14025 16405 14059
rect 16439 14056 16451 14059
rect 17313 14059 17371 14065
rect 17313 14056 17325 14059
rect 16439 14028 17325 14056
rect 16439 14025 16451 14028
rect 16393 14019 16451 14025
rect 17313 14025 17325 14028
rect 17359 14025 17371 14059
rect 17313 14019 17371 14025
rect 15194 13988 15200 14000
rect 14752 13960 15200 13988
rect 14752 13932 14780 13960
rect 15194 13948 15200 13960
rect 15252 13948 15258 14000
rect 15933 13991 15991 13997
rect 15933 13957 15945 13991
rect 15979 13957 15991 13991
rect 17328 13988 17356 14019
rect 17494 14016 17500 14068
rect 17552 14056 17558 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 17552 14028 18889 14056
rect 17552 14016 17558 14028
rect 18877 14025 18889 14028
rect 18923 14056 18935 14059
rect 19978 14056 19984 14068
rect 18923 14028 19984 14056
rect 18923 14025 18935 14028
rect 18877 14019 18935 14025
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20070 14016 20076 14068
rect 20128 14056 20134 14068
rect 20165 14059 20223 14065
rect 20165 14056 20177 14059
rect 20128 14028 20177 14056
rect 20128 14016 20134 14028
rect 20165 14025 20177 14028
rect 20211 14025 20223 14059
rect 20165 14019 20223 14025
rect 20625 14059 20683 14065
rect 20625 14025 20637 14059
rect 20671 14056 20683 14059
rect 20990 14056 20996 14068
rect 20671 14028 20996 14056
rect 20671 14025 20683 14028
rect 20625 14019 20683 14025
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 21232 14028 21312 14056
rect 21232 14016 21238 14028
rect 18506 13988 18512 14000
rect 17328 13960 18512 13988
rect 15933 13951 15991 13957
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 14090 13920 14096 13932
rect 12492 13892 14096 13920
rect 12492 13880 12498 13892
rect 14090 13880 14096 13892
rect 14148 13920 14154 13932
rect 14274 13920 14280 13932
rect 14148 13892 14280 13920
rect 14148 13880 14154 13892
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 14734 13880 14740 13932
rect 14792 13880 14798 13932
rect 14826 13880 14832 13932
rect 14884 13880 14890 13932
rect 14918 13880 14924 13932
rect 14976 13920 14982 13932
rect 15286 13920 15292 13932
rect 14976 13892 15292 13920
rect 14976 13880 14982 13892
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 15948 13920 15976 13951
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 21284 13997 21312 14028
rect 21726 14016 21732 14068
rect 21784 14056 21790 14068
rect 22097 14059 22155 14065
rect 22097 14056 22109 14059
rect 21784 14028 22109 14056
rect 21784 14016 21790 14028
rect 22097 14025 22109 14028
rect 22143 14056 22155 14059
rect 22278 14056 22284 14068
rect 22143 14028 22284 14056
rect 22143 14025 22155 14028
rect 22097 14019 22155 14025
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 22646 14016 22652 14068
rect 22704 14016 22710 14068
rect 22830 14016 22836 14068
rect 22888 14056 22894 14068
rect 23109 14059 23167 14065
rect 23109 14056 23121 14059
rect 22888 14028 23121 14056
rect 22888 14016 22894 14028
rect 23109 14025 23121 14028
rect 23155 14025 23167 14059
rect 23109 14019 23167 14025
rect 23201 14059 23259 14065
rect 23201 14025 23213 14059
rect 23247 14056 23259 14059
rect 23290 14056 23296 14068
rect 23247 14028 23296 14056
rect 23247 14025 23259 14028
rect 23201 14019 23259 14025
rect 23290 14016 23296 14028
rect 23348 14016 23354 14068
rect 23474 14016 23480 14068
rect 23532 14056 23538 14068
rect 24029 14059 24087 14065
rect 24029 14056 24041 14059
rect 23532 14028 24041 14056
rect 23532 14016 23538 14028
rect 24029 14025 24041 14028
rect 24075 14056 24087 14059
rect 24854 14056 24860 14068
rect 24075 14028 24860 14056
rect 24075 14025 24087 14028
rect 24029 14019 24087 14025
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 26786 14016 26792 14068
rect 26844 14016 26850 14068
rect 27617 14059 27675 14065
rect 27617 14025 27629 14059
rect 27663 14056 27675 14059
rect 27706 14056 27712 14068
rect 27663 14028 27712 14056
rect 27663 14025 27675 14028
rect 27617 14019 27675 14025
rect 27706 14016 27712 14028
rect 27764 14056 27770 14068
rect 27893 14059 27951 14065
rect 27893 14056 27905 14059
rect 27764 14028 27905 14056
rect 27764 14016 27770 14028
rect 27893 14025 27905 14028
rect 27939 14025 27951 14059
rect 27893 14019 27951 14025
rect 29362 14016 29368 14068
rect 29420 14016 29426 14068
rect 30926 14016 30932 14068
rect 30984 14016 30990 14068
rect 19061 13991 19119 13997
rect 19061 13957 19073 13991
rect 19107 13988 19119 13991
rect 19429 13991 19487 13997
rect 19429 13988 19441 13991
rect 19107 13960 19441 13988
rect 19107 13957 19119 13960
rect 19061 13951 19119 13957
rect 19429 13957 19441 13960
rect 19475 13957 19487 13991
rect 19429 13951 19487 13957
rect 19521 13991 19579 13997
rect 19521 13957 19533 13991
rect 19567 13988 19579 13991
rect 20441 13991 20499 13997
rect 20441 13988 20453 13991
rect 19567 13960 20453 13988
rect 19567 13957 19579 13960
rect 19521 13951 19579 13957
rect 20441 13957 20453 13960
rect 20487 13957 20499 13991
rect 21269 13991 21327 13997
rect 20441 13951 20499 13957
rect 20548 13960 20760 13988
rect 19613 13923 19671 13929
rect 19613 13920 19625 13923
rect 15948 13892 19625 13920
rect 19613 13889 19625 13892
rect 19659 13889 19671 13923
rect 20548 13920 20576 13960
rect 19613 13883 19671 13889
rect 19720 13892 20576 13920
rect 20732 13920 20760 13960
rect 21269 13957 21281 13991
rect 21315 13988 21327 13991
rect 22370 13988 22376 14000
rect 21315 13960 22376 13988
rect 21315 13957 21327 13960
rect 21269 13951 21327 13957
rect 22370 13948 22376 13960
rect 22428 13948 22434 14000
rect 22664 13988 22692 14016
rect 23017 13991 23075 13997
rect 23017 13988 23029 13991
rect 22664 13960 23029 13988
rect 23017 13957 23029 13960
rect 23063 13957 23075 13991
rect 23017 13951 23075 13957
rect 24581 13991 24639 13997
rect 24581 13957 24593 13991
rect 24627 13957 24639 13991
rect 24581 13951 24639 13957
rect 24596 13920 24624 13951
rect 26602 13920 26608 13932
rect 20732 13892 24624 13920
rect 25884 13892 26608 13920
rect 13265 13855 13323 13861
rect 13265 13852 13277 13855
rect 12820 13824 13277 13852
rect 12158 13744 12164 13796
rect 12216 13784 12222 13796
rect 12621 13787 12679 13793
rect 12621 13784 12633 13787
rect 12216 13756 12633 13784
rect 12216 13744 12222 13756
rect 12621 13753 12633 13756
rect 12667 13753 12679 13787
rect 12621 13747 12679 13753
rect 12713 13787 12771 13793
rect 12713 13753 12725 13787
rect 12759 13753 12771 13787
rect 12713 13747 12771 13753
rect 12728 13716 12756 13747
rect 12820 13728 12848 13824
rect 13265 13821 13277 13824
rect 13311 13821 13323 13855
rect 13265 13815 13323 13821
rect 13354 13812 13360 13864
rect 13412 13812 13418 13864
rect 13998 13852 14004 13864
rect 13556 13824 14004 13852
rect 12929 13787 12987 13793
rect 12929 13753 12941 13787
rect 12975 13784 12987 13787
rect 13556 13784 13584 13824
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 12975 13756 13584 13784
rect 12975 13753 12987 13756
rect 12929 13747 12987 13753
rect 13630 13744 13636 13796
rect 13688 13744 13694 13796
rect 13722 13744 13728 13796
rect 13780 13784 13786 13796
rect 14093 13787 14151 13793
rect 14093 13784 14105 13787
rect 13780 13756 14105 13784
rect 13780 13744 13786 13756
rect 14093 13753 14105 13756
rect 14139 13753 14151 13787
rect 14093 13747 14151 13753
rect 14309 13787 14367 13793
rect 14309 13753 14321 13787
rect 14355 13784 14367 13787
rect 14927 13784 14955 13880
rect 15304 13839 15332 13880
rect 16114 13852 16120 13864
rect 15288 13833 15346 13839
rect 15288 13799 15300 13833
rect 15334 13799 15346 13833
rect 15810 13827 16120 13852
rect 15102 13793 15108 13796
rect 14355 13756 14955 13784
rect 14987 13787 15045 13793
rect 14355 13753 14367 13756
rect 14309 13747 14367 13753
rect 14987 13753 14999 13787
rect 15033 13753 15045 13787
rect 14987 13747 15045 13753
rect 15080 13787 15108 13793
rect 15080 13753 15092 13787
rect 15080 13747 15108 13753
rect 11900 13688 12756 13716
rect 12802 13676 12808 13728
rect 12860 13676 12866 13728
rect 13078 13676 13084 13728
rect 13136 13676 13142 13728
rect 13170 13676 13176 13728
rect 13228 13716 13234 13728
rect 13833 13719 13891 13725
rect 13833 13716 13845 13719
rect 13228 13688 13845 13716
rect 13228 13676 13234 13688
rect 13833 13685 13845 13688
rect 13879 13685 13891 13719
rect 13833 13679 13891 13685
rect 13998 13676 14004 13728
rect 14056 13676 14062 13728
rect 14461 13719 14519 13725
rect 14461 13685 14473 13719
rect 14507 13716 14519 13719
rect 14826 13716 14832 13728
rect 14507 13688 14832 13716
rect 14507 13685 14519 13688
rect 14461 13679 14519 13685
rect 14826 13676 14832 13688
rect 14884 13676 14890 13728
rect 15002 13716 15030 13747
rect 15102 13744 15108 13747
rect 15160 13744 15166 13796
rect 15194 13744 15200 13796
rect 15252 13744 15258 13796
rect 15288 13793 15346 13799
rect 15795 13824 16120 13827
rect 15795 13821 15853 13824
rect 15378 13744 15384 13796
rect 15436 13784 15442 13796
rect 15473 13787 15531 13793
rect 15473 13784 15485 13787
rect 15436 13756 15485 13784
rect 15436 13744 15442 13756
rect 15473 13753 15485 13756
rect 15519 13753 15531 13787
rect 15473 13747 15531 13753
rect 15562 13744 15568 13796
rect 15620 13744 15626 13796
rect 15795 13787 15807 13821
rect 15841 13787 15853 13821
rect 16114 13812 16120 13824
rect 16172 13812 16178 13864
rect 16758 13852 16764 13864
rect 16316 13824 16764 13852
rect 15795 13781 15853 13787
rect 15930 13744 15936 13796
rect 15988 13784 15994 13796
rect 16209 13787 16267 13793
rect 16209 13784 16221 13787
rect 15988 13756 16221 13784
rect 15988 13744 15994 13756
rect 16209 13753 16221 13756
rect 16255 13753 16267 13787
rect 16209 13747 16267 13753
rect 16316 13716 16344 13824
rect 16758 13812 16764 13824
rect 16816 13852 16822 13864
rect 17770 13852 17776 13864
rect 16816 13824 17776 13852
rect 16816 13812 16822 13824
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 19720 13861 19748 13892
rect 19705 13855 19763 13861
rect 18616 13824 18828 13852
rect 16666 13744 16672 13796
rect 16724 13784 16730 13796
rect 17497 13787 17555 13793
rect 17497 13784 17509 13787
rect 16724 13756 17509 13784
rect 16724 13744 16730 13756
rect 17497 13753 17509 13756
rect 17543 13753 17555 13787
rect 17497 13747 17555 13753
rect 18046 13744 18052 13796
rect 18104 13784 18110 13796
rect 18616 13784 18644 13824
rect 18104 13756 18644 13784
rect 18104 13744 18110 13756
rect 18690 13744 18696 13796
rect 18748 13744 18754 13796
rect 18800 13784 18828 13824
rect 19705 13821 19717 13855
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 19889 13855 19947 13861
rect 19889 13821 19901 13855
rect 19935 13852 19947 13855
rect 20438 13852 20444 13864
rect 19935 13824 20444 13852
rect 19935 13821 19947 13824
rect 19889 13815 19947 13821
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 20898 13852 20904 13864
rect 20732 13824 20904 13852
rect 20732 13818 20760 13824
rect 19794 13784 19800 13796
rect 18800 13756 19800 13784
rect 19794 13744 19800 13756
rect 19852 13744 19858 13796
rect 20346 13744 20352 13796
rect 20404 13744 20410 13796
rect 20641 13793 20760 13818
rect 20898 13812 20904 13824
rect 20956 13812 20962 13864
rect 20990 13812 20996 13864
rect 21048 13812 21054 13864
rect 21082 13812 21088 13864
rect 21140 13852 21146 13864
rect 21358 13852 21364 13864
rect 21140 13824 21364 13852
rect 21140 13812 21146 13824
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 21450 13812 21456 13864
rect 21508 13812 21514 13864
rect 21542 13812 21548 13864
rect 21600 13812 21606 13864
rect 21637 13855 21695 13861
rect 21637 13821 21649 13855
rect 21683 13821 21695 13855
rect 21637 13815 21695 13821
rect 20609 13790 20760 13793
rect 20609 13787 20669 13790
rect 20609 13753 20621 13787
rect 20655 13756 20669 13787
rect 20655 13753 20667 13756
rect 20609 13747 20667 13753
rect 20806 13744 20812 13796
rect 20864 13744 20870 13796
rect 21008 13784 21036 13812
rect 21560 13784 21588 13812
rect 21008 13756 21588 13784
rect 15002 13688 16344 13716
rect 16390 13676 16396 13728
rect 16448 13725 16454 13728
rect 16448 13719 16472 13725
rect 16460 13685 16472 13719
rect 16448 13679 16472 13685
rect 16577 13719 16635 13725
rect 16577 13685 16589 13719
rect 16623 13716 16635 13719
rect 16942 13716 16948 13728
rect 16623 13688 16948 13716
rect 16623 13685 16635 13688
rect 16577 13679 16635 13685
rect 16448 13676 16454 13679
rect 16942 13676 16948 13688
rect 17000 13676 17006 13728
rect 17126 13676 17132 13728
rect 17184 13676 17190 13728
rect 17310 13725 17316 13728
rect 17297 13719 17316 13725
rect 17297 13685 17309 13719
rect 17297 13679 17316 13685
rect 17310 13676 17316 13679
rect 17368 13676 17374 13728
rect 17586 13676 17592 13728
rect 17644 13716 17650 13728
rect 18782 13716 18788 13728
rect 17644 13688 18788 13716
rect 17644 13676 17650 13688
rect 18782 13676 18788 13688
rect 18840 13676 18846 13728
rect 18874 13676 18880 13728
rect 18932 13725 18938 13728
rect 18932 13719 18951 13725
rect 18939 13685 18951 13719
rect 18932 13679 18951 13685
rect 19153 13719 19211 13725
rect 19153 13685 19165 13719
rect 19199 13716 19211 13719
rect 19242 13716 19248 13728
rect 19199 13688 19248 13716
rect 19199 13685 19211 13688
rect 19153 13679 19211 13685
rect 18932 13676 18938 13679
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 20162 13725 20168 13728
rect 19981 13719 20039 13725
rect 19981 13716 19993 13719
rect 19392 13688 19993 13716
rect 19392 13676 19398 13688
rect 19981 13685 19993 13688
rect 20027 13685 20039 13719
rect 19981 13679 20039 13685
rect 20149 13719 20168 13725
rect 20149 13685 20161 13719
rect 20220 13716 20226 13728
rect 21008 13716 21036 13756
rect 20220 13688 21036 13716
rect 20149 13679 20168 13685
rect 20162 13676 20168 13679
rect 20220 13676 20226 13688
rect 21174 13676 21180 13728
rect 21232 13716 21238 13728
rect 21652 13716 21680 13815
rect 21726 13812 21732 13864
rect 21784 13812 21790 13864
rect 22462 13812 22468 13864
rect 22520 13852 22526 13864
rect 22741 13855 22799 13861
rect 22741 13852 22753 13855
rect 22520 13824 22753 13852
rect 22520 13812 22526 13824
rect 22741 13821 22753 13824
rect 22787 13821 22799 13855
rect 22741 13815 22799 13821
rect 23014 13812 23020 13864
rect 23072 13852 23078 13864
rect 23477 13855 23535 13861
rect 23477 13852 23489 13855
rect 23072 13824 23489 13852
rect 23072 13812 23078 13824
rect 23477 13821 23489 13824
rect 23523 13821 23535 13855
rect 23477 13815 23535 13821
rect 23566 13812 23572 13864
rect 23624 13852 23630 13864
rect 25705 13855 25763 13861
rect 23624 13827 24118 13852
rect 23624 13824 24133 13827
rect 23624 13812 23630 13824
rect 24075 13821 24133 13824
rect 21913 13787 21971 13793
rect 21913 13753 21925 13787
rect 21959 13784 21971 13787
rect 22002 13784 22008 13796
rect 21959 13756 22008 13784
rect 21959 13753 21971 13756
rect 21913 13747 21971 13753
rect 22002 13744 22008 13756
rect 22060 13744 22066 13796
rect 22554 13784 22560 13796
rect 22128 13756 22560 13784
rect 22128 13725 22156 13756
rect 22554 13744 22560 13756
rect 22612 13744 22618 13796
rect 23842 13744 23848 13796
rect 23900 13744 23906 13796
rect 24075 13787 24087 13821
rect 24121 13787 24133 13821
rect 25705 13821 25717 13855
rect 25751 13852 25763 13855
rect 25884 13852 25912 13892
rect 26602 13880 26608 13892
rect 26660 13880 26666 13932
rect 26804 13920 26832 14016
rect 27065 13991 27123 13997
rect 27065 13957 27077 13991
rect 27111 13988 27123 13991
rect 27111 13960 27384 13988
rect 27111 13957 27123 13960
rect 27065 13951 27123 13957
rect 27356 13929 27384 13960
rect 28074 13948 28080 14000
rect 28132 13988 28138 14000
rect 30944 13988 30972 14016
rect 28132 13960 30972 13988
rect 28132 13948 28138 13960
rect 27341 13923 27399 13929
rect 26804 13892 27292 13920
rect 25751 13824 25912 13852
rect 25751 13821 25763 13824
rect 25705 13815 25763 13821
rect 25958 13812 25964 13864
rect 26016 13812 26022 13864
rect 26053 13855 26111 13861
rect 26053 13821 26065 13855
rect 26099 13821 26111 13855
rect 26053 13815 26111 13821
rect 26145 13855 26203 13861
rect 26145 13821 26157 13855
rect 26191 13852 26203 13855
rect 26421 13855 26479 13861
rect 26421 13852 26433 13855
rect 26191 13824 26433 13852
rect 26191 13821 26203 13824
rect 26145 13815 26203 13821
rect 26421 13821 26433 13824
rect 26467 13821 26479 13855
rect 26421 13815 26479 13821
rect 24075 13781 24133 13787
rect 22118 13719 22176 13725
rect 22118 13716 22130 13719
rect 21232 13688 22130 13716
rect 21232 13676 21238 13688
rect 22118 13685 22130 13688
rect 22164 13685 22176 13719
rect 22118 13679 22176 13685
rect 22278 13676 22284 13728
rect 22336 13676 22342 13728
rect 22370 13676 22376 13728
rect 22428 13716 22434 13728
rect 23198 13716 23204 13728
rect 22428 13688 23204 13716
rect 22428 13676 22434 13688
rect 23198 13676 23204 13688
rect 23256 13676 23262 13728
rect 23382 13676 23388 13728
rect 23440 13676 23446 13728
rect 24210 13676 24216 13728
rect 24268 13676 24274 13728
rect 25038 13676 25044 13728
rect 25096 13716 25102 13728
rect 26068 13716 26096 13815
rect 26436 13784 26464 13815
rect 26510 13812 26516 13864
rect 26568 13852 26574 13864
rect 27264 13861 27292 13892
rect 27341 13889 27353 13923
rect 27387 13920 27399 13923
rect 27798 13920 27804 13932
rect 27387 13892 27804 13920
rect 27387 13889 27399 13892
rect 27341 13883 27399 13889
rect 27798 13880 27804 13892
rect 27856 13920 27862 13932
rect 29178 13920 29184 13932
rect 27856 13892 28028 13920
rect 27856 13880 27862 13892
rect 28000 13861 28028 13892
rect 29012 13892 29184 13920
rect 29012 13861 29040 13892
rect 29178 13880 29184 13892
rect 29236 13880 29242 13932
rect 26697 13855 26755 13861
rect 26697 13852 26709 13855
rect 26568 13824 26709 13852
rect 26568 13812 26574 13824
rect 26697 13821 26709 13824
rect 26743 13821 26755 13855
rect 26697 13815 26755 13821
rect 26973 13855 27031 13861
rect 26973 13821 26985 13855
rect 27019 13821 27031 13855
rect 26973 13815 27031 13821
rect 27249 13855 27307 13861
rect 27249 13821 27261 13855
rect 27295 13821 27307 13855
rect 27249 13815 27307 13821
rect 27525 13855 27583 13861
rect 27525 13821 27537 13855
rect 27571 13821 27583 13855
rect 27525 13815 27583 13821
rect 27985 13855 28043 13861
rect 27985 13821 27997 13855
rect 28031 13821 28043 13855
rect 27985 13815 28043 13821
rect 28997 13855 29055 13861
rect 28997 13821 29009 13855
rect 29043 13821 29055 13855
rect 28997 13815 29055 13821
rect 26786 13784 26792 13796
rect 26436 13756 26792 13784
rect 26786 13744 26792 13756
rect 26844 13784 26850 13796
rect 26988 13784 27016 13815
rect 26844 13756 27016 13784
rect 26844 13744 26850 13756
rect 25096 13688 26096 13716
rect 26513 13719 26571 13725
rect 25096 13676 25102 13688
rect 26513 13685 26525 13719
rect 26559 13716 26571 13719
rect 26602 13716 26608 13728
rect 26559 13688 26608 13716
rect 26559 13685 26571 13688
rect 26513 13679 26571 13685
rect 26602 13676 26608 13688
rect 26660 13716 26666 13728
rect 27540 13716 27568 13815
rect 28000 13784 28028 13815
rect 29270 13812 29276 13864
rect 29328 13852 29334 13864
rect 29457 13855 29515 13861
rect 29457 13852 29469 13855
rect 29328 13824 29469 13852
rect 29328 13812 29334 13824
rect 29457 13821 29469 13824
rect 29503 13821 29515 13855
rect 29457 13815 29515 13821
rect 28074 13784 28080 13796
rect 28000 13756 28080 13784
rect 28074 13744 28080 13756
rect 28132 13744 28138 13796
rect 26660 13688 27568 13716
rect 29089 13719 29147 13725
rect 26660 13676 26666 13688
rect 29089 13685 29101 13719
rect 29135 13716 29147 13719
rect 29454 13716 29460 13728
rect 29135 13688 29460 13716
rect 29135 13685 29147 13688
rect 29089 13679 29147 13685
rect 29454 13676 29460 13688
rect 29512 13676 29518 13728
rect 552 13626 31531 13648
rect 552 13574 8102 13626
rect 8154 13574 8166 13626
rect 8218 13574 8230 13626
rect 8282 13574 8294 13626
rect 8346 13574 8358 13626
rect 8410 13574 15807 13626
rect 15859 13574 15871 13626
rect 15923 13574 15935 13626
rect 15987 13574 15999 13626
rect 16051 13574 16063 13626
rect 16115 13574 23512 13626
rect 23564 13574 23576 13626
rect 23628 13574 23640 13626
rect 23692 13574 23704 13626
rect 23756 13574 23768 13626
rect 23820 13574 31217 13626
rect 31269 13574 31281 13626
rect 31333 13574 31345 13626
rect 31397 13574 31409 13626
rect 31461 13574 31473 13626
rect 31525 13574 31531 13626
rect 552 13552 31531 13574
rect 1121 13515 1179 13521
rect 1121 13481 1133 13515
rect 1167 13512 1179 13515
rect 1210 13512 1216 13524
rect 1167 13484 1216 13512
rect 1167 13481 1179 13484
rect 1121 13475 1179 13481
rect 1210 13472 1216 13484
rect 1268 13472 1274 13524
rect 4065 13515 4123 13521
rect 4065 13481 4077 13515
rect 4111 13512 4123 13515
rect 4154 13512 4160 13524
rect 4111 13484 4160 13512
rect 4111 13481 4123 13484
rect 4065 13475 4123 13481
rect 4154 13472 4160 13484
rect 4212 13512 4218 13524
rect 4706 13512 4712 13524
rect 4212 13484 4712 13512
rect 4212 13472 4218 13484
rect 4706 13472 4712 13484
rect 4764 13512 4770 13524
rect 4893 13515 4951 13521
rect 4893 13512 4905 13515
rect 4764 13484 4905 13512
rect 4764 13472 4770 13484
rect 4893 13481 4905 13484
rect 4939 13481 4951 13515
rect 4893 13475 4951 13481
rect 5166 13472 5172 13524
rect 5224 13472 5230 13524
rect 8018 13472 8024 13524
rect 8076 13472 8082 13524
rect 9858 13472 9864 13524
rect 9916 13472 9922 13524
rect 10134 13472 10140 13524
rect 10192 13472 10198 13524
rect 11606 13472 11612 13524
rect 11664 13472 11670 13524
rect 12342 13512 12348 13524
rect 11716 13484 12348 13512
rect 1029 13379 1087 13385
rect 1029 13345 1041 13379
rect 1075 13345 1087 13379
rect 1228 13376 1256 13472
rect 1394 13404 1400 13456
rect 1452 13404 1458 13456
rect 8036 13444 8064 13472
rect 8113 13447 8171 13453
rect 8113 13444 8125 13447
rect 4448 13416 5028 13444
rect 1305 13379 1363 13385
rect 1305 13376 1317 13379
rect 1228 13348 1317 13376
rect 1029 13339 1087 13345
rect 1305 13345 1317 13348
rect 1351 13345 1363 13379
rect 1305 13339 1363 13345
rect 1044 13308 1072 13339
rect 1412 13308 1440 13404
rect 1762 13336 1768 13388
rect 1820 13376 1826 13388
rect 4448 13385 4476 13416
rect 5000 13388 5028 13416
rect 5828 13416 8125 13444
rect 1929 13379 1987 13385
rect 1929 13376 1941 13379
rect 1820 13348 1941 13376
rect 1820 13336 1826 13348
rect 1929 13345 1941 13348
rect 1975 13345 1987 13379
rect 1929 13339 1987 13345
rect 4157 13379 4215 13385
rect 4157 13345 4169 13379
rect 4203 13345 4215 13379
rect 4157 13339 4215 13345
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13345 4491 13379
rect 4433 13339 4491 13345
rect 4525 13379 4583 13385
rect 4525 13345 4537 13379
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 1044 13280 1440 13308
rect 1670 13268 1676 13320
rect 1728 13268 1734 13320
rect 4172 13308 4200 13339
rect 4540 13308 4568 13339
rect 4798 13336 4804 13388
rect 4856 13336 4862 13388
rect 4982 13336 4988 13388
rect 5040 13376 5046 13388
rect 5828 13385 5856 13416
rect 8113 13413 8125 13416
rect 8159 13413 8171 13447
rect 8113 13407 8171 13413
rect 9324 13416 9996 13444
rect 5077 13379 5135 13385
rect 5077 13376 5089 13379
rect 5040 13348 5089 13376
rect 5040 13336 5046 13348
rect 5077 13345 5089 13348
rect 5123 13345 5135 13379
rect 5077 13339 5135 13345
rect 5813 13379 5871 13385
rect 5813 13345 5825 13379
rect 5859 13345 5871 13379
rect 6069 13379 6127 13385
rect 6069 13376 6081 13379
rect 5813 13339 5871 13345
rect 5920 13348 6081 13376
rect 4172 13280 4568 13308
rect 4617 13311 4675 13317
rect 3050 13200 3056 13252
rect 3108 13200 3114 13252
rect 4172 13184 4200 13280
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 5442 13308 5448 13320
rect 4663 13280 5448 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 5442 13268 5448 13280
rect 5500 13308 5506 13320
rect 5920 13308 5948 13348
rect 6069 13345 6081 13348
rect 6115 13345 6127 13379
rect 6069 13339 6127 13345
rect 7285 13379 7343 13385
rect 7285 13345 7297 13379
rect 7331 13345 7343 13379
rect 7285 13339 7343 13345
rect 5500 13280 5948 13308
rect 5500 13268 5506 13280
rect 7300 13252 7328 13339
rect 7558 13336 7564 13388
rect 7616 13376 7622 13388
rect 8478 13376 8484 13388
rect 7616 13348 8484 13376
rect 7616 13336 7622 13348
rect 8478 13336 8484 13348
rect 8536 13336 8542 13388
rect 9324 13320 9352 13416
rect 9968 13385 9996 13416
rect 11624 13385 11652 13472
rect 11716 13453 11744 13484
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 13909 13515 13967 13521
rect 13909 13481 13921 13515
rect 13955 13512 13967 13515
rect 16574 13512 16580 13524
rect 13955 13484 16580 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 16758 13472 16764 13524
rect 16816 13472 16822 13524
rect 16850 13472 16856 13524
rect 16908 13512 16914 13524
rect 22830 13512 22836 13524
rect 16908 13484 17724 13512
rect 16908 13472 16914 13484
rect 11701 13447 11759 13453
rect 11701 13413 11713 13447
rect 11747 13413 11759 13447
rect 11701 13407 11759 13413
rect 11917 13447 11975 13453
rect 11917 13413 11929 13447
rect 11963 13444 11975 13447
rect 12986 13444 12992 13456
rect 11963 13416 12992 13444
rect 11963 13413 11975 13416
rect 11917 13407 11975 13413
rect 12986 13404 12992 13416
rect 13044 13404 13050 13456
rect 13630 13444 13636 13456
rect 13188 13416 13636 13444
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 9953 13379 10011 13385
rect 9953 13345 9965 13379
rect 9999 13376 10011 13379
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9999 13348 10057 13376
rect 9999 13345 10011 13348
rect 9953 13339 10011 13345
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 11609 13379 11667 13385
rect 11609 13345 11621 13379
rect 11655 13345 11667 13379
rect 12158 13376 12164 13388
rect 11609 13339 11667 13345
rect 11992 13348 12164 13376
rect 7650 13268 7656 13320
rect 7708 13308 7714 13320
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 7708 13280 8401 13308
rect 7708 13268 7714 13280
rect 8389 13277 8401 13280
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 9306 13268 9312 13320
rect 9364 13268 9370 13320
rect 9692 13308 9720 13339
rect 9766 13308 9772 13320
rect 9692 13280 9772 13308
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 11992 13308 12020 13348
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 13188 13385 13216 13416
rect 13630 13404 13636 13416
rect 13688 13444 13694 13456
rect 13688 13416 14044 13444
rect 13688 13404 13694 13416
rect 13173 13379 13231 13385
rect 13173 13345 13185 13379
rect 13219 13345 13231 13379
rect 13173 13339 13231 13345
rect 13357 13379 13415 13385
rect 13357 13345 13369 13379
rect 13403 13376 13415 13379
rect 13722 13376 13728 13388
rect 13403 13348 13728 13376
rect 13403 13345 13415 13348
rect 13357 13339 13415 13345
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14016 13376 14044 13416
rect 14200 13416 14955 13444
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 14016 13348 14105 13376
rect 14093 13345 14105 13348
rect 14139 13345 14151 13379
rect 14093 13339 14151 13345
rect 11532 13280 12020 13308
rect 7282 13200 7288 13252
rect 7340 13240 7346 13252
rect 11532 13240 11560 13280
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 12989 13311 13047 13317
rect 12989 13308 13001 13311
rect 12124 13280 13001 13308
rect 12124 13268 12130 13280
rect 12989 13277 13001 13280
rect 13035 13308 13047 13311
rect 13035 13280 14136 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 14108 13252 14136 13280
rect 12802 13240 12808 13252
rect 7340 13212 11560 13240
rect 11624 13212 12808 13240
rect 7340 13200 7346 13212
rect 11624 13184 11652 13212
rect 12802 13200 12808 13212
rect 12860 13200 12866 13252
rect 13078 13200 13084 13252
rect 13136 13240 13142 13252
rect 13541 13243 13599 13249
rect 13541 13240 13553 13243
rect 13136 13212 13553 13240
rect 13136 13200 13142 13212
rect 13541 13209 13553 13212
rect 13587 13209 13599 13243
rect 13541 13203 13599 13209
rect 14090 13200 14096 13252
rect 14148 13200 14154 13252
rect 1118 13132 1124 13184
rect 1176 13172 1182 13184
rect 1397 13175 1455 13181
rect 1397 13172 1409 13175
rect 1176 13144 1409 13172
rect 1176 13132 1182 13144
rect 1397 13141 1409 13144
rect 1443 13141 1455 13175
rect 1397 13135 1455 13141
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 4212 13144 4353 13172
rect 4212 13132 4218 13144
rect 4341 13141 4353 13144
rect 4387 13141 4399 13175
rect 4341 13135 4399 13141
rect 7193 13175 7251 13181
rect 7193 13141 7205 13175
rect 7239 13172 7251 13175
rect 7558 13172 7564 13184
rect 7239 13144 7564 13172
rect 7239 13141 7251 13144
rect 7193 13135 7251 13141
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 9306 13132 9312 13184
rect 9364 13172 9370 13184
rect 9585 13175 9643 13181
rect 9585 13172 9597 13175
rect 9364 13144 9597 13172
rect 9364 13132 9370 13144
rect 9585 13141 9597 13144
rect 9631 13141 9643 13175
rect 9585 13135 9643 13141
rect 11517 13175 11575 13181
rect 11517 13141 11529 13175
rect 11563 13172 11575 13175
rect 11606 13172 11612 13184
rect 11563 13144 11612 13172
rect 11563 13141 11575 13144
rect 11517 13135 11575 13141
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 11790 13132 11796 13184
rect 11848 13172 11854 13184
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11848 13144 11897 13172
rect 11848 13132 11854 13144
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 11885 13135 11943 13141
rect 12069 13175 12127 13181
rect 12069 13141 12081 13175
rect 12115 13172 12127 13175
rect 13449 13175 13507 13181
rect 13449 13172 13461 13175
rect 12115 13144 13461 13172
rect 12115 13141 12127 13144
rect 12069 13135 12127 13141
rect 13449 13141 13461 13144
rect 13495 13141 13507 13175
rect 13449 13135 13507 13141
rect 13633 13175 13691 13181
rect 13633 13141 13645 13175
rect 13679 13172 13691 13175
rect 14200 13172 14228 13416
rect 14274 13336 14280 13388
rect 14332 13336 14338 13388
rect 14366 13336 14372 13388
rect 14424 13336 14430 13388
rect 14553 13379 14611 13385
rect 14826 13382 14832 13388
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 14752 13376 14832 13382
rect 14599 13354 14832 13376
rect 14599 13348 14780 13354
rect 14824 13348 14832 13354
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 14927 13376 14955 13416
rect 15378 13404 15384 13456
rect 15436 13444 15442 13456
rect 15436 13416 17632 13444
rect 15436 13404 15442 13416
rect 14927 13348 15700 13376
rect 14384 13308 14412 13336
rect 15672 13308 15700 13348
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 16669 13379 16727 13385
rect 16669 13376 16681 13379
rect 15804 13348 16681 13376
rect 15804 13336 15810 13348
rect 16669 13345 16681 13348
rect 16715 13345 16727 13379
rect 16669 13339 16727 13345
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 16945 13379 17003 13385
rect 16945 13376 16957 13379
rect 16908 13348 16957 13376
rect 16908 13336 16914 13348
rect 16945 13345 16957 13348
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 17037 13379 17095 13385
rect 17037 13345 17049 13379
rect 17083 13376 17095 13379
rect 17126 13376 17132 13388
rect 17083 13348 17132 13376
rect 17083 13345 17095 13348
rect 17037 13339 17095 13345
rect 17126 13336 17132 13348
rect 17184 13336 17190 13388
rect 17604 13385 17632 13416
rect 17696 13385 17724 13484
rect 17972 13484 22836 13512
rect 17770 13404 17776 13456
rect 17828 13444 17834 13456
rect 17972 13453 18000 13484
rect 22830 13472 22836 13484
rect 22888 13472 22894 13524
rect 23382 13472 23388 13524
rect 23440 13512 23446 13524
rect 23477 13515 23535 13521
rect 23477 13512 23489 13515
rect 23440 13484 23489 13512
rect 23440 13472 23446 13484
rect 23477 13481 23489 13484
rect 23523 13481 23535 13515
rect 23477 13475 23535 13481
rect 24581 13515 24639 13521
rect 24581 13481 24593 13515
rect 24627 13512 24639 13515
rect 24857 13515 24915 13521
rect 24857 13512 24869 13515
rect 24627 13484 24869 13512
rect 24627 13481 24639 13484
rect 24581 13475 24639 13481
rect 24857 13481 24869 13484
rect 24903 13512 24915 13515
rect 26513 13515 26571 13521
rect 24903 13484 26464 13512
rect 24903 13481 24915 13484
rect 24857 13475 24915 13481
rect 17865 13447 17923 13453
rect 17865 13444 17877 13447
rect 17828 13416 17877 13444
rect 17828 13404 17834 13416
rect 17865 13413 17877 13416
rect 17911 13413 17923 13447
rect 17865 13407 17923 13413
rect 17957 13447 18015 13453
rect 17957 13413 17969 13447
rect 18003 13413 18015 13447
rect 17957 13407 18015 13413
rect 18322 13404 18328 13456
rect 18380 13444 18386 13456
rect 18874 13444 18880 13456
rect 18380 13416 18880 13444
rect 18380 13404 18386 13416
rect 18874 13404 18880 13416
rect 18932 13453 18938 13456
rect 18932 13447 18995 13453
rect 18932 13413 18949 13447
rect 18983 13413 18995 13447
rect 18932 13407 18995 13413
rect 18932 13404 18938 13407
rect 19150 13404 19156 13456
rect 19208 13404 19214 13456
rect 19797 13447 19855 13453
rect 19797 13413 19809 13447
rect 19843 13444 19855 13447
rect 21634 13444 21640 13456
rect 19843 13416 21640 13444
rect 19843 13413 19855 13416
rect 19797 13407 19855 13413
rect 17589 13379 17647 13385
rect 17589 13345 17601 13379
rect 17635 13345 17647 13379
rect 17589 13339 17647 13345
rect 17682 13379 17740 13385
rect 17682 13345 17694 13379
rect 17728 13345 17740 13379
rect 17682 13339 17740 13345
rect 18046 13336 18052 13388
rect 18104 13385 18110 13388
rect 18104 13376 18112 13385
rect 18598 13376 18604 13388
rect 18104 13348 18604 13376
rect 18104 13339 18112 13348
rect 18104 13336 18110 13339
rect 18598 13336 18604 13348
rect 18656 13336 18662 13388
rect 19334 13376 19340 13388
rect 18892 13348 19340 13376
rect 14384 13280 14504 13308
rect 15672 13280 18828 13308
rect 14476 13249 14504 13280
rect 18800 13249 18828 13280
rect 14461 13243 14519 13249
rect 14461 13209 14473 13243
rect 14507 13209 14519 13243
rect 18785 13243 18843 13249
rect 14461 13203 14519 13209
rect 14768 13212 18368 13240
rect 13679 13144 14228 13172
rect 14369 13175 14427 13181
rect 13679 13141 13691 13144
rect 13633 13135 13691 13141
rect 14369 13141 14381 13175
rect 14415 13172 14427 13175
rect 14768 13172 14796 13212
rect 14415 13144 14796 13172
rect 14415 13141 14427 13144
rect 14369 13135 14427 13141
rect 14826 13132 14832 13184
rect 14884 13132 14890 13184
rect 15194 13132 15200 13184
rect 15252 13172 15258 13184
rect 15470 13172 15476 13184
rect 15252 13144 15476 13172
rect 15252 13132 15258 13144
rect 15470 13132 15476 13144
rect 15528 13172 15534 13184
rect 16390 13172 16396 13184
rect 15528 13144 16396 13172
rect 15528 13132 15534 13144
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 16850 13132 16856 13184
rect 16908 13172 16914 13184
rect 17129 13175 17187 13181
rect 17129 13172 17141 13175
rect 16908 13144 17141 13172
rect 16908 13132 16914 13144
rect 17129 13141 17141 13144
rect 17175 13141 17187 13175
rect 17129 13135 17187 13141
rect 17218 13132 17224 13184
rect 17276 13172 17282 13184
rect 17405 13175 17463 13181
rect 17405 13172 17417 13175
rect 17276 13144 17417 13172
rect 17276 13132 17282 13144
rect 17405 13141 17417 13144
rect 17451 13141 17463 13175
rect 17405 13135 17463 13141
rect 17586 13132 17592 13184
rect 17644 13172 17650 13184
rect 18046 13172 18052 13184
rect 17644 13144 18052 13172
rect 17644 13132 17650 13144
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 18230 13132 18236 13184
rect 18288 13132 18294 13184
rect 18340 13172 18368 13212
rect 18785 13209 18797 13243
rect 18831 13209 18843 13243
rect 18785 13203 18843 13209
rect 18892 13172 18920 13348
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 20162 13376 20168 13388
rect 19484 13348 20168 13376
rect 19484 13336 19490 13348
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 19245 13311 19303 13317
rect 19245 13277 19257 13311
rect 19291 13308 19303 13311
rect 20070 13308 20076 13320
rect 19291 13280 20076 13308
rect 19291 13277 19303 13280
rect 19245 13271 19303 13277
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 20456 13308 20484 13416
rect 21634 13404 21640 13416
rect 21692 13444 21698 13456
rect 21692 13416 25176 13444
rect 21692 13404 21698 13416
rect 20530 13336 20536 13388
rect 20588 13376 20594 13388
rect 21174 13376 21180 13388
rect 20588 13348 21180 13376
rect 20588 13336 20594 13348
rect 21174 13336 21180 13348
rect 21232 13336 21238 13388
rect 21453 13379 21511 13385
rect 21453 13345 21465 13379
rect 21499 13376 21511 13379
rect 21542 13376 21548 13388
rect 21499 13348 21548 13376
rect 21499 13345 21511 13348
rect 21453 13339 21511 13345
rect 21542 13336 21548 13348
rect 21600 13336 21606 13388
rect 21818 13336 21824 13388
rect 21876 13376 21882 13388
rect 22186 13376 22192 13388
rect 21876 13348 22192 13376
rect 21876 13336 21882 13348
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 22364 13379 22422 13385
rect 22364 13345 22376 13379
rect 22410 13376 22422 13379
rect 24394 13376 24400 13388
rect 22410 13348 24400 13376
rect 22410 13345 22422 13348
rect 23011 13346 23060 13348
rect 22364 13339 22422 13345
rect 24394 13336 24400 13348
rect 24452 13376 24458 13388
rect 24489 13379 24547 13385
rect 24489 13376 24501 13379
rect 24452 13348 24501 13376
rect 24452 13336 24458 13348
rect 24489 13345 24501 13348
rect 24535 13345 24547 13379
rect 24489 13339 24547 13345
rect 24949 13379 25007 13385
rect 24949 13345 24961 13379
rect 24995 13376 25007 13379
rect 25038 13376 25044 13388
rect 24995 13348 25044 13376
rect 24995 13345 25007 13348
rect 24949 13339 25007 13345
rect 25038 13336 25044 13348
rect 25096 13336 25102 13388
rect 20456 13280 20576 13308
rect 20548 13252 20576 13280
rect 19150 13200 19156 13252
rect 19208 13240 19214 13252
rect 19613 13243 19671 13249
rect 19613 13240 19625 13243
rect 19208 13212 19625 13240
rect 19208 13200 19214 13212
rect 19613 13209 19625 13212
rect 19659 13209 19671 13243
rect 19613 13203 19671 13209
rect 20530 13200 20536 13252
rect 20588 13200 20594 13252
rect 21192 13240 21220 13336
rect 21269 13311 21327 13317
rect 21269 13277 21281 13311
rect 21315 13308 21327 13311
rect 21358 13308 21364 13320
rect 21315 13280 21364 13308
rect 21315 13277 21327 13280
rect 21269 13271 21327 13277
rect 21358 13268 21364 13280
rect 21416 13308 21422 13320
rect 21726 13308 21732 13320
rect 21416 13280 21732 13308
rect 21416 13268 21422 13280
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 22097 13311 22155 13317
rect 22097 13277 22109 13311
rect 22143 13277 22155 13311
rect 22097 13271 22155 13277
rect 22112 13240 22140 13271
rect 23474 13268 23480 13320
rect 23532 13308 23538 13320
rect 24578 13308 24584 13320
rect 23532 13280 24584 13308
rect 23532 13268 23538 13280
rect 24578 13268 24584 13280
rect 24636 13268 24642 13320
rect 25148 13308 25176 13416
rect 25240 13385 25268 13484
rect 26436 13385 26464 13484
rect 26513 13481 26525 13515
rect 26559 13512 26571 13515
rect 26602 13512 26608 13524
rect 26559 13484 26608 13512
rect 26559 13481 26571 13484
rect 26513 13475 26571 13481
rect 26602 13472 26608 13484
rect 26660 13472 26666 13524
rect 26786 13472 26792 13524
rect 26844 13472 26850 13524
rect 27706 13472 27712 13524
rect 27764 13512 27770 13524
rect 28445 13515 28503 13521
rect 28445 13512 28457 13515
rect 27764 13484 28457 13512
rect 27764 13472 27770 13484
rect 28445 13481 28457 13484
rect 28491 13481 28503 13515
rect 28445 13475 28503 13481
rect 28074 13404 28080 13456
rect 28132 13453 28138 13456
rect 28132 13407 28144 13453
rect 28132 13404 28138 13407
rect 29270 13404 29276 13456
rect 29328 13444 29334 13456
rect 29558 13447 29616 13453
rect 29558 13444 29570 13447
rect 29328 13416 29570 13444
rect 29328 13404 29334 13416
rect 29558 13413 29570 13416
rect 29604 13413 29616 13447
rect 29558 13407 29616 13413
rect 25225 13379 25283 13385
rect 25225 13345 25237 13379
rect 25271 13345 25283 13379
rect 25225 13339 25283 13345
rect 25317 13379 25375 13385
rect 25317 13345 25329 13379
rect 25363 13345 25375 13379
rect 25317 13339 25375 13345
rect 26421 13379 26479 13385
rect 26421 13345 26433 13379
rect 26467 13345 26479 13379
rect 26421 13339 26479 13345
rect 25332 13308 25360 13339
rect 26510 13336 26516 13388
rect 26568 13376 26574 13388
rect 26697 13379 26755 13385
rect 26697 13376 26709 13379
rect 26568 13348 26709 13376
rect 26568 13336 26574 13348
rect 26697 13345 26709 13348
rect 26743 13345 26755 13379
rect 28353 13379 28411 13385
rect 28353 13376 28365 13379
rect 26697 13339 26755 13345
rect 26804 13348 28365 13376
rect 25406 13308 25412 13320
rect 25148 13280 25412 13308
rect 25406 13268 25412 13280
rect 25464 13268 25470 13320
rect 25682 13268 25688 13320
rect 25740 13308 25746 13320
rect 25958 13308 25964 13320
rect 25740 13280 25964 13308
rect 25740 13268 25746 13280
rect 25958 13268 25964 13280
rect 26016 13308 26022 13320
rect 26053 13311 26111 13317
rect 26053 13308 26065 13311
rect 26016 13280 26065 13308
rect 26016 13268 26022 13280
rect 26053 13277 26065 13280
rect 26099 13308 26111 13311
rect 26804 13308 26832 13348
rect 28353 13345 28365 13348
rect 28399 13345 28411 13379
rect 28353 13339 28411 13345
rect 26099 13280 26832 13308
rect 29825 13311 29883 13317
rect 26099 13277 26111 13280
rect 26053 13271 26111 13277
rect 29825 13277 29837 13311
rect 29871 13277 29883 13311
rect 29825 13271 29883 13277
rect 21192 13212 22140 13240
rect 23290 13200 23296 13252
rect 23348 13240 23354 13252
rect 23348 13212 25268 13240
rect 23348 13200 23354 13212
rect 18340 13144 18920 13172
rect 18969 13175 19027 13181
rect 18969 13141 18981 13175
rect 19015 13172 19027 13175
rect 19058 13172 19064 13184
rect 19015 13144 19064 13172
rect 19015 13141 19027 13144
rect 18969 13135 19027 13141
rect 19058 13132 19064 13144
rect 19116 13172 19122 13184
rect 19426 13172 19432 13184
rect 19116 13144 19432 13172
rect 19116 13132 19122 13144
rect 19426 13132 19432 13144
rect 19484 13132 19490 13184
rect 20438 13132 20444 13184
rect 20496 13172 20502 13184
rect 21634 13172 21640 13184
rect 20496 13144 21640 13172
rect 20496 13132 20502 13144
rect 21634 13132 21640 13144
rect 21692 13132 21698 13184
rect 25038 13132 25044 13184
rect 25096 13172 25102 13184
rect 25133 13175 25191 13181
rect 25133 13172 25145 13175
rect 25096 13144 25145 13172
rect 25096 13132 25102 13144
rect 25133 13141 25145 13144
rect 25179 13141 25191 13175
rect 25240 13172 25268 13212
rect 26973 13175 27031 13181
rect 26973 13172 26985 13175
rect 25240 13144 26985 13172
rect 25133 13135 25191 13141
rect 26973 13141 26985 13144
rect 27019 13141 27031 13175
rect 26973 13135 27031 13141
rect 29086 13132 29092 13184
rect 29144 13172 29150 13184
rect 29840 13172 29868 13271
rect 29144 13144 29868 13172
rect 29144 13132 29150 13144
rect 552 13082 31372 13104
rect 552 13030 4250 13082
rect 4302 13030 4314 13082
rect 4366 13030 4378 13082
rect 4430 13030 4442 13082
rect 4494 13030 4506 13082
rect 4558 13030 11955 13082
rect 12007 13030 12019 13082
rect 12071 13030 12083 13082
rect 12135 13030 12147 13082
rect 12199 13030 12211 13082
rect 12263 13030 19660 13082
rect 19712 13030 19724 13082
rect 19776 13030 19788 13082
rect 19840 13030 19852 13082
rect 19904 13030 19916 13082
rect 19968 13030 27365 13082
rect 27417 13030 27429 13082
rect 27481 13030 27493 13082
rect 27545 13030 27557 13082
rect 27609 13030 27621 13082
rect 27673 13030 31372 13082
rect 552 13008 31372 13030
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 4433 12971 4491 12977
rect 4433 12968 4445 12971
rect 4212 12940 4445 12968
rect 4212 12928 4218 12940
rect 4433 12937 4445 12940
rect 4479 12937 4491 12971
rect 4433 12931 4491 12937
rect 7282 12928 7288 12980
rect 7340 12928 7346 12980
rect 7466 12928 7472 12980
rect 7524 12928 7530 12980
rect 9306 12928 9312 12980
rect 9364 12928 9370 12980
rect 10042 12968 10048 12980
rect 9876 12940 10048 12968
rect 4798 12832 4804 12844
rect 4632 12804 4804 12832
rect 1029 12767 1087 12773
rect 1029 12733 1041 12767
rect 1075 12733 1087 12767
rect 1029 12727 1087 12733
rect 1121 12767 1179 12773
rect 1121 12733 1133 12767
rect 1167 12764 1179 12767
rect 1302 12764 1308 12776
rect 1167 12736 1308 12764
rect 1167 12733 1179 12736
rect 1121 12727 1179 12733
rect 1044 12696 1072 12727
rect 1302 12724 1308 12736
rect 1360 12724 1366 12776
rect 1394 12724 1400 12776
rect 1452 12724 1458 12776
rect 1670 12724 1676 12776
rect 1728 12724 1734 12776
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 4632 12773 4660 12804
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 4249 12767 4307 12773
rect 4249 12764 4261 12767
rect 4212 12736 4261 12764
rect 4212 12724 4218 12736
rect 4249 12733 4261 12736
rect 4295 12764 4307 12767
rect 4341 12767 4399 12773
rect 4341 12764 4353 12767
rect 4295 12736 4353 12764
rect 4295 12733 4307 12736
rect 4249 12727 4307 12733
rect 4341 12733 4353 12736
rect 4387 12733 4399 12767
rect 4341 12727 4399 12733
rect 4617 12767 4675 12773
rect 4617 12733 4629 12767
rect 4663 12733 4675 12767
rect 4617 12727 4675 12733
rect 1412 12696 1440 12724
rect 1918 12699 1976 12705
rect 1918 12696 1930 12699
rect 1044 12668 1930 12696
rect 1918 12665 1930 12668
rect 1964 12665 1976 12699
rect 1918 12659 1976 12665
rect 1118 12588 1124 12640
rect 1176 12628 1182 12640
rect 1397 12631 1455 12637
rect 1397 12628 1409 12631
rect 1176 12600 1409 12628
rect 1176 12588 1182 12600
rect 1397 12597 1409 12600
rect 1443 12597 1455 12631
rect 1397 12591 1455 12597
rect 3050 12588 3056 12640
rect 3108 12588 3114 12640
rect 4157 12631 4215 12637
rect 4157 12597 4169 12631
rect 4203 12628 4215 12631
rect 4246 12628 4252 12640
rect 4203 12600 4252 12628
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 4246 12588 4252 12600
rect 4304 12628 4310 12640
rect 4632 12628 4660 12727
rect 6086 12724 6092 12776
rect 6144 12724 6150 12776
rect 6181 12767 6239 12773
rect 6181 12733 6193 12767
rect 6227 12733 6239 12767
rect 6181 12727 6239 12733
rect 6457 12767 6515 12773
rect 6457 12733 6469 12767
rect 6503 12764 6515 12767
rect 7300 12764 7328 12928
rect 7484 12832 7512 12928
rect 7926 12832 7932 12844
rect 7484 12804 7932 12832
rect 7926 12792 7932 12804
rect 7984 12832 7990 12844
rect 9876 12841 9904 12940
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11848 12940 11989 12968
rect 11848 12928 11854 12940
rect 11977 12937 11989 12940
rect 12023 12968 12035 12971
rect 13170 12968 13176 12980
rect 12023 12940 13176 12968
rect 12023 12937 12035 12940
rect 11977 12931 12035 12937
rect 13170 12928 13176 12940
rect 13228 12928 13234 12980
rect 13998 12928 14004 12980
rect 14056 12928 14062 12980
rect 14182 12928 14188 12980
rect 14240 12928 14246 12980
rect 14277 12971 14335 12977
rect 14277 12937 14289 12971
rect 14323 12968 14335 12971
rect 16482 12968 16488 12980
rect 14323 12940 16488 12968
rect 14323 12937 14335 12940
rect 14277 12931 14335 12937
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 16666 12968 16672 12980
rect 16724 12977 16730 12980
rect 16724 12971 16749 12977
rect 16592 12940 16672 12968
rect 13357 12903 13415 12909
rect 13357 12869 13369 12903
rect 13403 12900 13415 12903
rect 13817 12903 13875 12909
rect 13817 12900 13829 12903
rect 13403 12872 13829 12900
rect 13403 12869 13415 12872
rect 13357 12863 13415 12869
rect 13817 12869 13829 12872
rect 13863 12869 13875 12903
rect 13817 12863 13875 12869
rect 9861 12835 9919 12841
rect 7984 12804 8156 12832
rect 7984 12792 7990 12804
rect 6503 12736 7328 12764
rect 6503 12733 6515 12736
rect 6457 12727 6515 12733
rect 5997 12699 6055 12705
rect 5997 12665 6009 12699
rect 6043 12696 6055 12699
rect 6196 12696 6224 12727
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 8128 12773 8156 12804
rect 9861 12801 9873 12835
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 10962 12792 10968 12844
rect 11020 12832 11026 12844
rect 14200 12832 14228 12928
rect 14642 12860 14648 12912
rect 14700 12900 14706 12912
rect 14918 12900 14924 12912
rect 14700 12872 14924 12900
rect 14700 12860 14706 12872
rect 14918 12860 14924 12872
rect 14976 12860 14982 12912
rect 16206 12860 16212 12912
rect 16264 12900 16270 12912
rect 16592 12900 16620 12940
rect 16666 12928 16672 12940
rect 16737 12968 16749 12971
rect 17678 12968 17684 12980
rect 16737 12940 17684 12968
rect 16737 12937 16749 12940
rect 16724 12931 16749 12937
rect 16724 12928 16730 12931
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 18877 12971 18935 12977
rect 18877 12937 18889 12971
rect 18923 12968 18935 12971
rect 19058 12968 19064 12980
rect 18923 12940 19064 12968
rect 18923 12937 18935 12940
rect 18877 12931 18935 12937
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 19245 12971 19303 12977
rect 19245 12937 19257 12971
rect 19291 12937 19303 12971
rect 21818 12968 21824 12980
rect 19245 12931 19303 12937
rect 19628 12940 21824 12968
rect 17494 12900 17500 12912
rect 16264 12872 16620 12900
rect 17312 12872 17500 12900
rect 16264 12860 16270 12872
rect 17312 12832 17340 12872
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 17770 12860 17776 12912
rect 17828 12900 17834 12912
rect 19260 12900 19288 12931
rect 17828 12872 19288 12900
rect 17828 12860 17834 12872
rect 11020 12804 13768 12832
rect 14200 12804 15036 12832
rect 11020 12792 11026 12804
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7708 12736 7849 12764
rect 7708 12724 7714 12736
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 8113 12767 8171 12773
rect 8113 12733 8125 12767
rect 8159 12733 8171 12767
rect 8113 12727 8171 12733
rect 9214 12724 9220 12776
rect 9272 12724 9278 12776
rect 9674 12724 9680 12776
rect 9732 12724 9738 12776
rect 12434 12724 12440 12776
rect 12492 12724 12498 12776
rect 13538 12724 13544 12776
rect 13596 12724 13602 12776
rect 13740 12773 13768 12804
rect 13725 12767 13783 12773
rect 13725 12733 13737 12767
rect 13771 12733 13783 12767
rect 13725 12727 13783 12733
rect 13906 12724 13912 12776
rect 13964 12724 13970 12776
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14240 12736 14933 12764
rect 14240 12724 14246 12736
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 15008 12764 15036 12804
rect 16132 12804 17340 12832
rect 15188 12767 15246 12773
rect 15188 12764 15200 12767
rect 15008 12736 15200 12764
rect 14921 12727 14979 12733
rect 15188 12733 15200 12736
rect 15234 12733 15246 12767
rect 15188 12727 15246 12733
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 15746 12764 15752 12776
rect 15528 12736 15752 12764
rect 15528 12724 15534 12736
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 7098 12696 7104 12708
rect 6043 12668 7104 12696
rect 6043 12665 6055 12668
rect 5997 12659 6055 12665
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 7190 12656 7196 12708
rect 7248 12656 7254 12708
rect 9585 12699 9643 12705
rect 9585 12665 9597 12699
rect 9631 12696 9643 12699
rect 9858 12696 9864 12708
rect 9631 12668 9864 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 9858 12656 9864 12668
rect 9916 12696 9922 12708
rect 10106 12699 10164 12705
rect 10106 12696 10118 12699
rect 9916 12668 10118 12696
rect 9916 12656 9922 12668
rect 10106 12665 10118 12668
rect 10152 12665 10164 12699
rect 11793 12699 11851 12705
rect 11793 12696 11805 12699
rect 10106 12659 10164 12665
rect 11256 12668 11805 12696
rect 4304 12600 4660 12628
rect 4709 12631 4767 12637
rect 4304 12588 4310 12600
rect 4709 12597 4721 12631
rect 4755 12628 4767 12631
rect 4982 12628 4988 12640
rect 4755 12600 4988 12628
rect 4755 12597 4767 12600
rect 4709 12591 4767 12597
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 6273 12631 6331 12637
rect 6273 12597 6285 12631
rect 6319 12628 6331 12631
rect 7466 12628 7472 12640
rect 6319 12600 7472 12628
rect 6319 12597 6331 12600
rect 6273 12591 6331 12597
rect 7466 12588 7472 12600
rect 7524 12628 7530 12640
rect 7745 12631 7803 12637
rect 7745 12628 7757 12631
rect 7524 12600 7757 12628
rect 7524 12588 7530 12600
rect 7745 12597 7757 12600
rect 7791 12597 7803 12631
rect 7745 12591 7803 12597
rect 8018 12588 8024 12640
rect 8076 12588 8082 12640
rect 11256 12637 11284 12668
rect 11793 12665 11805 12668
rect 11839 12665 11851 12699
rect 11793 12659 11851 12665
rect 12989 12699 13047 12705
rect 12989 12665 13001 12699
rect 13035 12696 13047 12699
rect 13035 12668 13308 12696
rect 13035 12665 13047 12668
rect 12989 12659 13047 12665
rect 11241 12631 11299 12637
rect 11241 12597 11253 12631
rect 11287 12597 11299 12631
rect 11241 12591 11299 12597
rect 11974 12588 11980 12640
rect 12032 12637 12038 12640
rect 12032 12631 12061 12637
rect 12049 12597 12061 12631
rect 12032 12591 12061 12597
rect 12032 12588 12038 12591
rect 12158 12588 12164 12640
rect 12216 12588 12222 12640
rect 12250 12588 12256 12640
rect 12308 12628 12314 12640
rect 12345 12631 12403 12637
rect 12345 12628 12357 12631
rect 12308 12600 12357 12628
rect 12308 12588 12314 12600
rect 12345 12597 12357 12600
rect 12391 12597 12403 12631
rect 12345 12591 12403 12597
rect 13078 12588 13084 12640
rect 13136 12628 13142 12640
rect 13189 12631 13247 12637
rect 13189 12628 13201 12631
rect 13136 12600 13201 12628
rect 13136 12588 13142 12600
rect 13189 12597 13201 12600
rect 13235 12597 13247 12631
rect 13280 12628 13308 12668
rect 14734 12656 14740 12708
rect 14792 12696 14798 12708
rect 16132 12696 16160 12804
rect 16700 12705 16728 12804
rect 17402 12792 17408 12844
rect 17460 12832 17466 12844
rect 17460 12804 18036 12832
rect 17460 12792 17466 12804
rect 17034 12724 17040 12776
rect 17092 12764 17098 12776
rect 17635 12767 17693 12773
rect 17635 12764 17647 12767
rect 17092 12736 17647 12764
rect 17092 12724 17098 12736
rect 17624 12733 17647 12736
rect 17681 12733 17693 12767
rect 17624 12727 17693 12733
rect 14792 12668 16160 12696
rect 16485 12699 16543 12705
rect 14792 12656 14798 12668
rect 16485 12665 16497 12699
rect 16531 12665 16543 12699
rect 16485 12659 16543 12665
rect 16685 12699 16743 12705
rect 16685 12665 16697 12699
rect 16731 12665 16743 12699
rect 16685 12659 16743 12665
rect 13446 12628 13452 12640
rect 13280 12600 13452 12628
rect 13189 12591 13247 12597
rect 13446 12588 13452 12600
rect 13504 12588 13510 12640
rect 16301 12631 16359 12637
rect 16301 12597 16313 12631
rect 16347 12628 16359 12631
rect 16500 12628 16528 12659
rect 16347 12600 16528 12628
rect 16347 12597 16359 12600
rect 16301 12591 16359 12597
rect 16850 12588 16856 12640
rect 16908 12588 16914 12640
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 17497 12631 17555 12637
rect 17497 12628 17509 12631
rect 17460 12600 17509 12628
rect 17460 12588 17466 12600
rect 17497 12597 17509 12600
rect 17543 12597 17555 12631
rect 17624 12628 17652 12727
rect 17770 12724 17776 12776
rect 17828 12724 17834 12776
rect 17862 12724 17868 12776
rect 17920 12724 17926 12776
rect 18008 12773 18036 12804
rect 18598 12792 18604 12844
rect 18656 12832 18662 12844
rect 19150 12832 19156 12844
rect 18656 12804 19156 12832
rect 18656 12792 18662 12804
rect 19150 12792 19156 12804
rect 19208 12832 19214 12844
rect 19628 12832 19656 12940
rect 21818 12928 21824 12940
rect 21876 12928 21882 12980
rect 22204 12940 23244 12968
rect 19705 12903 19763 12909
rect 19705 12869 19717 12903
rect 19751 12869 19763 12903
rect 19705 12863 19763 12869
rect 19208 12804 19656 12832
rect 19720 12832 19748 12863
rect 19720 12804 20576 12832
rect 19208 12792 19214 12804
rect 17993 12767 18051 12773
rect 17993 12733 18005 12767
rect 18039 12733 18051 12767
rect 17993 12727 18051 12733
rect 18138 12724 18144 12776
rect 18196 12724 18202 12776
rect 19242 12724 19248 12776
rect 19300 12724 19306 12776
rect 19426 12724 19432 12776
rect 19484 12724 19490 12776
rect 19521 12767 19579 12773
rect 19521 12733 19533 12767
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 20070 12764 20076 12776
rect 19843 12736 20076 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 17788 12668 18736 12696
rect 17788 12628 17816 12668
rect 17624 12600 17816 12628
rect 18708 12628 18736 12668
rect 18782 12656 18788 12708
rect 18840 12656 18846 12708
rect 19536 12696 19564 12727
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 20162 12724 20168 12776
rect 20220 12724 20226 12776
rect 20548 12773 20576 12804
rect 20622 12792 20628 12844
rect 20680 12832 20686 12844
rect 21453 12835 21511 12841
rect 21453 12832 21465 12835
rect 20680 12804 21465 12832
rect 20680 12792 20686 12804
rect 21453 12801 21465 12804
rect 21499 12801 21511 12835
rect 21453 12795 21511 12801
rect 20441 12767 20499 12773
rect 20441 12733 20453 12767
rect 20487 12733 20499 12767
rect 20441 12727 20499 12733
rect 20533 12767 20591 12773
rect 20533 12733 20545 12767
rect 20579 12733 20591 12767
rect 20533 12727 20591 12733
rect 20254 12696 20260 12708
rect 19536 12668 20260 12696
rect 20254 12656 20260 12668
rect 20312 12656 20318 12708
rect 20456 12696 20484 12727
rect 20898 12724 20904 12776
rect 20956 12724 20962 12776
rect 21154 12767 21212 12773
rect 21154 12733 21166 12767
rect 21200 12764 21212 12767
rect 22204 12764 22232 12940
rect 23216 12900 23244 12940
rect 23382 12928 23388 12980
rect 23440 12968 23446 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 23440 12940 24777 12968
rect 23440 12928 23446 12940
rect 24765 12937 24777 12940
rect 24811 12968 24823 12971
rect 24946 12968 24952 12980
rect 24811 12940 24952 12968
rect 24811 12937 24823 12940
rect 24765 12931 24823 12937
rect 24946 12928 24952 12940
rect 25004 12928 25010 12980
rect 25038 12928 25044 12980
rect 25096 12928 25102 12980
rect 25148 12940 29224 12968
rect 25148 12900 25176 12940
rect 23216 12872 25176 12900
rect 29196 12844 29224 12940
rect 30742 12928 30748 12980
rect 30800 12928 30806 12980
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12832 23259 12835
rect 25682 12832 25688 12844
rect 23247 12804 25688 12832
rect 23247 12801 23259 12804
rect 23201 12795 23259 12801
rect 25682 12792 25688 12804
rect 25740 12792 25746 12844
rect 29178 12792 29184 12844
rect 29236 12792 29242 12844
rect 21200 12736 22232 12764
rect 21200 12733 21212 12736
rect 21154 12727 21212 12733
rect 22554 12724 22560 12776
rect 22612 12764 22618 12776
rect 22945 12767 23003 12773
rect 22945 12764 22957 12767
rect 22612 12736 22957 12764
rect 22612 12724 22618 12736
rect 22945 12733 22957 12736
rect 22991 12764 23003 12767
rect 23382 12764 23388 12776
rect 22991 12736 23388 12764
rect 22991 12733 23003 12736
rect 22945 12727 23003 12733
rect 23382 12724 23388 12736
rect 23440 12724 23446 12776
rect 23842 12724 23848 12776
rect 23900 12764 23906 12776
rect 24029 12767 24087 12773
rect 24029 12764 24041 12767
rect 23900 12736 24041 12764
rect 23900 12724 23906 12736
rect 24029 12733 24041 12736
rect 24075 12733 24087 12767
rect 24029 12727 24087 12733
rect 24394 12724 24400 12776
rect 24452 12724 24458 12776
rect 24857 12767 24915 12773
rect 24857 12733 24869 12767
rect 24903 12764 24915 12767
rect 24949 12767 25007 12773
rect 24949 12764 24961 12767
rect 24903 12736 24961 12764
rect 24903 12733 24915 12736
rect 24857 12727 24915 12733
rect 24949 12733 24961 12736
rect 24995 12733 25007 12767
rect 24949 12727 25007 12733
rect 22738 12696 22744 12708
rect 20456 12668 22744 12696
rect 22738 12656 22744 12668
rect 22796 12656 22802 12708
rect 24121 12699 24179 12705
rect 24121 12665 24133 12699
rect 24167 12696 24179 12699
rect 24489 12699 24547 12705
rect 24489 12696 24501 12699
rect 24167 12668 24501 12696
rect 24167 12665 24179 12668
rect 24121 12659 24179 12665
rect 24489 12665 24501 12668
rect 24535 12696 24547 12699
rect 24872 12696 24900 12727
rect 25038 12724 25044 12776
rect 25096 12724 25102 12776
rect 25700 12764 25728 12792
rect 26697 12767 26755 12773
rect 26697 12764 26709 12767
rect 25700 12736 26709 12764
rect 26697 12733 26709 12736
rect 26743 12733 26755 12767
rect 26697 12727 26755 12733
rect 28994 12724 29000 12776
rect 29052 12724 29058 12776
rect 29086 12724 29092 12776
rect 29144 12764 29150 12776
rect 29365 12767 29423 12773
rect 29365 12764 29377 12767
rect 29144 12736 29377 12764
rect 29144 12724 29150 12736
rect 29365 12733 29377 12736
rect 29411 12733 29423 12767
rect 29365 12727 29423 12733
rect 29454 12724 29460 12776
rect 29512 12764 29518 12776
rect 29621 12767 29679 12773
rect 29621 12764 29633 12767
rect 29512 12736 29633 12764
rect 29512 12724 29518 12736
rect 29621 12733 29633 12736
rect 29667 12733 29679 12767
rect 29621 12727 29679 12733
rect 24535 12668 24900 12696
rect 25056 12696 25084 12724
rect 26418 12696 26424 12708
rect 26476 12705 26482 12708
rect 25056 12668 26424 12696
rect 24535 12665 24547 12668
rect 24489 12659 24547 12665
rect 26418 12656 26424 12668
rect 26476 12659 26488 12705
rect 26789 12699 26847 12705
rect 26789 12665 26801 12699
rect 26835 12665 26847 12699
rect 26789 12659 26847 12665
rect 26476 12656 26482 12659
rect 18966 12628 18972 12640
rect 18708 12600 18972 12628
rect 17497 12591 17555 12597
rect 18966 12588 18972 12600
rect 19024 12588 19030 12640
rect 19242 12588 19248 12640
rect 19300 12628 19306 12640
rect 19981 12631 20039 12637
rect 19981 12628 19993 12631
rect 19300 12600 19993 12628
rect 19300 12588 19306 12600
rect 19981 12597 19993 12600
rect 20027 12628 20039 12631
rect 20622 12628 20628 12640
rect 20027 12600 20628 12628
rect 20027 12597 20039 12600
rect 19981 12591 20039 12597
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 21821 12631 21879 12637
rect 21821 12597 21833 12631
rect 21867 12628 21879 12631
rect 22830 12628 22836 12640
rect 21867 12600 22836 12628
rect 21867 12597 21879 12600
rect 21821 12591 21879 12597
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 23014 12588 23020 12640
rect 23072 12628 23078 12640
rect 23382 12628 23388 12640
rect 23072 12600 23388 12628
rect 23072 12588 23078 12600
rect 23382 12588 23388 12600
rect 23440 12588 23446 12640
rect 25314 12588 25320 12640
rect 25372 12588 25378 12640
rect 25406 12588 25412 12640
rect 25464 12628 25470 12640
rect 26804 12628 26832 12659
rect 26970 12656 26976 12708
rect 27028 12696 27034 12708
rect 27525 12699 27583 12705
rect 27525 12696 27537 12699
rect 27028 12668 27537 12696
rect 27028 12656 27034 12668
rect 27525 12665 27537 12668
rect 27571 12665 27583 12699
rect 29012 12696 29040 12724
rect 29012 12668 29592 12696
rect 27525 12659 27583 12665
rect 25464 12600 26832 12628
rect 29089 12631 29147 12637
rect 25464 12588 25470 12600
rect 29089 12597 29101 12631
rect 29135 12628 29147 12631
rect 29270 12628 29276 12640
rect 29135 12600 29276 12628
rect 29135 12597 29147 12600
rect 29089 12591 29147 12597
rect 29270 12588 29276 12600
rect 29328 12588 29334 12640
rect 29564 12628 29592 12668
rect 29914 12628 29920 12640
rect 29564 12600 29920 12628
rect 29914 12588 29920 12600
rect 29972 12588 29978 12640
rect 552 12538 31531 12560
rect 552 12486 8102 12538
rect 8154 12486 8166 12538
rect 8218 12486 8230 12538
rect 8282 12486 8294 12538
rect 8346 12486 8358 12538
rect 8410 12486 15807 12538
rect 15859 12486 15871 12538
rect 15923 12486 15935 12538
rect 15987 12486 15999 12538
rect 16051 12486 16063 12538
rect 16115 12486 23512 12538
rect 23564 12486 23576 12538
rect 23628 12486 23640 12538
rect 23692 12486 23704 12538
rect 23756 12486 23768 12538
rect 23820 12486 31217 12538
rect 31269 12486 31281 12538
rect 31333 12486 31345 12538
rect 31397 12486 31409 12538
rect 31461 12486 31473 12538
rect 31525 12486 31531 12538
rect 552 12464 31531 12486
rect 1394 12384 1400 12436
rect 1452 12424 1458 12436
rect 1765 12427 1823 12433
rect 1765 12424 1777 12427
rect 1452 12396 1777 12424
rect 1452 12384 1458 12396
rect 1765 12393 1777 12396
rect 1811 12393 1823 12427
rect 1765 12387 1823 12393
rect 3973 12427 4031 12433
rect 3973 12393 3985 12427
rect 4019 12424 4031 12427
rect 4246 12424 4252 12436
rect 4019 12396 4252 12424
rect 4019 12393 4031 12396
rect 3973 12387 4031 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 5629 12427 5687 12433
rect 5629 12393 5641 12427
rect 5675 12393 5687 12427
rect 5629 12387 5687 12393
rect 6472 12396 6684 12424
rect 1578 12316 1584 12368
rect 1636 12356 1642 12368
rect 5644 12356 5672 12387
rect 6472 12365 6500 12396
rect 6457 12359 6515 12365
rect 1636 12328 1992 12356
rect 5644 12328 6316 12356
rect 1636 12316 1642 12328
rect 1596 12287 1624 12316
rect 1964 12297 1992 12328
rect 1857 12291 1915 12297
rect 1581 12281 1639 12287
rect 1581 12247 1593 12281
rect 1627 12247 1639 12281
rect 1857 12257 1869 12291
rect 1903 12257 1915 12291
rect 1857 12251 1915 12257
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12257 2007 12291
rect 1949 12251 2007 12257
rect 1581 12241 1639 12247
rect 1872 12220 1900 12251
rect 3694 12248 3700 12300
rect 3752 12288 3758 12300
rect 4522 12297 4528 12300
rect 3881 12291 3939 12297
rect 3881 12288 3893 12291
rect 3752 12260 3893 12288
rect 3752 12248 3758 12260
rect 3881 12257 3893 12260
rect 3927 12257 3939 12291
rect 4516 12288 4528 12297
rect 4483 12260 4528 12288
rect 3881 12251 3939 12257
rect 4516 12251 4528 12260
rect 4522 12248 4528 12251
rect 4580 12248 4586 12300
rect 6288 12297 6316 12328
rect 6457 12325 6469 12359
rect 6503 12325 6515 12359
rect 6457 12319 6515 12325
rect 6546 12316 6552 12368
rect 6604 12316 6610 12368
rect 6656 12356 6684 12396
rect 6822 12384 6828 12436
rect 6880 12384 6886 12436
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 8018 12424 8024 12436
rect 7156 12396 8024 12424
rect 7156 12384 7162 12396
rect 8018 12384 8024 12396
rect 8076 12384 8082 12436
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 9674 12424 9680 12436
rect 9447 12396 9680 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 9674 12384 9680 12396
rect 9732 12424 9738 12436
rect 9953 12427 10011 12433
rect 9953 12424 9965 12427
rect 9732 12396 9965 12424
rect 9732 12384 9738 12396
rect 9953 12393 9965 12396
rect 9999 12424 10011 12427
rect 9999 12396 10180 12424
rect 9999 12393 10011 12396
rect 9953 12387 10011 12393
rect 6914 12356 6920 12368
rect 6656 12328 6920 12356
rect 6914 12316 6920 12328
rect 6972 12316 6978 12368
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12257 6239 12291
rect 6181 12251 6239 12257
rect 6274 12291 6332 12297
rect 6274 12257 6286 12291
rect 6320 12257 6332 12291
rect 6274 12251 6332 12257
rect 6687 12291 6745 12297
rect 6687 12257 6699 12291
rect 6733 12288 6745 12291
rect 6822 12288 6828 12300
rect 6733 12260 6828 12288
rect 6733 12257 6745 12260
rect 6687 12251 6745 12257
rect 2041 12223 2099 12229
rect 2041 12220 2053 12223
rect 1872 12192 2053 12220
rect 1302 12112 1308 12164
rect 1360 12152 1366 12164
rect 1872 12152 1900 12192
rect 2041 12189 2053 12192
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12189 4307 12223
rect 6196 12220 6224 12251
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 7116 12286 7144 12384
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 7622 12359 7680 12365
rect 7622 12356 7634 12359
rect 7524 12328 7634 12356
rect 7524 12316 7530 12328
rect 7622 12325 7634 12328
rect 7668 12325 7680 12359
rect 7622 12319 7680 12325
rect 7742 12316 7748 12368
rect 7800 12356 7806 12368
rect 10042 12356 10048 12368
rect 7800 12328 10048 12356
rect 7800 12316 7806 12328
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 7185 12289 7243 12295
rect 7185 12286 7197 12289
rect 7116 12258 7197 12286
rect 7185 12255 7197 12258
rect 7231 12255 7243 12289
rect 7185 12249 7243 12255
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 9309 12291 9367 12297
rect 9309 12288 9321 12291
rect 9180 12260 9321 12288
rect 9180 12248 9186 12260
rect 9309 12257 9321 12260
rect 9355 12257 9367 12291
rect 9309 12251 9367 12257
rect 9582 12248 9588 12300
rect 9640 12248 9646 12300
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12288 9735 12291
rect 9766 12288 9772 12300
rect 9723 12260 9772 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 9858 12248 9864 12300
rect 9916 12248 9922 12300
rect 10152 12297 10180 12396
rect 11514 12384 11520 12436
rect 11572 12384 11578 12436
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 12250 12424 12256 12436
rect 11940 12396 12256 12424
rect 11940 12384 11946 12396
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 12618 12384 12624 12436
rect 12676 12424 12682 12436
rect 15378 12424 15384 12436
rect 12676 12396 15384 12424
rect 12676 12384 12682 12396
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 15528 12396 17172 12424
rect 15528 12384 15534 12396
rect 11532 12356 11560 12384
rect 11977 12359 12035 12365
rect 11977 12356 11989 12359
rect 11532 12328 11989 12356
rect 11977 12325 11989 12328
rect 12023 12325 12035 12359
rect 11977 12319 12035 12325
rect 12066 12316 12072 12368
rect 12124 12356 12130 12368
rect 12124 12328 12434 12356
rect 12124 12316 12130 12328
rect 10137 12291 10195 12297
rect 10137 12257 10149 12291
rect 10183 12257 10195 12291
rect 10137 12251 10195 12257
rect 11882 12248 11888 12300
rect 11940 12248 11946 12300
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12257 12219 12291
rect 12406 12288 12434 12328
rect 12986 12316 12992 12368
rect 13044 12316 13050 12368
rect 13078 12316 13084 12368
rect 13136 12356 13142 12368
rect 13189 12359 13247 12365
rect 13189 12356 13201 12359
rect 13136 12328 13201 12356
rect 13136 12316 13142 12328
rect 13189 12325 13201 12328
rect 13235 12325 13247 12359
rect 13189 12319 13247 12325
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 14369 12359 14427 12365
rect 14369 12356 14381 12359
rect 13780 12328 14381 12356
rect 13780 12316 13786 12328
rect 14369 12325 14381 12328
rect 14415 12356 14427 12359
rect 17034 12356 17040 12368
rect 14415 12328 17040 12356
rect 14415 12325 14427 12328
rect 14369 12319 14427 12325
rect 17034 12316 17040 12328
rect 17092 12316 17098 12368
rect 17144 12356 17172 12396
rect 17678 12384 17684 12436
rect 17736 12424 17742 12436
rect 18049 12427 18107 12433
rect 17736 12396 17908 12424
rect 17736 12384 17742 12396
rect 17563 12359 17621 12365
rect 17563 12356 17575 12359
rect 17144 12328 17575 12356
rect 17563 12325 17575 12328
rect 17609 12325 17621 12359
rect 17563 12319 17621 12325
rect 17770 12316 17776 12368
rect 17828 12316 17834 12368
rect 13096 12288 13124 12316
rect 12406 12260 13124 12288
rect 12161 12251 12219 12257
rect 7006 12220 7012 12232
rect 6196 12192 7012 12220
rect 4249 12183 4307 12189
rect 1360 12124 1900 12152
rect 1360 12112 1366 12124
rect 1486 12044 1492 12096
rect 1544 12044 1550 12096
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4264 12084 4292 12183
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 7208 12192 7389 12220
rect 7208 12164 7236 12192
rect 7377 12189 7389 12192
rect 7423 12189 7435 12223
rect 9784 12220 9812 12248
rect 10226 12220 10232 12232
rect 9784 12192 10232 12220
rect 7377 12183 7435 12189
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10962 12180 10968 12232
rect 11020 12180 11026 12232
rect 12176 12220 12204 12251
rect 11624 12192 12204 12220
rect 7190 12152 7196 12164
rect 5184 12124 7196 12152
rect 5184 12084 5212 12124
rect 7190 12112 7196 12124
rect 7248 12112 7254 12164
rect 8757 12155 8815 12161
rect 8757 12121 8769 12155
rect 8803 12152 8815 12155
rect 10980 12152 11008 12180
rect 11624 12164 11652 12192
rect 8803 12124 11008 12152
rect 8803 12121 8815 12124
rect 8757 12115 8815 12121
rect 11606 12112 11612 12164
rect 11664 12112 11670 12164
rect 13740 12152 13768 12316
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12288 14243 12291
rect 15194 12288 15200 12300
rect 14231 12260 15200 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 14936 12232 14964 12260
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15286 12248 15292 12300
rect 15344 12248 15350 12300
rect 15437 12291 15495 12297
rect 15437 12257 15449 12291
rect 15483 12288 15495 12291
rect 15483 12257 15516 12288
rect 15437 12251 15516 12257
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14001 12223 14059 12229
rect 14001 12220 14013 12223
rect 13872 12192 14013 12220
rect 13872 12180 13878 12192
rect 14001 12189 14013 12192
rect 14047 12189 14059 12223
rect 14001 12183 14059 12189
rect 13096 12124 13768 12152
rect 14016 12152 14044 12183
rect 14918 12180 14924 12232
rect 14976 12180 14982 12232
rect 15488 12220 15516 12251
rect 15562 12248 15568 12300
rect 15620 12248 15626 12300
rect 15654 12248 15660 12300
rect 15712 12248 15718 12300
rect 15746 12248 15752 12300
rect 15804 12297 15810 12300
rect 15804 12291 15853 12297
rect 15804 12257 15807 12291
rect 15841 12288 15853 12291
rect 16390 12288 16396 12300
rect 15841 12260 16396 12288
rect 15841 12257 15853 12260
rect 15804 12251 15853 12257
rect 15804 12248 15810 12251
rect 16390 12248 16396 12260
rect 16448 12248 16454 12300
rect 16574 12248 16580 12300
rect 16632 12288 16638 12300
rect 16758 12288 16764 12300
rect 16632 12260 16764 12288
rect 16632 12248 16638 12260
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 16850 12248 16856 12300
rect 16908 12294 16914 12300
rect 16945 12294 17003 12297
rect 16908 12291 17003 12294
rect 16908 12266 16957 12291
rect 16908 12248 16914 12266
rect 16945 12257 16957 12266
rect 16991 12257 17003 12291
rect 17129 12291 17187 12297
rect 17129 12288 17141 12291
rect 16945 12251 17003 12257
rect 17052 12260 17141 12288
rect 17052 12232 17080 12260
rect 17129 12257 17141 12260
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 17313 12291 17371 12297
rect 17313 12257 17325 12291
rect 17359 12288 17371 12291
rect 17359 12286 17451 12288
rect 17359 12260 17540 12286
rect 17359 12257 17371 12260
rect 17423 12258 17540 12260
rect 17313 12251 17371 12257
rect 16482 12220 16488 12232
rect 15488 12192 16488 12220
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 17034 12180 17040 12232
rect 17092 12180 17098 12232
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12189 17463 12223
rect 17405 12183 17463 12189
rect 15194 12152 15200 12164
rect 14016 12124 15200 12152
rect 4212 12056 5212 12084
rect 4212 12044 4218 12056
rect 7098 12044 7104 12096
rect 7156 12044 7162 12096
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 13096 12084 13124 12124
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 15930 12112 15936 12164
rect 15988 12112 15994 12164
rect 16022 12112 16028 12164
rect 16080 12152 16086 12164
rect 17411 12152 17439 12183
rect 16080 12124 17439 12152
rect 17512 12152 17540 12258
rect 17678 12248 17684 12300
rect 17736 12248 17742 12300
rect 17880 12297 17908 12396
rect 18049 12393 18061 12427
rect 18095 12424 18107 12427
rect 18138 12424 18144 12436
rect 18095 12396 18144 12424
rect 18095 12393 18107 12396
rect 18049 12387 18107 12393
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 18506 12384 18512 12436
rect 18564 12424 18570 12436
rect 18782 12424 18788 12436
rect 18564 12396 18788 12424
rect 18564 12384 18570 12396
rect 18782 12384 18788 12396
rect 18840 12424 18846 12436
rect 19334 12424 19340 12436
rect 18840 12396 19340 12424
rect 18840 12384 18846 12396
rect 19334 12384 19340 12396
rect 19392 12384 19398 12436
rect 19518 12384 19524 12436
rect 19576 12384 19582 12436
rect 21634 12384 21640 12436
rect 21692 12424 21698 12436
rect 23385 12427 23443 12433
rect 21692 12396 23060 12424
rect 21692 12384 21698 12396
rect 18230 12316 18236 12368
rect 18288 12356 18294 12368
rect 19058 12356 19064 12368
rect 18288 12328 19064 12356
rect 18288 12316 18294 12328
rect 19058 12316 19064 12328
rect 19116 12316 19122 12368
rect 19242 12316 19248 12368
rect 19300 12316 19306 12368
rect 19536 12356 19564 12384
rect 23032 12368 23060 12396
rect 23385 12393 23397 12427
rect 23431 12393 23443 12427
rect 23385 12387 23443 12393
rect 19536 12328 20116 12356
rect 17865 12291 17923 12297
rect 17865 12257 17877 12291
rect 17911 12288 17923 12291
rect 19260 12288 19288 12316
rect 17911 12260 19288 12288
rect 17911 12257 17923 12260
rect 17865 12251 17923 12257
rect 19334 12248 19340 12300
rect 19392 12248 19398 12300
rect 19429 12291 19487 12297
rect 19429 12257 19441 12291
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 19444 12220 19472 12251
rect 19610 12248 19616 12300
rect 19668 12248 19674 12300
rect 19981 12291 20039 12297
rect 19981 12257 19993 12291
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 18196 12192 19472 12220
rect 18196 12180 18202 12192
rect 17862 12152 17868 12164
rect 17512 12124 17868 12152
rect 16080 12112 16086 12124
rect 17862 12112 17868 12124
rect 17920 12112 17926 12164
rect 18598 12112 18604 12164
rect 18656 12152 18662 12164
rect 19886 12152 19892 12164
rect 18656 12124 19892 12152
rect 18656 12112 18662 12124
rect 19886 12112 19892 12124
rect 19944 12112 19950 12164
rect 19996 12152 20024 12251
rect 20088 12220 20116 12328
rect 20530 12316 20536 12368
rect 20588 12356 20594 12368
rect 21450 12356 21456 12368
rect 20588 12328 21456 12356
rect 20588 12316 20594 12328
rect 21450 12316 21456 12328
rect 21508 12316 21514 12368
rect 23014 12316 23020 12368
rect 23072 12316 23078 12368
rect 23106 12316 23112 12368
rect 23164 12316 23170 12368
rect 23400 12356 23428 12387
rect 23474 12384 23480 12436
rect 23532 12424 23538 12436
rect 23569 12427 23627 12433
rect 23569 12424 23581 12427
rect 23532 12396 23581 12424
rect 23532 12384 23538 12396
rect 23569 12393 23581 12396
rect 23615 12424 23627 12427
rect 24394 12424 24400 12436
rect 23615 12396 24400 12424
rect 23615 12393 23627 12396
rect 23569 12387 23627 12393
rect 24394 12384 24400 12396
rect 24452 12384 24458 12436
rect 24854 12424 24860 12436
rect 24780 12396 24860 12424
rect 24780 12356 24808 12396
rect 24854 12384 24860 12396
rect 24912 12384 24918 12436
rect 28626 12424 28632 12436
rect 25516 12396 28632 12424
rect 25516 12365 25544 12396
rect 28626 12384 28632 12396
rect 28684 12384 28690 12436
rect 23400 12328 24164 12356
rect 20234 12291 20292 12297
rect 20234 12257 20246 12291
rect 20280 12288 20292 12291
rect 22649 12291 22707 12297
rect 20280 12260 22508 12288
rect 20280 12257 20292 12260
rect 20234 12251 20292 12257
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 20088 12192 20545 12220
rect 20533 12189 20545 12192
rect 20579 12189 20591 12223
rect 20533 12183 20591 12189
rect 20898 12180 20904 12232
rect 20956 12180 20962 12232
rect 20070 12152 20076 12164
rect 19996 12124 20076 12152
rect 20070 12112 20076 12124
rect 20128 12152 20134 12164
rect 20916 12152 20944 12180
rect 20128 12124 20944 12152
rect 20128 12112 20134 12124
rect 8076 12056 13124 12084
rect 8076 12044 8082 12056
rect 13170 12044 13176 12096
rect 13228 12044 13234 12096
rect 13354 12044 13360 12096
rect 13412 12044 13418 12096
rect 16574 12044 16580 12096
rect 16632 12044 16638 12096
rect 16850 12044 16856 12096
rect 16908 12044 16914 12096
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17037 12087 17095 12093
rect 17037 12084 17049 12087
rect 17000 12056 17049 12084
rect 17000 12044 17006 12056
rect 17037 12053 17049 12056
rect 17083 12053 17095 12087
rect 17037 12047 17095 12053
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 22370 12084 22376 12096
rect 18288 12056 22376 12084
rect 18288 12044 18294 12056
rect 22370 12044 22376 12056
rect 22428 12044 22434 12096
rect 22480 12084 22508 12260
rect 22649 12257 22661 12291
rect 22695 12257 22707 12291
rect 22649 12251 22707 12257
rect 22664 12220 22692 12251
rect 22738 12248 22744 12300
rect 22796 12248 22802 12300
rect 22830 12248 22836 12300
rect 22888 12248 22894 12300
rect 23198 12248 23204 12300
rect 23256 12297 23262 12300
rect 23256 12288 23264 12297
rect 23477 12291 23535 12297
rect 23256 12260 23301 12288
rect 23256 12251 23264 12260
rect 23477 12257 23489 12291
rect 23523 12288 23535 12291
rect 23523 12260 23612 12288
rect 23523 12257 23535 12260
rect 23477 12251 23535 12257
rect 23256 12248 23262 12251
rect 22664 12192 22876 12220
rect 22848 12164 22876 12192
rect 23584 12164 23612 12260
rect 24026 12248 24032 12300
rect 24084 12248 24090 12300
rect 24136 12297 24164 12328
rect 24320 12328 24808 12356
rect 25501 12359 25559 12365
rect 24320 12297 24348 12328
rect 25501 12325 25513 12359
rect 25547 12325 25559 12359
rect 25501 12319 25559 12325
rect 26970 12316 26976 12368
rect 27028 12356 27034 12368
rect 29086 12356 29092 12368
rect 27028 12328 29092 12356
rect 27028 12316 27034 12328
rect 24121 12291 24179 12297
rect 24121 12257 24133 12291
rect 24167 12257 24179 12291
rect 24121 12251 24179 12257
rect 24305 12291 24363 12297
rect 24305 12257 24317 12291
rect 24351 12257 24363 12291
rect 24305 12251 24363 12257
rect 24670 12248 24676 12300
rect 24728 12248 24734 12300
rect 24926 12291 24984 12297
rect 24926 12257 24938 12291
rect 24972 12288 24984 12291
rect 28005 12291 28063 12297
rect 24972 12260 26924 12288
rect 24972 12257 24984 12260
rect 24926 12251 24984 12257
rect 22557 12155 22615 12161
rect 22557 12121 22569 12155
rect 22603 12152 22615 12155
rect 22646 12152 22652 12164
rect 22603 12124 22652 12152
rect 22603 12121 22615 12124
rect 22557 12115 22615 12121
rect 22646 12112 22652 12124
rect 22704 12112 22710 12164
rect 22830 12112 22836 12164
rect 22888 12112 22894 12164
rect 23566 12112 23572 12164
rect 23624 12112 23630 12164
rect 26896 12161 26924 12260
rect 28005 12257 28017 12291
rect 28051 12288 28063 12291
rect 28166 12288 28172 12300
rect 28051 12260 28172 12288
rect 28051 12257 28063 12260
rect 28005 12251 28063 12257
rect 28166 12248 28172 12260
rect 28224 12248 28230 12300
rect 28276 12297 28304 12328
rect 29086 12316 29092 12328
rect 29144 12356 29150 12368
rect 29144 12328 29868 12356
rect 29144 12316 29150 12328
rect 29840 12300 29868 12328
rect 28261 12291 28319 12297
rect 28261 12257 28273 12291
rect 28307 12257 28319 12291
rect 28261 12251 28319 12257
rect 29270 12248 29276 12300
rect 29328 12288 29334 12300
rect 29558 12291 29616 12297
rect 29558 12288 29570 12291
rect 29328 12260 29570 12288
rect 29328 12248 29334 12260
rect 29558 12257 29570 12260
rect 29604 12257 29616 12291
rect 29558 12251 29616 12257
rect 29822 12248 29828 12300
rect 29880 12248 29886 12300
rect 29914 12248 29920 12300
rect 29972 12248 29978 12300
rect 26881 12155 26939 12161
rect 26881 12121 26893 12155
rect 26927 12121 26939 12155
rect 26881 12115 26939 12121
rect 28445 12155 28503 12161
rect 28445 12121 28457 12155
rect 28491 12121 28503 12155
rect 28445 12115 28503 12121
rect 28460 12084 28488 12115
rect 22480 12056 28488 12084
rect 30009 12087 30067 12093
rect 30009 12053 30021 12087
rect 30055 12084 30067 12087
rect 30374 12084 30380 12096
rect 30055 12056 30380 12084
rect 30055 12053 30067 12056
rect 30009 12047 30067 12053
rect 30374 12044 30380 12056
rect 30432 12044 30438 12096
rect 552 11994 31372 12016
rect 552 11942 4250 11994
rect 4302 11942 4314 11994
rect 4366 11942 4378 11994
rect 4430 11942 4442 11994
rect 4494 11942 4506 11994
rect 4558 11942 11955 11994
rect 12007 11942 12019 11994
rect 12071 11942 12083 11994
rect 12135 11942 12147 11994
rect 12199 11942 12211 11994
rect 12263 11942 19660 11994
rect 19712 11942 19724 11994
rect 19776 11942 19788 11994
rect 19840 11942 19852 11994
rect 19904 11942 19916 11994
rect 19968 11942 27365 11994
rect 27417 11942 27429 11994
rect 27481 11942 27493 11994
rect 27545 11942 27557 11994
rect 27609 11942 27621 11994
rect 27673 11942 31372 11994
rect 552 11920 31372 11942
rect 1213 11883 1271 11889
rect 1213 11849 1225 11883
rect 1259 11880 1271 11883
rect 1394 11880 1400 11892
rect 1259 11852 1400 11880
rect 1259 11849 1271 11852
rect 1213 11843 1271 11849
rect 1394 11840 1400 11852
rect 1452 11840 1458 11892
rect 1486 11840 1492 11892
rect 1544 11840 1550 11892
rect 4154 11880 4160 11892
rect 3436 11852 4160 11880
rect 937 11747 995 11753
rect 937 11713 949 11747
rect 983 11744 995 11747
rect 983 11716 1164 11744
rect 983 11713 995 11716
rect 937 11707 995 11713
rect 1136 11685 1164 11716
rect 1029 11679 1087 11685
rect 1029 11645 1041 11679
rect 1075 11645 1087 11679
rect 1029 11639 1087 11645
rect 1121 11679 1179 11685
rect 1121 11645 1133 11679
rect 1167 11676 1179 11679
rect 1397 11679 1455 11685
rect 1397 11676 1409 11679
rect 1167 11648 1409 11676
rect 1167 11645 1179 11648
rect 1121 11639 1179 11645
rect 1397 11645 1409 11648
rect 1443 11676 1455 11679
rect 1504 11676 1532 11840
rect 1670 11704 1676 11756
rect 1728 11704 1734 11756
rect 3326 11744 3332 11756
rect 2746 11716 3332 11744
rect 1443 11648 1532 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1044 11552 1072 11639
rect 1578 11636 1584 11688
rect 1636 11636 1642 11688
rect 1688 11676 1716 11704
rect 2746 11676 2774 11716
rect 3326 11704 3332 11716
rect 3384 11744 3390 11756
rect 3436 11753 3464 11852
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 7742 11880 7748 11892
rect 5316 11852 7748 11880
rect 5316 11840 5322 11852
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 9401 11883 9459 11889
rect 9401 11849 9413 11883
rect 9447 11880 9459 11883
rect 9582 11880 9588 11892
rect 9447 11852 9588 11880
rect 9447 11849 9459 11852
rect 9401 11843 9459 11849
rect 4801 11815 4859 11821
rect 4801 11781 4813 11815
rect 4847 11781 4859 11815
rect 6086 11812 6092 11824
rect 4801 11775 4859 11781
rect 5920 11784 6092 11812
rect 3421 11747 3479 11753
rect 3421 11744 3433 11747
rect 3384 11716 3433 11744
rect 3384 11704 3390 11716
rect 3421 11713 3433 11716
rect 3467 11713 3479 11747
rect 4816 11744 4844 11775
rect 4816 11716 5764 11744
rect 3421 11707 3479 11713
rect 3694 11685 3700 11688
rect 3688 11676 3700 11685
rect 1688 11648 2774 11676
rect 3655 11648 3700 11676
rect 3688 11639 3700 11648
rect 3694 11636 3700 11639
rect 3752 11636 3758 11688
rect 5626 11636 5632 11688
rect 5684 11636 5690 11688
rect 5736 11685 5764 11716
rect 5920 11685 5948 11784
rect 6086 11772 6092 11784
rect 6144 11812 6150 11824
rect 6914 11812 6920 11824
rect 6144 11784 6920 11812
rect 6144 11772 6150 11784
rect 6914 11772 6920 11784
rect 6972 11812 6978 11824
rect 7650 11812 7656 11824
rect 6972 11784 7656 11812
rect 6972 11772 6978 11784
rect 7650 11772 7656 11784
rect 7708 11772 7714 11824
rect 9416 11744 9444 11843
rect 9582 11840 9588 11852
rect 9640 11880 9646 11892
rect 9677 11883 9735 11889
rect 9677 11880 9689 11883
rect 9640 11852 9689 11880
rect 9640 11840 9646 11852
rect 9677 11849 9689 11852
rect 9723 11849 9735 11883
rect 9677 11843 9735 11849
rect 9766 11840 9772 11892
rect 9824 11840 9830 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 9876 11852 14657 11880
rect 9784 11744 9812 11840
rect 7484 11716 9168 11744
rect 5722 11679 5780 11685
rect 5722 11645 5734 11679
rect 5768 11645 5780 11679
rect 5722 11639 5780 11645
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 5994 11636 6000 11688
rect 6052 11636 6058 11688
rect 7484 11685 7512 11716
rect 6135 11679 6193 11685
rect 6135 11645 6147 11679
rect 6181 11676 6193 11679
rect 7469 11679 7527 11685
rect 6181 11648 6592 11676
rect 6181 11645 6193 11648
rect 6135 11639 6193 11645
rect 1596 11608 1624 11636
rect 1918 11611 1976 11617
rect 1918 11608 1930 11611
rect 1596 11580 1930 11608
rect 1918 11577 1930 11580
rect 1964 11577 1976 11611
rect 1918 11571 1976 11577
rect 1026 11500 1032 11552
rect 1084 11500 1090 11552
rect 1489 11543 1547 11549
rect 1489 11509 1501 11543
rect 1535 11540 1547 11543
rect 1762 11540 1768 11552
rect 1535 11512 1768 11540
rect 1535 11509 1547 11512
rect 1489 11503 1547 11509
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 3053 11543 3111 11549
rect 3053 11509 3065 11543
rect 3099 11540 3111 11543
rect 4246 11540 4252 11552
rect 3099 11512 4252 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 6270 11500 6276 11552
rect 6328 11500 6334 11552
rect 6564 11540 6592 11648
rect 7469 11645 7481 11679
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 7562 11679 7620 11685
rect 7562 11645 7574 11679
rect 7608 11645 7620 11679
rect 7562 11639 7620 11645
rect 6638 11568 6644 11620
rect 6696 11608 6702 11620
rect 7576 11608 7604 11639
rect 7834 11636 7840 11688
rect 7892 11636 7898 11688
rect 8018 11685 8024 11688
rect 7975 11679 8024 11685
rect 7975 11645 7987 11679
rect 8021 11645 8024 11679
rect 7975 11639 8024 11645
rect 7990 11636 8024 11639
rect 8076 11636 8082 11688
rect 6696 11580 7604 11608
rect 6696 11568 6702 11580
rect 7742 11568 7748 11620
rect 7800 11568 7806 11620
rect 6822 11540 6828 11552
rect 6564 11512 6828 11540
rect 6822 11500 6828 11512
rect 6880 11540 6886 11552
rect 7990 11540 8018 11636
rect 9140 11608 9168 11716
rect 9232 11716 9444 11744
rect 9646 11716 9812 11744
rect 9232 11685 9260 11716
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11645 9275 11679
rect 9217 11639 9275 11645
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11676 9367 11679
rect 9490 11676 9496 11688
rect 9355 11648 9496 11676
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 9490 11636 9496 11648
rect 9548 11676 9554 11688
rect 9646 11676 9674 11716
rect 9548 11648 9674 11676
rect 9548 11636 9554 11648
rect 9766 11636 9772 11688
rect 9824 11636 9830 11688
rect 9876 11608 9904 11852
rect 14645 11849 14657 11852
rect 14691 11849 14703 11883
rect 14645 11843 14703 11849
rect 14826 11840 14832 11892
rect 14884 11880 14890 11892
rect 16577 11883 16635 11889
rect 16577 11880 16589 11883
rect 14884 11852 16589 11880
rect 14884 11840 14890 11852
rect 16577 11849 16589 11852
rect 16623 11849 16635 11883
rect 16577 11843 16635 11849
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 18049 11883 18107 11889
rect 18049 11880 18061 11883
rect 16816 11852 18061 11880
rect 16816 11840 16822 11852
rect 18049 11849 18061 11852
rect 18095 11849 18107 11883
rect 18049 11843 18107 11849
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 19610 11880 19616 11892
rect 19116 11852 19616 11880
rect 19116 11840 19122 11852
rect 19610 11840 19616 11852
rect 19668 11840 19674 11892
rect 19904 11852 20760 11880
rect 11793 11815 11851 11821
rect 11793 11781 11805 11815
rect 11839 11812 11851 11815
rect 11974 11812 11980 11824
rect 11839 11784 11980 11812
rect 11839 11781 11851 11784
rect 11793 11775 11851 11781
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 16482 11772 16488 11824
rect 16540 11812 16546 11824
rect 16942 11812 16948 11824
rect 16540 11784 16948 11812
rect 16540 11772 16546 11784
rect 16942 11772 16948 11784
rect 17000 11772 17006 11824
rect 17037 11815 17095 11821
rect 17037 11781 17049 11815
rect 17083 11812 17095 11815
rect 19904 11812 19932 11852
rect 17083 11784 19932 11812
rect 17083 11781 17095 11784
rect 17037 11775 17095 11781
rect 13280 11716 13768 11744
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 11790 11676 11796 11688
rect 10008 11648 11796 11676
rect 10008 11636 10014 11648
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 11882 11636 11888 11688
rect 11940 11636 11946 11688
rect 11974 11636 11980 11688
rect 12032 11636 12038 11688
rect 13280 11676 13308 11716
rect 13740 11685 13768 11716
rect 14090 11704 14096 11756
rect 14148 11744 14154 11756
rect 14148 11716 15056 11744
rect 14148 11704 14154 11716
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 12084 11648 13308 11676
rect 13372 11648 13553 11676
rect 10226 11617 10232 11620
rect 10220 11608 10232 11617
rect 9140 11580 9904 11608
rect 10187 11580 10232 11608
rect 10220 11571 10232 11580
rect 10226 11568 10232 11571
rect 10284 11568 10290 11620
rect 11422 11568 11428 11620
rect 11480 11608 11486 11620
rect 12084 11608 12112 11648
rect 12244 11611 12302 11617
rect 12244 11608 12256 11611
rect 11480 11580 12112 11608
rect 12156 11580 12256 11608
rect 11480 11568 11486 11580
rect 6880 11512 8018 11540
rect 6880 11500 6886 11512
rect 8110 11500 8116 11552
rect 8168 11500 8174 11552
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 9122 11540 9128 11552
rect 8536 11512 9128 11540
rect 8536 11500 8542 11512
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 11296 11512 11345 11540
rect 11296 11500 11302 11512
rect 11333 11509 11345 11512
rect 11379 11509 11391 11543
rect 11333 11503 11391 11509
rect 11514 11500 11520 11552
rect 11572 11540 11578 11552
rect 12156 11540 12184 11580
rect 12244 11577 12256 11580
rect 12290 11608 12302 11611
rect 12894 11608 12900 11620
rect 12290 11580 12900 11608
rect 12290 11577 12302 11580
rect 12244 11571 12302 11577
rect 12894 11568 12900 11580
rect 12952 11568 12958 11620
rect 13372 11549 13400 11648
rect 13541 11645 13553 11648
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 13740 11608 13768 11639
rect 13814 11636 13820 11688
rect 13872 11636 13878 11688
rect 13906 11636 13912 11688
rect 13964 11636 13970 11688
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 14642 11676 14648 11688
rect 14056 11648 14648 11676
rect 14056 11636 14062 11648
rect 14642 11636 14648 11648
rect 14700 11676 14706 11688
rect 15028 11685 15056 11716
rect 15166 11716 15608 11744
rect 15166 11685 15194 11716
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 14700 11648 14841 11676
rect 14700 11636 14706 11648
rect 14829 11645 14841 11648
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 15013 11679 15071 11685
rect 15013 11645 15025 11679
rect 15059 11645 15071 11679
rect 15013 11639 15071 11645
rect 15131 11679 15194 11685
rect 15131 11645 15143 11679
rect 15177 11648 15194 11679
rect 15289 11679 15347 11685
rect 15177 11645 15189 11648
rect 15131 11639 15189 11645
rect 15289 11645 15301 11679
rect 15335 11645 15347 11679
rect 15289 11639 15347 11645
rect 14274 11608 14280 11620
rect 13740 11580 14280 11608
rect 14274 11568 14280 11580
rect 14332 11568 14338 11620
rect 14734 11568 14740 11620
rect 14792 11608 14798 11620
rect 14921 11611 14979 11617
rect 14921 11608 14933 11611
rect 14792 11580 14933 11608
rect 14792 11568 14798 11580
rect 14921 11577 14933 11580
rect 14967 11577 14979 11611
rect 14921 11571 14979 11577
rect 11572 11512 12184 11540
rect 13357 11543 13415 11549
rect 11572 11500 11578 11512
rect 13357 11509 13369 11543
rect 13403 11509 13415 11543
rect 13357 11503 13415 11509
rect 14093 11543 14151 11549
rect 14093 11509 14105 11543
rect 14139 11540 14151 11543
rect 15010 11540 15016 11552
rect 14139 11512 15016 11540
rect 14139 11509 14151 11512
rect 14093 11503 14151 11509
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15304 11540 15332 11639
rect 15580 11620 15608 11716
rect 16574 11704 16580 11756
rect 16632 11704 16638 11756
rect 16761 11747 16819 11753
rect 16761 11713 16773 11747
rect 16807 11744 16819 11747
rect 17218 11744 17224 11756
rect 16807 11716 17224 11744
rect 16807 11713 16819 11716
rect 16761 11707 16819 11713
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11744 18199 11747
rect 18598 11744 18604 11756
rect 18187 11716 18604 11744
rect 18187 11713 18199 11716
rect 18141 11707 18199 11713
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 19150 11704 19156 11756
rect 19208 11744 19214 11756
rect 20073 11747 20131 11753
rect 19208 11716 19840 11744
rect 19208 11704 19214 11716
rect 15562 11568 15568 11620
rect 15620 11568 15626 11620
rect 16592 11617 16620 11704
rect 16853 11679 16911 11685
rect 16853 11645 16865 11679
rect 16899 11676 16911 11679
rect 16942 11676 16948 11688
rect 16899 11648 16948 11676
rect 16899 11645 16911 11648
rect 16853 11639 16911 11645
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11676 18107 11679
rect 18230 11676 18236 11688
rect 18095 11648 18236 11676
rect 18095 11645 18107 11648
rect 18049 11639 18107 11645
rect 18230 11636 18236 11648
rect 18288 11636 18294 11688
rect 18325 11679 18383 11685
rect 18325 11645 18337 11679
rect 18371 11645 18383 11679
rect 18325 11639 18383 11645
rect 16577 11611 16635 11617
rect 16577 11577 16589 11611
rect 16623 11577 16635 11611
rect 16577 11571 16635 11577
rect 17402 11568 17408 11620
rect 17460 11608 17466 11620
rect 17954 11608 17960 11620
rect 17460 11580 17960 11608
rect 17460 11568 17466 11580
rect 17954 11568 17960 11580
rect 18012 11568 18018 11620
rect 18340 11608 18368 11639
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 18472 11648 18705 11676
rect 18472 11636 18478 11648
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 18874 11636 18880 11688
rect 18932 11636 18938 11688
rect 19702 11685 19708 11688
rect 19061 11679 19119 11685
rect 19061 11645 19073 11679
rect 19107 11645 19119 11679
rect 19429 11679 19487 11685
rect 19429 11676 19441 11679
rect 19061 11639 19119 11645
rect 19168 11648 19441 11676
rect 19076 11608 19104 11639
rect 18340 11580 18460 11608
rect 18432 11552 18460 11580
rect 18524 11580 19104 11608
rect 17862 11540 17868 11552
rect 15304 11512 17868 11540
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 18414 11500 18420 11552
rect 18472 11500 18478 11552
rect 18524 11549 18552 11580
rect 19168 11552 19196 11648
rect 19429 11645 19441 11648
rect 19475 11645 19487 11679
rect 19429 11639 19487 11645
rect 19682 11679 19708 11685
rect 19682 11645 19694 11679
rect 19682 11639 19708 11645
rect 19444 11608 19472 11639
rect 19702 11636 19708 11639
rect 19760 11636 19766 11688
rect 19812 11678 19840 11716
rect 20073 11713 20085 11747
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 19812 11670 19932 11678
rect 20088 11670 20116 11707
rect 19812 11650 20116 11670
rect 19904 11642 20116 11650
rect 20346 11636 20352 11688
rect 20404 11636 20410 11688
rect 20732 11685 20760 11852
rect 20806 11840 20812 11892
rect 20864 11880 20870 11892
rect 26145 11883 26203 11889
rect 26145 11880 26157 11883
rect 20864 11852 26157 11880
rect 20864 11840 20870 11852
rect 26145 11849 26157 11852
rect 26191 11849 26203 11883
rect 26145 11843 26203 11849
rect 28353 11883 28411 11889
rect 28353 11849 28365 11883
rect 28399 11880 28411 11883
rect 28629 11883 28687 11889
rect 28629 11880 28641 11883
rect 28399 11852 28641 11880
rect 28399 11849 28411 11852
rect 28353 11843 28411 11849
rect 28629 11849 28641 11852
rect 28675 11880 28687 11883
rect 28994 11880 29000 11892
rect 28675 11852 29000 11880
rect 28675 11849 28687 11852
rect 28629 11843 28687 11849
rect 28994 11840 29000 11852
rect 29052 11840 29058 11892
rect 29178 11840 29184 11892
rect 29236 11880 29242 11892
rect 29549 11883 29607 11889
rect 29549 11880 29561 11883
rect 29236 11852 29561 11880
rect 29236 11840 29242 11852
rect 29549 11849 29561 11852
rect 29595 11849 29607 11883
rect 29549 11843 29607 11849
rect 22002 11812 22008 11824
rect 21353 11784 22008 11812
rect 20533 11679 20591 11685
rect 20533 11645 20545 11679
rect 20579 11645 20591 11679
rect 20533 11639 20591 11645
rect 20717 11679 20775 11685
rect 20717 11645 20729 11679
rect 20763 11645 20775 11679
rect 20717 11639 20775 11645
rect 19794 11608 19800 11620
rect 19444 11580 19800 11608
rect 19794 11568 19800 11580
rect 19852 11568 19858 11620
rect 18509 11543 18567 11549
rect 18509 11509 18521 11543
rect 18555 11509 18567 11543
rect 18509 11503 18567 11509
rect 19150 11500 19156 11552
rect 19208 11500 19214 11552
rect 19610 11500 19616 11552
rect 19668 11540 19674 11552
rect 20548 11540 20576 11639
rect 20898 11636 20904 11688
rect 20956 11676 20962 11688
rect 21353 11685 21381 11784
rect 22002 11772 22008 11784
rect 22060 11772 22066 11824
rect 22830 11772 22836 11824
rect 22888 11812 22894 11824
rect 23017 11815 23075 11821
rect 23017 11812 23029 11815
rect 22888 11784 23029 11812
rect 22888 11772 22894 11784
rect 23017 11781 23029 11784
rect 23063 11781 23075 11815
rect 23017 11775 23075 11781
rect 21634 11704 21640 11756
rect 21692 11704 21698 11756
rect 23032 11744 23060 11775
rect 23290 11772 23296 11824
rect 23348 11812 23354 11824
rect 23937 11815 23995 11821
rect 23937 11812 23949 11815
rect 23348 11784 23949 11812
rect 23348 11772 23354 11784
rect 23937 11781 23949 11784
rect 23983 11781 23995 11815
rect 23937 11775 23995 11781
rect 24026 11772 24032 11824
rect 24084 11812 24090 11824
rect 24673 11815 24731 11821
rect 24673 11812 24685 11815
rect 24084 11784 24685 11812
rect 24084 11772 24090 11784
rect 24673 11781 24685 11784
rect 24719 11781 24731 11815
rect 24673 11775 24731 11781
rect 23566 11744 23572 11756
rect 22572 11716 22968 11744
rect 23032 11716 23572 11744
rect 22572 11688 22600 11716
rect 21085 11679 21143 11685
rect 21085 11676 21097 11679
rect 20956 11648 21097 11676
rect 20956 11636 20962 11648
rect 21085 11645 21097 11648
rect 21131 11645 21143 11679
rect 21085 11639 21143 11645
rect 21338 11679 21396 11685
rect 21338 11645 21350 11679
rect 21384 11645 21396 11679
rect 21338 11639 21396 11645
rect 21100 11608 21128 11639
rect 21450 11636 21456 11688
rect 21508 11636 21514 11688
rect 22097 11679 22155 11685
rect 22097 11645 22109 11679
rect 22143 11645 22155 11679
rect 22097 11639 22155 11645
rect 22189 11679 22247 11685
rect 22189 11645 22201 11679
rect 22235 11676 22247 11679
rect 22465 11679 22523 11685
rect 22465 11676 22477 11679
rect 22235 11648 22477 11676
rect 22235 11645 22247 11648
rect 22189 11639 22247 11645
rect 22465 11645 22477 11648
rect 22511 11676 22523 11679
rect 22511 11645 22524 11676
rect 22465 11639 22524 11645
rect 21468 11608 21496 11636
rect 21100 11580 21496 11608
rect 19668 11512 20576 11540
rect 22112 11540 22140 11639
rect 22496 11608 22524 11639
rect 22554 11636 22560 11688
rect 22612 11636 22618 11688
rect 22940 11685 22968 11716
rect 23566 11704 23572 11716
rect 23624 11704 23630 11756
rect 23842 11744 23848 11756
rect 23676 11716 23848 11744
rect 22833 11679 22891 11685
rect 22833 11645 22845 11679
rect 22879 11645 22891 11679
rect 22833 11639 22891 11645
rect 22925 11679 22983 11685
rect 22925 11645 22937 11679
rect 22971 11645 22983 11679
rect 22925 11639 22983 11645
rect 23201 11679 23259 11685
rect 23201 11645 23213 11679
rect 23247 11645 23259 11679
rect 23201 11639 23259 11645
rect 23293 11679 23351 11685
rect 23293 11645 23305 11679
rect 23339 11676 23351 11679
rect 23474 11676 23480 11688
rect 23339 11648 23480 11676
rect 23339 11645 23351 11648
rect 23293 11639 23351 11645
rect 22849 11608 22877 11639
rect 23216 11608 23244 11639
rect 23474 11636 23480 11648
rect 23532 11636 23538 11688
rect 23676 11685 23704 11716
rect 23842 11704 23848 11716
rect 23900 11704 23906 11756
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11744 24639 11747
rect 24762 11744 24768 11756
rect 24627 11716 24768 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 24762 11704 24768 11716
rect 24820 11704 24826 11756
rect 28166 11704 28172 11756
rect 28224 11744 28230 11756
rect 28224 11716 28764 11744
rect 28224 11704 28230 11716
rect 23661 11679 23719 11685
rect 23661 11645 23673 11679
rect 23707 11645 23719 11679
rect 23661 11639 23719 11645
rect 22496 11580 23244 11608
rect 22278 11540 22284 11552
rect 22112 11512 22284 11540
rect 19668 11500 19674 11512
rect 22278 11500 22284 11512
rect 22336 11500 22342 11552
rect 22741 11543 22799 11549
rect 22741 11509 22753 11543
rect 22787 11540 22799 11543
rect 22830 11540 22836 11552
rect 22787 11512 22836 11540
rect 22787 11509 22799 11512
rect 22741 11503 22799 11509
rect 22830 11500 22836 11512
rect 22888 11540 22894 11552
rect 23676 11540 23704 11639
rect 23934 11636 23940 11688
rect 23992 11676 23998 11688
rect 24121 11679 24179 11685
rect 24121 11676 24133 11679
rect 23992 11648 24133 11676
rect 23992 11636 23998 11648
rect 24121 11645 24133 11648
rect 24167 11645 24179 11679
rect 24121 11639 24179 11645
rect 24305 11679 24363 11685
rect 24305 11645 24317 11679
rect 24351 11676 24363 11679
rect 26053 11679 26111 11685
rect 24351 11648 25728 11676
rect 24351 11645 24363 11648
rect 24305 11639 24363 11645
rect 22888 11512 23704 11540
rect 23961 11540 23989 11636
rect 24026 11568 24032 11620
rect 24084 11608 24090 11620
rect 24213 11611 24271 11617
rect 24213 11608 24225 11611
rect 24084 11580 24225 11608
rect 24084 11568 24090 11580
rect 24213 11577 24225 11580
rect 24259 11577 24271 11611
rect 24213 11571 24271 11577
rect 24443 11611 24501 11617
rect 24443 11577 24455 11611
rect 24489 11608 24501 11611
rect 24578 11608 24584 11620
rect 24489 11580 24584 11608
rect 24489 11577 24501 11580
rect 24443 11571 24501 11577
rect 24578 11568 24584 11580
rect 24636 11568 24642 11620
rect 24854 11540 24860 11552
rect 23961 11512 24860 11540
rect 22888 11500 22894 11512
rect 24854 11500 24860 11512
rect 24912 11500 24918 11552
rect 25700 11540 25728 11648
rect 26053 11645 26065 11679
rect 26099 11676 26111 11679
rect 26234 11676 26240 11688
rect 26099 11648 26240 11676
rect 26099 11645 26111 11648
rect 26053 11639 26111 11645
rect 26234 11636 26240 11648
rect 26292 11676 26298 11688
rect 26970 11676 26976 11688
rect 26292 11648 26976 11676
rect 26292 11636 26298 11648
rect 26970 11636 26976 11648
rect 27028 11676 27034 11688
rect 28736 11685 28764 11716
rect 29270 11704 29276 11756
rect 29328 11744 29334 11756
rect 29328 11716 29500 11744
rect 29328 11704 29334 11716
rect 29472 11685 29500 11716
rect 27525 11679 27583 11685
rect 27525 11676 27537 11679
rect 27028 11648 27537 11676
rect 27028 11636 27034 11648
rect 27525 11645 27537 11648
rect 27571 11645 27583 11679
rect 27525 11639 27583 11645
rect 28261 11679 28319 11685
rect 28261 11645 28273 11679
rect 28307 11645 28319 11679
rect 28261 11639 28319 11645
rect 28721 11679 28779 11685
rect 28721 11645 28733 11679
rect 28767 11676 28779 11679
rect 28997 11679 29055 11685
rect 28997 11676 29009 11679
rect 28767 11648 29009 11676
rect 28767 11645 28779 11648
rect 28721 11639 28779 11645
rect 28997 11645 29009 11648
rect 29043 11645 29055 11679
rect 28997 11639 29055 11645
rect 29457 11679 29515 11685
rect 29457 11645 29469 11679
rect 29503 11645 29515 11679
rect 29457 11639 29515 11645
rect 25808 11611 25866 11617
rect 25808 11577 25820 11611
rect 25854 11608 25866 11611
rect 25958 11608 25964 11620
rect 25854 11580 25964 11608
rect 25854 11577 25866 11580
rect 25808 11571 25866 11577
rect 25958 11568 25964 11580
rect 26016 11568 26022 11620
rect 27246 11568 27252 11620
rect 27304 11617 27310 11620
rect 27304 11608 27316 11617
rect 27982 11608 27988 11620
rect 27304 11580 27988 11608
rect 27304 11571 27316 11580
rect 27304 11568 27310 11571
rect 27982 11568 27988 11580
rect 28040 11608 28046 11620
rect 28276 11608 28304 11639
rect 29822 11636 29828 11688
rect 29880 11676 29886 11688
rect 30282 11676 30288 11688
rect 29880 11648 30288 11676
rect 29880 11636 29886 11648
rect 30282 11636 30288 11648
rect 30340 11676 30346 11688
rect 30929 11679 30987 11685
rect 30929 11676 30941 11679
rect 30340 11648 30941 11676
rect 30340 11636 30346 11648
rect 30929 11645 30941 11648
rect 30975 11645 30987 11679
rect 30929 11639 30987 11645
rect 28040 11580 28304 11608
rect 28040 11568 28046 11580
rect 30374 11568 30380 11620
rect 30432 11608 30438 11620
rect 30662 11611 30720 11617
rect 30662 11608 30674 11611
rect 30432 11580 30674 11608
rect 30432 11568 30438 11580
rect 30662 11577 30674 11580
rect 30708 11577 30720 11611
rect 30662 11571 30720 11577
rect 28442 11540 28448 11552
rect 25700 11512 28448 11540
rect 28442 11500 28448 11512
rect 28500 11500 28506 11552
rect 28994 11500 29000 11552
rect 29052 11540 29058 11552
rect 29089 11543 29147 11549
rect 29089 11540 29101 11543
rect 29052 11512 29101 11540
rect 29052 11500 29058 11512
rect 29089 11509 29101 11512
rect 29135 11540 29147 11543
rect 29365 11543 29423 11549
rect 29365 11540 29377 11543
rect 29135 11512 29377 11540
rect 29135 11509 29147 11512
rect 29089 11503 29147 11509
rect 29365 11509 29377 11512
rect 29411 11509 29423 11543
rect 29365 11503 29423 11509
rect 552 11450 31531 11472
rect 552 11398 8102 11450
rect 8154 11398 8166 11450
rect 8218 11398 8230 11450
rect 8282 11398 8294 11450
rect 8346 11398 8358 11450
rect 8410 11398 15807 11450
rect 15859 11398 15871 11450
rect 15923 11398 15935 11450
rect 15987 11398 15999 11450
rect 16051 11398 16063 11450
rect 16115 11398 23512 11450
rect 23564 11398 23576 11450
rect 23628 11398 23640 11450
rect 23692 11398 23704 11450
rect 23756 11398 23768 11450
rect 23820 11398 31217 11450
rect 31269 11398 31281 11450
rect 31333 11398 31345 11450
rect 31397 11398 31409 11450
rect 31461 11398 31473 11450
rect 31525 11398 31531 11450
rect 552 11376 31531 11398
rect 1670 11296 1676 11348
rect 1728 11296 1734 11348
rect 3326 11296 3332 11348
rect 3384 11296 3390 11348
rect 4246 11296 4252 11348
rect 4304 11296 4310 11348
rect 6086 11296 6092 11348
rect 6144 11296 6150 11348
rect 6454 11296 6460 11348
rect 6512 11296 6518 11348
rect 7006 11296 7012 11348
rect 7064 11336 7070 11348
rect 9033 11339 9091 11345
rect 9033 11336 9045 11339
rect 7064 11308 9045 11336
rect 7064 11296 7070 11308
rect 9033 11305 9045 11308
rect 9079 11305 9091 11339
rect 9033 11299 9091 11305
rect 11624 11308 12296 11336
rect 1688 11268 1716 11296
rect 1320 11240 1716 11268
rect 1320 11209 1348 11240
rect 1305 11203 1363 11209
rect 1305 11169 1317 11203
rect 1351 11169 1363 11203
rect 1305 11163 1363 11169
rect 1394 11160 1400 11212
rect 1452 11200 1458 11212
rect 3344 11209 3372 11296
rect 4264 11268 4292 11296
rect 5353 11271 5411 11277
rect 5353 11268 5365 11271
rect 4264 11240 5365 11268
rect 5353 11237 5365 11240
rect 5399 11237 5411 11271
rect 5353 11231 5411 11237
rect 5445 11271 5503 11277
rect 5445 11237 5457 11271
rect 5491 11268 5503 11271
rect 5491 11240 6040 11268
rect 5491 11237 5503 11240
rect 5445 11231 5503 11237
rect 3602 11209 3608 11212
rect 1561 11203 1619 11209
rect 1561 11200 1573 11203
rect 1452 11172 1573 11200
rect 1452 11160 1458 11172
rect 1561 11169 1573 11172
rect 1607 11169 1619 11203
rect 1561 11163 1619 11169
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11169 3387 11203
rect 3329 11163 3387 11169
rect 3596 11163 3608 11209
rect 3602 11160 3608 11163
rect 3660 11160 3666 11212
rect 5258 11160 5264 11212
rect 5316 11160 5322 11212
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11200 5687 11203
rect 5718 11200 5724 11212
rect 5675 11172 5724 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 5906 11203 5964 11209
rect 5906 11169 5918 11203
rect 5952 11169 5964 11203
rect 5906 11163 5964 11169
rect 5077 11067 5135 11073
rect 5077 11033 5089 11067
rect 5123 11064 5135 11067
rect 5828 11064 5856 11163
rect 5123 11036 5856 11064
rect 5123 11033 5135 11036
rect 5077 11027 5135 11033
rect 2682 10956 2688 11008
rect 2740 10956 2746 11008
rect 4709 10999 4767 11005
rect 4709 10965 4721 10999
rect 4755 10996 4767 10999
rect 5920 10996 5948 11163
rect 6012 11132 6040 11240
rect 6104 11209 6132 11296
rect 11624 11280 11652 11308
rect 6178 11228 6184 11280
rect 6236 11228 6242 11280
rect 7276 11271 7334 11277
rect 7276 11237 7288 11271
rect 7322 11268 7334 11271
rect 8294 11268 8300 11280
rect 7322 11240 8300 11268
rect 7322 11237 7334 11240
rect 7276 11231 7334 11237
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11237 8815 11271
rect 11330 11268 11336 11280
rect 8757 11231 8815 11237
rect 8864 11240 11336 11268
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 6319 11203 6377 11209
rect 6319 11169 6331 11203
rect 6365 11200 6377 11203
rect 6822 11200 6828 11212
rect 6365 11172 6828 11200
rect 6365 11169 6377 11172
rect 6319 11163 6377 11169
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 6932 11172 8064 11200
rect 6932 11132 6960 11172
rect 6012 11104 6960 11132
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11101 7067 11135
rect 8036 11132 8064 11172
rect 8110 11160 8116 11212
rect 8168 11200 8174 11212
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 8168 11172 8493 11200
rect 8168 11160 8174 11172
rect 8481 11169 8493 11172
rect 8527 11169 8539 11203
rect 8481 11163 8539 11169
rect 8665 11203 8723 11209
rect 8665 11169 8677 11203
rect 8711 11169 8723 11203
rect 8665 11163 8723 11169
rect 8570 11132 8576 11144
rect 8036 11104 8576 11132
rect 7009 11095 7067 11101
rect 4755 10968 5948 10996
rect 7024 10996 7052 11095
rect 8570 11092 8576 11104
rect 8628 11132 8634 11144
rect 8680 11132 8708 11163
rect 8628 11104 8708 11132
rect 8628 11092 8634 11104
rect 8389 11067 8447 11073
rect 8389 11033 8401 11067
rect 8435 11064 8447 11067
rect 8772 11064 8800 11231
rect 8864 11209 8892 11240
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 11606 11228 11612 11280
rect 11664 11228 11670 11280
rect 12268 11268 12296 11308
rect 14274 11296 14280 11348
rect 14332 11336 14338 11348
rect 16022 11336 16028 11348
rect 14332 11308 16028 11336
rect 14332 11296 14338 11308
rect 16022 11296 16028 11308
rect 16080 11336 16086 11348
rect 16209 11339 16267 11345
rect 16209 11336 16221 11339
rect 16080 11308 16221 11336
rect 16080 11296 16086 11308
rect 16209 11305 16221 11308
rect 16255 11305 16267 11339
rect 16666 11336 16672 11348
rect 16209 11299 16267 11305
rect 16546 11308 16672 11336
rect 14430 11271 14488 11277
rect 14430 11268 14442 11271
rect 12268 11240 12480 11268
rect 8849 11203 8907 11209
rect 8849 11169 8861 11203
rect 8895 11169 8907 11203
rect 8849 11163 8907 11169
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11200 9459 11203
rect 9677 11203 9735 11209
rect 9447 11172 9628 11200
rect 9447 11169 9459 11172
rect 9401 11163 9459 11169
rect 9600 11076 9628 11172
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 9953 11203 10011 11209
rect 9953 11169 9965 11203
rect 9999 11200 10011 11203
rect 10229 11203 10287 11209
rect 10229 11200 10241 11203
rect 9999 11172 10241 11200
rect 9999 11169 10011 11172
rect 9953 11163 10011 11169
rect 10229 11169 10241 11172
rect 10275 11169 10287 11203
rect 10229 11163 10287 11169
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11200 10563 11203
rect 10551 11172 10732 11200
rect 10551 11169 10563 11172
rect 10505 11163 10563 11169
rect 9692 11132 9720 11163
rect 9766 11132 9772 11144
rect 9692 11104 9772 11132
rect 9766 11092 9772 11104
rect 9824 11132 9830 11144
rect 10134 11132 10140 11144
rect 9824 11104 10140 11132
rect 9824 11092 9830 11104
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 8435 11036 8800 11064
rect 9309 11067 9367 11073
rect 8435 11033 8447 11036
rect 8389 11027 8447 11033
rect 9309 11033 9321 11067
rect 9355 11064 9367 11067
rect 9490 11064 9496 11076
rect 9355 11036 9496 11064
rect 9355 11033 9367 11036
rect 9309 11027 9367 11033
rect 9490 11024 9496 11036
rect 9548 11024 9554 11076
rect 9582 11024 9588 11076
rect 9640 11064 9646 11076
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 9640 11036 9873 11064
rect 9640 11024 9646 11036
rect 9861 11033 9873 11036
rect 9907 11033 9919 11067
rect 10244 11064 10272 11163
rect 10704 11141 10732 11172
rect 10778 11160 10784 11212
rect 10836 11160 10842 11212
rect 11241 11203 11299 11209
rect 11241 11169 11253 11203
rect 11287 11200 11299 11203
rect 11425 11203 11483 11209
rect 11425 11200 11437 11203
rect 11287 11172 11437 11200
rect 11287 11169 11299 11172
rect 11241 11163 11299 11169
rect 11425 11169 11437 11172
rect 11471 11169 11483 11203
rect 11425 11163 11483 11169
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11132 10747 11135
rect 11256 11132 11284 11163
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 12452 11209 12480 11240
rect 13004 11240 14442 11268
rect 11885 11203 11943 11209
rect 11624 11172 11836 11200
rect 10735 11104 11284 11132
rect 10735 11101 10747 11104
rect 10689 11095 10747 11101
rect 11149 11067 11207 11073
rect 11149 11064 11161 11067
rect 10244 11036 11161 11064
rect 9861 11027 9919 11033
rect 11149 11033 11161 11036
rect 11195 11064 11207 11067
rect 11624 11064 11652 11172
rect 11808 11141 11836 11172
rect 11885 11169 11897 11203
rect 11931 11200 11943 11203
rect 12153 11206 12211 11209
rect 12153 11203 12287 11206
rect 12153 11200 12165 11203
rect 11931 11172 12165 11200
rect 11931 11169 11943 11172
rect 11885 11163 11943 11169
rect 12153 11169 12165 11172
rect 12199 11200 12287 11203
rect 12437 11203 12495 11209
rect 12199 11178 12388 11200
rect 12199 11169 12211 11178
rect 12259 11172 12388 11178
rect 12153 11163 12211 11169
rect 12360 11141 12388 11172
rect 12437 11169 12449 11203
rect 12483 11169 12495 11203
rect 12437 11163 12495 11169
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11200 12587 11203
rect 12894 11200 12900 11212
rect 12575 11172 12900 11200
rect 12575 11169 12587 11172
rect 12529 11163 12587 11169
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11132 11851 11135
rect 12345 11135 12403 11141
rect 11839 11104 12204 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 11195 11036 11652 11064
rect 11195 11033 11207 11036
rect 11149 11027 11207 11033
rect 7190 10996 7196 11008
rect 7024 10968 7196 10996
rect 4755 10965 4767 10968
rect 4709 10959 4767 10965
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 9398 10956 9404 11008
rect 9456 10996 9462 11008
rect 10042 10996 10048 11008
rect 9456 10968 10048 10996
rect 9456 10956 9462 10968
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 10134 10956 10140 11008
rect 10192 10956 10198 11008
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 10413 10999 10471 11005
rect 10413 10996 10425 10999
rect 10284 10968 10425 10996
rect 10284 10956 10290 10968
rect 10413 10965 10425 10968
rect 10459 10965 10471 10999
rect 10413 10959 10471 10965
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 12066 10996 12072 11008
rect 11940 10968 12072 10996
rect 11940 10956 11946 10968
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 12176 10996 12204 11104
rect 12345 11101 12357 11135
rect 12391 11132 12403 11135
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 12391 11104 12633 11132
rect 12391 11101 12403 11104
rect 12345 11095 12403 11101
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 13004 10996 13032 11240
rect 14430 11237 14442 11240
rect 14476 11237 14488 11271
rect 16546 11268 16574 11308
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 17218 11296 17224 11348
rect 17276 11296 17282 11348
rect 17313 11339 17371 11345
rect 17313 11305 17325 11339
rect 17359 11305 17371 11339
rect 17313 11299 17371 11305
rect 16945 11271 17003 11277
rect 14430 11231 14488 11237
rect 16316 11240 16620 11268
rect 14182 11160 14188 11212
rect 14240 11160 14246 11212
rect 16316 11200 16344 11240
rect 16592 11209 16620 11240
rect 16945 11237 16957 11271
rect 16991 11268 17003 11271
rect 17236 11268 17264 11296
rect 16991 11240 17264 11268
rect 17328 11268 17356 11299
rect 17494 11296 17500 11348
rect 17552 11336 17558 11348
rect 17678 11336 17684 11348
rect 17552 11308 17684 11336
rect 17552 11296 17558 11308
rect 17678 11296 17684 11308
rect 17736 11296 17742 11348
rect 17770 11296 17776 11348
rect 17828 11296 17834 11348
rect 17862 11296 17868 11348
rect 17920 11336 17926 11348
rect 20070 11336 20076 11348
rect 17920 11308 20076 11336
rect 17920 11296 17926 11308
rect 20070 11296 20076 11308
rect 20128 11296 20134 11348
rect 23017 11339 23075 11345
rect 23017 11336 23029 11339
rect 20364 11308 23029 11336
rect 17788 11268 17816 11296
rect 18046 11268 18052 11280
rect 17328 11240 17632 11268
rect 17788 11240 18052 11268
rect 16991 11237 17003 11240
rect 16945 11231 17003 11237
rect 14292 11172 16344 11200
rect 16393 11203 16451 11209
rect 13538 11092 13544 11144
rect 13596 11132 13602 11144
rect 14292 11132 14320 11172
rect 16393 11169 16405 11203
rect 16439 11190 16451 11203
rect 16577 11203 16635 11209
rect 16439 11169 16508 11190
rect 16393 11163 16508 11169
rect 16577 11169 16589 11203
rect 16623 11169 16635 11203
rect 16577 11163 16635 11169
rect 16413 11162 16508 11163
rect 16413 11132 16441 11162
rect 13596 11104 14320 11132
rect 16399 11104 16441 11132
rect 13596 11092 13602 11104
rect 15565 11067 15623 11073
rect 15565 11033 15577 11067
rect 15611 11064 15623 11067
rect 15838 11064 15844 11076
rect 15611 11036 15844 11064
rect 15611 11033 15623 11036
rect 15565 11027 15623 11033
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 16399 11064 16427 11104
rect 15948 11036 16427 11064
rect 16480 11064 16508 11162
rect 16666 11160 16672 11212
rect 16724 11160 16730 11212
rect 16850 11209 16856 11212
rect 16807 11203 16856 11209
rect 16807 11169 16819 11203
rect 16853 11169 16856 11203
rect 16807 11163 16856 11169
rect 16850 11160 16856 11163
rect 16908 11160 16914 11212
rect 17034 11160 17040 11212
rect 17092 11160 17098 11212
rect 17175 11203 17233 11209
rect 17175 11169 17187 11203
rect 17221 11169 17233 11203
rect 17175 11163 17233 11169
rect 17190 11132 17218 11163
rect 17402 11160 17408 11212
rect 17460 11160 17466 11212
rect 17604 11209 17632 11240
rect 18046 11228 18052 11240
rect 18104 11228 18110 11280
rect 19150 11268 19156 11280
rect 18248 11240 19156 11268
rect 18248 11212 18276 11240
rect 19150 11228 19156 11240
rect 19208 11228 19214 11280
rect 17589 11203 17647 11209
rect 17589 11169 17601 11203
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 17862 11160 17868 11212
rect 17920 11160 17926 11212
rect 18141 11203 18199 11209
rect 18141 11169 18153 11203
rect 18187 11200 18199 11203
rect 18230 11200 18236 11212
rect 18187 11172 18236 11200
rect 18187 11169 18199 11172
rect 18141 11163 18199 11169
rect 18230 11160 18236 11172
rect 18288 11160 18294 11212
rect 18394 11203 18452 11209
rect 18394 11169 18406 11203
rect 18440 11200 18452 11203
rect 20364 11200 20392 11308
rect 23017 11305 23029 11308
rect 23063 11305 23075 11339
rect 23017 11299 23075 11305
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 24394 11336 24400 11348
rect 23256 11308 24400 11336
rect 23256 11296 23262 11308
rect 24394 11296 24400 11308
rect 24452 11296 24458 11348
rect 27246 11296 27252 11348
rect 27304 11296 27310 11348
rect 28166 11296 28172 11348
rect 28224 11336 28230 11348
rect 28353 11339 28411 11345
rect 28353 11336 28365 11339
rect 28224 11308 28365 11336
rect 28224 11296 28230 11308
rect 28353 11305 28365 11308
rect 28399 11305 28411 11339
rect 28353 11299 28411 11305
rect 28442 11296 28448 11348
rect 28500 11336 28506 11348
rect 29181 11339 29239 11345
rect 28500 11308 28672 11336
rect 28500 11296 28506 11308
rect 20564 11271 20622 11277
rect 20564 11237 20576 11271
rect 20610 11268 20622 11271
rect 21266 11268 21272 11280
rect 20610 11240 21272 11268
rect 20610 11237 20622 11240
rect 20564 11231 20622 11237
rect 21266 11228 21272 11240
rect 21324 11228 21330 11280
rect 22186 11228 22192 11280
rect 22244 11268 22250 11280
rect 26234 11268 26240 11280
rect 22244 11240 26240 11268
rect 22244 11228 22250 11240
rect 18440 11172 20392 11200
rect 20809 11203 20867 11209
rect 18440 11169 18452 11172
rect 18394 11163 18452 11169
rect 20809 11169 20821 11203
rect 20855 11200 20867 11203
rect 20990 11200 20996 11212
rect 20855 11172 20996 11200
rect 20855 11169 20867 11172
rect 20809 11163 20867 11169
rect 20990 11160 20996 11172
rect 21048 11160 21054 11212
rect 22002 11160 22008 11212
rect 22060 11200 22066 11212
rect 22382 11203 22440 11209
rect 22382 11200 22394 11203
rect 22060 11172 22394 11200
rect 22060 11160 22066 11172
rect 22382 11169 22394 11172
rect 22428 11200 22440 11203
rect 22554 11200 22560 11212
rect 22428 11172 22560 11200
rect 22428 11169 22440 11172
rect 22382 11163 22440 11169
rect 22554 11160 22560 11172
rect 22612 11160 22618 11212
rect 22664 11209 22692 11240
rect 22649 11203 22707 11209
rect 22649 11169 22661 11203
rect 22695 11169 22707 11203
rect 22649 11163 22707 11169
rect 22738 11160 22744 11212
rect 22796 11160 22802 11212
rect 24412 11209 24440 11240
rect 26234 11228 26240 11240
rect 26292 11228 26298 11280
rect 28074 11268 28080 11280
rect 26896 11240 27476 11268
rect 24141 11203 24199 11209
rect 24141 11169 24153 11203
rect 24187 11200 24199 11203
rect 24397 11203 24455 11209
rect 24187 11172 24348 11200
rect 24187 11169 24199 11172
rect 24141 11163 24199 11169
rect 17494 11132 17500 11144
rect 17190 11104 17500 11132
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 18690 11092 18696 11144
rect 18748 11092 18754 11144
rect 18966 11092 18972 11144
rect 19024 11132 19030 11144
rect 19150 11132 19156 11144
rect 19024 11104 19156 11132
rect 19024 11092 19030 11104
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 22563 11132 22591 11160
rect 22833 11135 22891 11141
rect 22833 11132 22845 11135
rect 22563 11104 22845 11132
rect 22833 11101 22845 11104
rect 22879 11101 22891 11135
rect 24320 11132 24348 11172
rect 24397 11169 24409 11203
rect 24443 11169 24455 11203
rect 24397 11163 24455 11169
rect 25498 11160 25504 11212
rect 25556 11160 25562 11212
rect 26896 11209 26924 11240
rect 27448 11209 27476 11240
rect 27908 11240 28080 11268
rect 27908 11209 27936 11240
rect 28074 11228 28080 11240
rect 28132 11268 28138 11280
rect 28644 11268 28672 11308
rect 29181 11305 29193 11339
rect 29227 11336 29239 11339
rect 29270 11336 29276 11348
rect 29227 11308 29276 11336
rect 29227 11305 29239 11308
rect 29181 11299 29239 11305
rect 29270 11296 29276 11308
rect 29328 11296 29334 11348
rect 29549 11339 29607 11345
rect 29549 11305 29561 11339
rect 29595 11305 29607 11339
rect 29549 11299 29607 11305
rect 29564 11268 29592 11299
rect 28132 11240 28580 11268
rect 28644 11240 29592 11268
rect 30300 11240 30972 11268
rect 28132 11228 28138 11240
rect 28552 11209 28580 11240
rect 30300 11212 30328 11240
rect 26881 11203 26939 11209
rect 26881 11200 26893 11203
rect 26436 11172 26893 11200
rect 26436 11144 26464 11172
rect 26881 11169 26893 11172
rect 26927 11169 26939 11203
rect 26881 11163 26939 11169
rect 27157 11203 27215 11209
rect 27157 11169 27169 11203
rect 27203 11169 27215 11203
rect 27157 11163 27215 11169
rect 27433 11203 27491 11209
rect 27433 11169 27445 11203
rect 27479 11169 27491 11203
rect 27433 11163 27491 11169
rect 27893 11203 27951 11209
rect 27893 11169 27905 11203
rect 27939 11169 27951 11203
rect 27893 11163 27951 11169
rect 28169 11203 28227 11209
rect 28169 11169 28181 11203
rect 28215 11200 28227 11203
rect 28261 11203 28319 11209
rect 28261 11200 28273 11203
rect 28215 11172 28273 11200
rect 28215 11169 28227 11172
rect 28169 11163 28227 11169
rect 28261 11169 28273 11172
rect 28307 11169 28319 11203
rect 28261 11163 28319 11169
rect 28537 11203 28595 11209
rect 28537 11169 28549 11203
rect 28583 11169 28595 11203
rect 28537 11163 28595 11169
rect 28813 11203 28871 11209
rect 28813 11169 28825 11203
rect 28859 11169 28871 11203
rect 29089 11203 29147 11209
rect 29089 11200 29101 11203
rect 28813 11163 28871 11169
rect 28920 11172 29101 11200
rect 26418 11132 26424 11144
rect 24320 11104 26424 11132
rect 22833 11095 22891 11101
rect 26418 11092 26424 11104
rect 26476 11092 26482 11144
rect 26973 11135 27031 11141
rect 26973 11101 26985 11135
rect 27019 11132 27031 11135
rect 27172 11132 27200 11163
rect 27246 11132 27252 11144
rect 27019 11104 27252 11132
rect 27019 11101 27031 11104
rect 26973 11095 27031 11101
rect 27246 11092 27252 11104
rect 27304 11092 27310 11144
rect 28184 11132 28212 11163
rect 27816 11104 28212 11132
rect 17034 11064 17040 11076
rect 16480 11036 17040 11064
rect 12176 10968 13032 10996
rect 14458 10956 14464 11008
rect 14516 10996 14522 11008
rect 15948 10996 15976 11036
rect 17034 11024 17040 11036
rect 17092 11024 17098 11076
rect 20806 11024 20812 11076
rect 20864 11024 20870 11076
rect 24670 11024 24676 11076
rect 24728 11024 24734 11076
rect 27816 11073 27844 11104
rect 27525 11067 27583 11073
rect 27525 11033 27537 11067
rect 27571 11064 27583 11067
rect 27801 11067 27859 11073
rect 27801 11064 27813 11067
rect 27571 11036 27813 11064
rect 27571 11033 27583 11036
rect 27525 11027 27583 11033
rect 27801 11033 27813 11036
rect 27847 11033 27859 11067
rect 27801 11027 27859 11033
rect 27982 11024 27988 11076
rect 28040 11064 28046 11076
rect 28077 11067 28135 11073
rect 28077 11064 28089 11067
rect 28040 11036 28089 11064
rect 28040 11024 28046 11036
rect 28077 11033 28089 11036
rect 28123 11064 28135 11067
rect 28828 11064 28856 11163
rect 28123 11036 28856 11064
rect 28123 11033 28135 11036
rect 28077 11027 28135 11033
rect 14516 10968 15976 10996
rect 14516 10956 14522 10968
rect 16022 10956 16028 11008
rect 16080 10996 16086 11008
rect 16298 10996 16304 11008
rect 16080 10968 16304 10996
rect 16080 10956 16086 10968
rect 16298 10956 16304 10968
rect 16356 10956 16362 11008
rect 18322 10956 18328 11008
rect 18380 10996 18386 11008
rect 18966 10996 18972 11008
rect 18380 10968 18972 10996
rect 18380 10956 18386 10968
rect 18966 10956 18972 10968
rect 19024 10956 19030 11008
rect 19429 10999 19487 11005
rect 19429 10965 19441 10999
rect 19475 10996 19487 10999
rect 20070 10996 20076 11008
rect 19475 10968 20076 10996
rect 19475 10965 19487 10968
rect 19429 10959 19487 10965
rect 20070 10956 20076 10968
rect 20128 10956 20134 11008
rect 20824 10996 20852 11024
rect 21269 10999 21327 11005
rect 21269 10996 21281 10999
rect 20824 10968 21281 10996
rect 21269 10965 21281 10968
rect 21315 10965 21327 10999
rect 21269 10959 21327 10965
rect 21450 10956 21456 11008
rect 21508 10996 21514 11008
rect 24688 10996 24716 11024
rect 21508 10968 24716 10996
rect 21508 10956 21514 10968
rect 25590 10956 25596 11008
rect 25648 10996 25654 11008
rect 26786 10996 26792 11008
rect 25648 10968 26792 10996
rect 25648 10956 25654 10968
rect 26786 10956 26792 10968
rect 26844 10956 26850 11008
rect 28442 10956 28448 11008
rect 28500 10996 28506 11008
rect 28920 11005 28948 11172
rect 29089 11169 29101 11172
rect 29135 11169 29147 11203
rect 29089 11163 29147 11169
rect 30282 11160 30288 11212
rect 30340 11160 30346 11212
rect 30650 11160 30656 11212
rect 30708 11209 30714 11212
rect 30944 11209 30972 11240
rect 30708 11163 30720 11209
rect 30929 11203 30987 11209
rect 30929 11169 30941 11203
rect 30975 11169 30987 11203
rect 30929 11163 30987 11169
rect 30708 11160 30714 11163
rect 28629 10999 28687 11005
rect 28629 10996 28641 10999
rect 28500 10968 28641 10996
rect 28500 10956 28506 10968
rect 28629 10965 28641 10968
rect 28675 10996 28687 10999
rect 28905 10999 28963 11005
rect 28905 10996 28917 10999
rect 28675 10968 28917 10996
rect 28675 10965 28687 10968
rect 28629 10959 28687 10965
rect 28905 10965 28917 10968
rect 28951 10965 28963 10999
rect 28905 10959 28963 10965
rect 552 10906 31372 10928
rect 552 10854 4250 10906
rect 4302 10854 4314 10906
rect 4366 10854 4378 10906
rect 4430 10854 4442 10906
rect 4494 10854 4506 10906
rect 4558 10854 11955 10906
rect 12007 10854 12019 10906
rect 12071 10854 12083 10906
rect 12135 10854 12147 10906
rect 12199 10854 12211 10906
rect 12263 10854 19660 10906
rect 19712 10854 19724 10906
rect 19776 10854 19788 10906
rect 19840 10854 19852 10906
rect 19904 10854 19916 10906
rect 19968 10854 27365 10906
rect 27417 10854 27429 10906
rect 27481 10854 27493 10906
rect 27545 10854 27557 10906
rect 27609 10854 27621 10906
rect 27673 10854 31372 10906
rect 552 10832 31372 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 1762 10792 1768 10804
rect 1627 10764 1768 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 5258 10752 5264 10804
rect 5316 10752 5322 10804
rect 5537 10795 5595 10801
rect 5537 10761 5549 10795
rect 5583 10792 5595 10795
rect 5626 10792 5632 10804
rect 5583 10764 5632 10792
rect 5583 10761 5595 10764
rect 5537 10755 5595 10761
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 5736 10764 8892 10792
rect 5276 10724 5304 10752
rect 1044 10696 2084 10724
rect 5276 10696 5396 10724
rect 1044 10668 1072 10696
rect 1026 10616 1032 10668
rect 1084 10616 1090 10668
rect 1394 10616 1400 10668
rect 1452 10656 1458 10668
rect 1452 10628 1808 10656
rect 1452 10616 1458 10628
rect 1780 10597 1808 10628
rect 2056 10597 2084 10696
rect 2700 10628 5304 10656
rect 2700 10600 2728 10628
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10557 1731 10591
rect 1673 10551 1731 10557
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10557 2099 10591
rect 2041 10551 2099 10557
rect 1486 10480 1492 10532
rect 1544 10520 1550 10532
rect 1688 10520 1716 10551
rect 2682 10548 2688 10600
rect 2740 10548 2746 10600
rect 4246 10548 4252 10600
rect 4304 10548 4310 10600
rect 5276 10597 5304 10628
rect 5368 10597 5396 10696
rect 5442 10684 5448 10736
rect 5500 10724 5506 10736
rect 5736 10724 5764 10764
rect 5500 10696 5764 10724
rect 5500 10684 5506 10696
rect 7742 10684 7748 10736
rect 7800 10724 7806 10736
rect 7800 10696 8800 10724
rect 7800 10684 7806 10696
rect 4985 10591 5043 10597
rect 4985 10557 4997 10591
rect 5031 10557 5043 10591
rect 4985 10551 5043 10557
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10557 5411 10591
rect 5353 10551 5411 10557
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7190 10588 7196 10600
rect 6687 10560 7196 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 1544 10492 1900 10520
rect 1544 10480 1550 10492
rect 1872 10461 1900 10492
rect 3510 10480 3516 10532
rect 3568 10520 3574 10532
rect 5000 10520 5028 10551
rect 7190 10548 7196 10560
rect 7248 10588 7254 10600
rect 7742 10588 7748 10600
rect 7248 10560 7748 10588
rect 7248 10548 7254 10560
rect 7742 10548 7748 10560
rect 7800 10548 7806 10600
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 8036 10560 8401 10588
rect 3568 10492 5028 10520
rect 5169 10523 5227 10529
rect 3568 10480 3574 10492
rect 5169 10489 5181 10523
rect 5215 10489 5227 10523
rect 5169 10483 5227 10489
rect 6908 10523 6966 10529
rect 6908 10489 6920 10523
rect 6954 10520 6966 10523
rect 7098 10520 7104 10532
rect 6954 10492 7104 10520
rect 6954 10489 6966 10492
rect 6908 10483 6966 10489
rect 1857 10455 1915 10461
rect 1857 10421 1869 10455
rect 1903 10452 1915 10455
rect 2133 10455 2191 10461
rect 2133 10452 2145 10455
rect 1903 10424 2145 10452
rect 1903 10421 1915 10424
rect 1857 10415 1915 10421
rect 2133 10421 2145 10424
rect 2179 10421 2191 10455
rect 2133 10415 2191 10421
rect 4154 10412 4160 10464
rect 4212 10452 4218 10464
rect 4522 10452 4528 10464
rect 4212 10424 4528 10452
rect 4212 10412 4218 10424
rect 4522 10412 4528 10424
rect 4580 10412 4586 10464
rect 5184 10452 5212 10483
rect 7098 10480 7104 10492
rect 7156 10480 7162 10532
rect 7926 10452 7932 10464
rect 5184 10424 7932 10452
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 8036 10461 8064 10560
rect 8389 10557 8401 10560
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 8570 10548 8576 10600
rect 8628 10548 8634 10600
rect 8772 10597 8800 10696
rect 8864 10656 8892 10764
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 9861 10795 9919 10801
rect 9861 10792 9873 10795
rect 9548 10764 9873 10792
rect 9548 10752 9554 10764
rect 9861 10761 9873 10764
rect 9907 10761 9919 10795
rect 9861 10755 9919 10761
rect 12713 10795 12771 10801
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 13170 10792 13176 10804
rect 12759 10764 13176 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 13170 10752 13176 10764
rect 13228 10792 13234 10804
rect 14277 10795 14335 10801
rect 14277 10792 14289 10795
rect 13228 10764 14289 10792
rect 13228 10752 13234 10764
rect 14277 10761 14289 10764
rect 14323 10792 14335 10795
rect 14458 10792 14464 10804
rect 14323 10764 14464 10792
rect 14323 10761 14335 10764
rect 14277 10755 14335 10761
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 14734 10752 14740 10804
rect 14792 10752 14798 10804
rect 14918 10752 14924 10804
rect 14976 10792 14982 10804
rect 15197 10795 15255 10801
rect 15197 10792 15209 10795
rect 14976 10764 15209 10792
rect 14976 10752 14982 10764
rect 15197 10761 15209 10764
rect 15243 10792 15255 10795
rect 15654 10792 15660 10804
rect 15243 10764 15660 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 16390 10792 16396 10804
rect 16080 10764 16396 10792
rect 16080 10752 16086 10764
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 16577 10795 16635 10801
rect 16577 10761 16589 10795
rect 16623 10792 16635 10795
rect 16666 10792 16672 10804
rect 16623 10764 16672 10792
rect 16623 10761 16635 10764
rect 16577 10755 16635 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 16853 10795 16911 10801
rect 16853 10761 16865 10795
rect 16899 10792 16911 10795
rect 17034 10792 17040 10804
rect 16899 10764 17040 10792
rect 16899 10761 16911 10764
rect 16853 10755 16911 10761
rect 17034 10752 17040 10764
rect 17092 10792 17098 10804
rect 17310 10792 17316 10804
rect 17092 10764 17316 10792
rect 17092 10752 17098 10764
rect 17310 10752 17316 10764
rect 17368 10792 17374 10804
rect 17497 10795 17555 10801
rect 17497 10792 17509 10795
rect 17368 10764 17509 10792
rect 17368 10752 17374 10764
rect 17497 10761 17509 10764
rect 17543 10761 17555 10795
rect 17497 10755 17555 10761
rect 17678 10752 17684 10804
rect 17736 10752 17742 10804
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10792 18383 10795
rect 18782 10792 18788 10804
rect 18371 10764 18788 10792
rect 18371 10761 18383 10764
rect 18325 10755 18383 10761
rect 18782 10752 18788 10764
rect 18840 10752 18846 10804
rect 20346 10752 20352 10804
rect 20404 10752 20410 10804
rect 21453 10795 21511 10801
rect 21453 10761 21465 10795
rect 21499 10792 21511 10795
rect 22094 10792 22100 10804
rect 21499 10764 22100 10792
rect 21499 10761 21511 10764
rect 21453 10755 21511 10761
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 25041 10795 25099 10801
rect 25041 10761 25053 10795
rect 25087 10792 25099 10795
rect 25682 10792 25688 10804
rect 25087 10764 25688 10792
rect 25087 10761 25099 10764
rect 25041 10755 25099 10761
rect 25682 10752 25688 10764
rect 25740 10752 25746 10804
rect 25958 10752 25964 10804
rect 26016 10752 26022 10804
rect 26418 10752 26424 10804
rect 26476 10752 26482 10804
rect 27246 10752 27252 10804
rect 27304 10752 27310 10804
rect 27801 10795 27859 10801
rect 27801 10761 27813 10795
rect 27847 10792 27859 10795
rect 28074 10792 28080 10804
rect 27847 10764 28080 10792
rect 27847 10761 27859 10764
rect 27801 10755 27859 10761
rect 28074 10752 28080 10764
rect 28132 10752 28138 10804
rect 28166 10752 28172 10804
rect 28224 10792 28230 10804
rect 28353 10795 28411 10801
rect 28353 10792 28365 10795
rect 28224 10764 28365 10792
rect 28224 10752 28230 10764
rect 28353 10761 28365 10764
rect 28399 10761 28411 10795
rect 28353 10755 28411 10761
rect 28721 10795 28779 10801
rect 28721 10761 28733 10795
rect 28767 10792 28779 10795
rect 28810 10792 28816 10804
rect 28767 10764 28816 10792
rect 28767 10761 28779 10764
rect 28721 10755 28779 10761
rect 28810 10752 28816 10764
rect 28868 10792 28874 10804
rect 29454 10792 29460 10804
rect 28868 10764 29460 10792
rect 28868 10752 28874 10764
rect 29454 10752 29460 10764
rect 29512 10792 29518 10804
rect 30650 10792 30656 10804
rect 29512 10764 30656 10792
rect 29512 10752 29518 10764
rect 30650 10752 30656 10764
rect 30708 10752 30714 10804
rect 9646 10696 13860 10724
rect 9646 10656 9674 10696
rect 8864 10628 9674 10656
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 10192 10628 10701 10656
rect 10192 10616 10198 10628
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 8662 10480 8668 10532
rect 8720 10480 8726 10532
rect 8772 10464 8800 10551
rect 9122 10548 9128 10600
rect 9180 10588 9186 10600
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 9180 10560 9505 10588
rect 9180 10548 9186 10560
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 9582 10548 9588 10600
rect 9640 10548 9646 10600
rect 10336 10597 10364 10628
rect 10689 10625 10701 10628
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10588 10011 10591
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 9999 10560 10333 10588
rect 9999 10557 10011 10560
rect 9953 10551 10011 10557
rect 10321 10557 10333 10560
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 10778 10548 10784 10600
rect 10836 10588 10842 10600
rect 11882 10588 11888 10600
rect 10836 10560 11888 10588
rect 10836 10548 10842 10560
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 13832 10588 13860 10696
rect 13906 10684 13912 10736
rect 13964 10724 13970 10736
rect 14752 10724 14780 10752
rect 13964 10696 14780 10724
rect 15841 10727 15899 10733
rect 13964 10684 13970 10696
rect 15841 10693 15853 10727
rect 15887 10724 15899 10727
rect 17126 10724 17132 10736
rect 15887 10696 17132 10724
rect 15887 10693 15899 10696
rect 15841 10687 15899 10693
rect 17126 10684 17132 10696
rect 17184 10684 17190 10736
rect 17696 10724 17724 10752
rect 18877 10727 18935 10733
rect 18877 10724 18889 10727
rect 17696 10696 18889 10724
rect 18877 10693 18889 10696
rect 18923 10693 18935 10727
rect 18877 10687 18935 10693
rect 25516 10696 30512 10724
rect 16114 10656 16120 10668
rect 16041 10628 16120 10656
rect 12452 10560 12664 10588
rect 13832 10560 15056 10588
rect 12452 10520 12480 10560
rect 12636 10532 12664 10560
rect 8956 10492 12480 10520
rect 8021 10455 8079 10461
rect 8021 10421 8033 10455
rect 8067 10421 8079 10455
rect 8021 10415 8079 10421
rect 8754 10412 8760 10464
rect 8812 10412 8818 10464
rect 8956 10461 8984 10492
rect 12526 10480 12532 10532
rect 12584 10480 12590 10532
rect 12618 10480 12624 10532
rect 12676 10480 12682 10532
rect 12745 10523 12803 10529
rect 12745 10489 12757 10523
rect 12791 10520 12803 10523
rect 12791 10492 14304 10520
rect 12791 10489 12803 10492
rect 12745 10483 12803 10489
rect 8941 10455 8999 10461
rect 8941 10421 8953 10455
rect 8987 10421 8999 10455
rect 8941 10415 8999 10421
rect 10226 10412 10232 10464
rect 10284 10412 10290 10464
rect 12894 10412 12900 10464
rect 12952 10412 12958 10464
rect 14090 10412 14096 10464
rect 14148 10412 14154 10464
rect 14276 10461 14304 10492
rect 14366 10480 14372 10532
rect 14424 10520 14430 10532
rect 14461 10523 14519 10529
rect 14461 10520 14473 10523
rect 14424 10492 14473 10520
rect 14424 10480 14430 10492
rect 14461 10489 14473 10492
rect 14507 10489 14519 10523
rect 14461 10483 14519 10489
rect 14550 10480 14556 10532
rect 14608 10480 14614 10532
rect 14734 10480 14740 10532
rect 14792 10529 14798 10532
rect 15028 10529 15056 10560
rect 15838 10548 15844 10600
rect 15896 10548 15902 10600
rect 15930 10548 15936 10600
rect 15988 10548 15994 10600
rect 16041 10597 16069 10628
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 16850 10616 16856 10668
rect 16908 10616 16914 10668
rect 17402 10616 17408 10668
rect 17460 10656 17466 10668
rect 17460 10628 18828 10656
rect 17460 10616 17466 10628
rect 16026 10591 16084 10597
rect 16026 10557 16038 10591
rect 16072 10557 16084 10591
rect 16301 10591 16359 10597
rect 16301 10590 16313 10591
rect 16224 10588 16313 10590
rect 16026 10551 16084 10557
rect 16132 10562 16313 10588
rect 16132 10560 16252 10562
rect 14792 10523 14811 10529
rect 14799 10489 14811 10523
rect 14792 10483 14811 10489
rect 15013 10523 15071 10529
rect 15013 10489 15025 10523
rect 15059 10489 15071 10523
rect 15013 10483 15071 10489
rect 14792 10480 14798 10483
rect 15470 10480 15476 10532
rect 15528 10480 15534 10532
rect 15856 10520 15884 10548
rect 16132 10520 16160 10560
rect 16301 10557 16313 10562
rect 16347 10557 16359 10591
rect 16301 10551 16359 10557
rect 16390 10548 16396 10600
rect 16448 10597 16454 10600
rect 16448 10588 16456 10597
rect 16868 10588 16896 10616
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 16448 10560 16493 10588
rect 16592 10560 17356 10588
rect 16448 10551 16456 10560
rect 16448 10548 16454 10551
rect 15856 10492 16160 10520
rect 16209 10523 16267 10529
rect 16209 10489 16221 10523
rect 16255 10520 16267 10523
rect 16592 10520 16620 10560
rect 16255 10492 16620 10520
rect 16255 10489 16267 10492
rect 16209 10483 16267 10489
rect 16666 10480 16672 10532
rect 16724 10480 16730 10532
rect 16885 10523 16943 10529
rect 16885 10489 16897 10523
rect 16931 10520 16943 10523
rect 16931 10492 17264 10520
rect 16931 10489 16943 10492
rect 16885 10483 16943 10489
rect 14261 10455 14319 10461
rect 14261 10421 14273 10455
rect 14307 10452 14319 10455
rect 14752 10452 14780 10480
rect 17236 10464 17264 10492
rect 17328 10464 17356 10560
rect 18356 10560 18705 10588
rect 17589 10523 17647 10529
rect 17589 10489 17601 10523
rect 17635 10489 17647 10523
rect 17589 10483 17647 10489
rect 14307 10424 14780 10452
rect 14307 10421 14319 10424
rect 14261 10415 14319 10421
rect 14918 10412 14924 10464
rect 14976 10412 14982 10464
rect 15194 10412 15200 10464
rect 15252 10461 15258 10464
rect 15252 10455 15271 10461
rect 15259 10421 15271 10455
rect 15252 10415 15271 10421
rect 15252 10412 15258 10415
rect 15378 10412 15384 10464
rect 15436 10412 15442 10464
rect 15683 10455 15741 10461
rect 15683 10421 15695 10455
rect 15729 10452 15741 10455
rect 16298 10452 16304 10464
rect 15729 10424 16304 10452
rect 15729 10421 15741 10424
rect 15683 10415 15741 10421
rect 16298 10412 16304 10424
rect 16356 10412 16362 10464
rect 17034 10412 17040 10464
rect 17092 10412 17098 10464
rect 17218 10412 17224 10464
rect 17276 10412 17282 10464
rect 17310 10412 17316 10464
rect 17368 10412 17374 10464
rect 17604 10452 17632 10483
rect 18138 10480 18144 10532
rect 18196 10480 18202 10532
rect 17770 10452 17776 10464
rect 17604 10424 17776 10452
rect 17770 10412 17776 10424
rect 17828 10452 17834 10464
rect 18356 10461 18384 10560
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18800 10588 18828 10628
rect 19242 10616 19248 10668
rect 19300 10656 19306 10668
rect 19300 10628 20213 10656
rect 19300 10616 19306 10628
rect 18800 10560 19656 10588
rect 18693 10551 18751 10557
rect 19628 10520 19656 10560
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 19794 10548 19800 10600
rect 19852 10548 19858 10600
rect 20070 10548 20076 10600
rect 20128 10548 20134 10600
rect 20185 10597 20213 10628
rect 21266 10616 21272 10668
rect 21324 10656 21330 10668
rect 21324 10628 21404 10656
rect 21324 10616 21330 10628
rect 21376 10597 21404 10628
rect 22186 10616 22192 10668
rect 22244 10656 22250 10668
rect 22281 10659 22339 10665
rect 22281 10656 22293 10659
rect 22244 10628 22293 10656
rect 22244 10616 22250 10628
rect 22281 10625 22293 10628
rect 22327 10625 22339 10659
rect 22281 10619 22339 10625
rect 20185 10591 20269 10597
rect 20185 10560 20223 10591
rect 20211 10557 20223 10560
rect 20257 10588 20269 10591
rect 21361 10591 21419 10597
rect 20257 10560 21312 10588
rect 20257 10557 20269 10560
rect 20211 10551 20269 10557
rect 19981 10523 20039 10529
rect 19981 10520 19993 10523
rect 19628 10492 19993 10520
rect 19981 10489 19993 10492
rect 20027 10489 20039 10523
rect 21284 10520 21312 10560
rect 21361 10557 21373 10591
rect 21407 10588 21419 10591
rect 21637 10591 21695 10597
rect 21637 10588 21649 10591
rect 21407 10560 21649 10588
rect 21407 10557 21419 10560
rect 21361 10551 21419 10557
rect 21637 10557 21649 10560
rect 21683 10557 21695 10591
rect 21913 10591 21971 10597
rect 21913 10588 21925 10591
rect 21637 10551 21695 10557
rect 21744 10560 21925 10588
rect 21744 10532 21772 10560
rect 21913 10557 21925 10560
rect 21959 10557 21971 10591
rect 21913 10551 21971 10557
rect 22548 10591 22606 10597
rect 22548 10557 22560 10591
rect 22594 10588 22606 10591
rect 22830 10588 22836 10600
rect 22594 10560 22836 10588
rect 22594 10557 22606 10560
rect 22548 10551 22606 10557
rect 22830 10548 22836 10560
rect 22888 10548 22894 10600
rect 25133 10591 25191 10597
rect 25133 10557 25145 10591
rect 25179 10588 25191 10591
rect 25406 10588 25412 10600
rect 25179 10560 25412 10588
rect 25179 10557 25191 10560
rect 25133 10551 25191 10557
rect 25406 10548 25412 10560
rect 25464 10588 25470 10600
rect 25516 10597 25544 10696
rect 25958 10656 25964 10668
rect 25792 10628 25964 10656
rect 25792 10597 25820 10628
rect 25958 10616 25964 10628
rect 26016 10656 26022 10668
rect 26016 10628 26648 10656
rect 26016 10616 26022 10628
rect 25501 10591 25559 10597
rect 25501 10588 25513 10591
rect 25464 10560 25513 10588
rect 25464 10548 25470 10560
rect 25501 10557 25513 10560
rect 25547 10557 25559 10591
rect 25501 10551 25559 10557
rect 25777 10591 25835 10597
rect 25777 10557 25789 10591
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 25869 10591 25927 10597
rect 25869 10557 25881 10591
rect 25915 10557 25927 10591
rect 25869 10551 25927 10557
rect 26329 10591 26387 10597
rect 26329 10557 26341 10591
rect 26375 10557 26387 10591
rect 26329 10551 26387 10557
rect 21542 10520 21548 10532
rect 21284 10492 21548 10520
rect 19981 10483 20039 10489
rect 21542 10480 21548 10492
rect 21600 10480 21606 10532
rect 21726 10480 21732 10532
rect 21784 10480 21790 10532
rect 25884 10520 25912 10551
rect 25516 10492 25912 10520
rect 25516 10464 25544 10492
rect 18346 10455 18404 10461
rect 18346 10452 18358 10455
rect 17828 10424 18358 10452
rect 17828 10412 17834 10424
rect 18346 10421 18358 10424
rect 18392 10421 18404 10455
rect 18346 10415 18404 10421
rect 18506 10412 18512 10464
rect 18564 10412 18570 10464
rect 22005 10455 22063 10461
rect 22005 10421 22017 10455
rect 22051 10452 22063 10455
rect 22186 10452 22192 10464
rect 22051 10424 22192 10452
rect 22051 10421 22063 10424
rect 22005 10415 22063 10421
rect 22186 10412 22192 10424
rect 22244 10412 22250 10464
rect 23661 10455 23719 10461
rect 23661 10421 23673 10455
rect 23707 10452 23719 10455
rect 23842 10452 23848 10464
rect 23707 10424 23848 10452
rect 23707 10421 23719 10424
rect 23661 10415 23719 10421
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 25498 10412 25504 10464
rect 25556 10412 25562 10464
rect 25682 10412 25688 10464
rect 25740 10452 25746 10464
rect 26344 10452 26372 10551
rect 26418 10548 26424 10600
rect 26476 10548 26482 10600
rect 26620 10597 26648 10628
rect 27246 10616 27252 10668
rect 27304 10656 27310 10668
rect 30374 10656 30380 10668
rect 27304 10628 28028 10656
rect 27304 10616 27310 10628
rect 26605 10591 26663 10597
rect 26605 10557 26617 10591
rect 26651 10557 26663 10591
rect 26605 10551 26663 10557
rect 26786 10548 26792 10600
rect 26844 10588 26850 10600
rect 28000 10597 28028 10628
rect 29840 10628 30380 10656
rect 27065 10591 27123 10597
rect 27065 10588 27077 10591
rect 26844 10560 27077 10588
rect 26844 10548 26850 10560
rect 27065 10557 27077 10560
rect 27111 10588 27123 10591
rect 27157 10591 27215 10597
rect 27157 10588 27169 10591
rect 27111 10560 27169 10588
rect 27111 10557 27123 10560
rect 27065 10551 27123 10557
rect 27157 10557 27169 10560
rect 27203 10557 27215 10591
rect 27157 10551 27215 10557
rect 27617 10591 27675 10597
rect 27617 10557 27629 10591
rect 27663 10588 27675 10591
rect 27709 10591 27767 10597
rect 27709 10588 27721 10591
rect 27663 10560 27721 10588
rect 27663 10557 27675 10560
rect 27617 10551 27675 10557
rect 27709 10557 27721 10560
rect 27755 10557 27767 10591
rect 27709 10551 27767 10557
rect 27985 10591 28043 10597
rect 27985 10557 27997 10591
rect 28031 10557 28043 10591
rect 27985 10551 28043 10557
rect 25740 10424 26372 10452
rect 26436 10452 26464 10548
rect 26697 10523 26755 10529
rect 26697 10489 26709 10523
rect 26743 10520 26755 10523
rect 26973 10523 27031 10529
rect 26973 10520 26985 10523
rect 26743 10492 26985 10520
rect 26743 10489 26755 10492
rect 26697 10483 26755 10489
rect 26973 10489 26985 10492
rect 27019 10520 27031 10523
rect 27632 10520 27660 10551
rect 28442 10548 28448 10600
rect 28500 10548 28506 10600
rect 28813 10591 28871 10597
rect 28813 10557 28825 10591
rect 28859 10557 28871 10591
rect 28813 10551 28871 10557
rect 27019 10492 27660 10520
rect 28828 10520 28856 10551
rect 29086 10548 29092 10600
rect 29144 10548 29150 10600
rect 29181 10591 29239 10597
rect 29181 10557 29193 10591
rect 29227 10588 29239 10591
rect 29270 10588 29276 10600
rect 29227 10560 29276 10588
rect 29227 10557 29239 10560
rect 29181 10551 29239 10557
rect 29270 10548 29276 10560
rect 29328 10588 29334 10600
rect 29840 10597 29868 10628
rect 30374 10616 30380 10628
rect 30432 10616 30438 10668
rect 30484 10665 30512 10696
rect 30469 10659 30527 10665
rect 30469 10625 30481 10659
rect 30515 10625 30527 10659
rect 30469 10619 30527 10625
rect 29365 10591 29423 10597
rect 29365 10588 29377 10591
rect 29328 10560 29377 10588
rect 29328 10548 29334 10560
rect 29365 10557 29377 10560
rect 29411 10588 29423 10591
rect 29733 10591 29791 10597
rect 29733 10588 29745 10591
rect 29411 10560 29745 10588
rect 29411 10557 29423 10560
rect 29365 10551 29423 10557
rect 29733 10557 29745 10560
rect 29779 10557 29791 10591
rect 29733 10551 29791 10557
rect 29825 10591 29883 10597
rect 29825 10557 29837 10591
rect 29871 10557 29883 10591
rect 29825 10551 29883 10557
rect 30929 10591 30987 10597
rect 30929 10557 30941 10591
rect 30975 10588 30987 10591
rect 31662 10588 31668 10600
rect 30975 10560 31668 10588
rect 30975 10557 30987 10560
rect 30929 10551 30987 10557
rect 31662 10548 31668 10560
rect 31720 10548 31726 10600
rect 28994 10520 29000 10532
rect 28828 10492 29000 10520
rect 27019 10489 27031 10492
rect 26973 10483 27031 10489
rect 28994 10480 29000 10492
rect 29052 10520 29058 10532
rect 29914 10520 29920 10532
rect 29052 10492 29920 10520
rect 29052 10480 29058 10492
rect 29914 10480 29920 10492
rect 29972 10480 29978 10532
rect 27525 10455 27583 10461
rect 27525 10452 27537 10455
rect 26436 10424 27537 10452
rect 25740 10412 25746 10424
rect 27525 10421 27537 10424
rect 27571 10421 27583 10455
rect 27525 10415 27583 10421
rect 552 10362 31531 10384
rect 552 10310 8102 10362
rect 8154 10310 8166 10362
rect 8218 10310 8230 10362
rect 8282 10310 8294 10362
rect 8346 10310 8358 10362
rect 8410 10310 15807 10362
rect 15859 10310 15871 10362
rect 15923 10310 15935 10362
rect 15987 10310 15999 10362
rect 16051 10310 16063 10362
rect 16115 10310 23512 10362
rect 23564 10310 23576 10362
rect 23628 10310 23640 10362
rect 23692 10310 23704 10362
rect 23756 10310 23768 10362
rect 23820 10310 31217 10362
rect 31269 10310 31281 10362
rect 31333 10310 31345 10362
rect 31397 10310 31409 10362
rect 31461 10310 31473 10362
rect 31525 10310 31531 10362
rect 552 10288 31531 10310
rect 1394 10248 1400 10260
rect 1228 10220 1400 10248
rect 1228 10121 1256 10220
rect 1394 10208 1400 10220
rect 1452 10208 1458 10260
rect 19613 10251 19671 10257
rect 19613 10248 19625 10251
rect 2746 10220 16160 10248
rect 1302 10140 1308 10192
rect 1360 10180 1366 10192
rect 2746 10180 2774 10220
rect 3602 10180 3608 10192
rect 1360 10152 2774 10180
rect 3344 10152 3608 10180
rect 1360 10140 1366 10152
rect 1213 10115 1271 10121
rect 1213 10081 1225 10115
rect 1259 10081 1271 10115
rect 1213 10075 1271 10081
rect 1486 10072 1492 10124
rect 1544 10072 1550 10124
rect 1670 10072 1676 10124
rect 1728 10112 1734 10124
rect 3344 10121 3372 10152
rect 3602 10140 3608 10152
rect 3660 10140 3666 10192
rect 3694 10140 3700 10192
rect 3752 10180 3758 10192
rect 3752 10152 4016 10180
rect 3752 10140 3758 10152
rect 1857 10115 1915 10121
rect 1857 10112 1869 10115
rect 1728 10084 1869 10112
rect 1728 10072 1734 10084
rect 1857 10081 1869 10084
rect 1903 10081 1915 10115
rect 2113 10115 2171 10121
rect 2113 10112 2125 10115
rect 1857 10075 1915 10081
rect 1964 10084 2125 10112
rect 1964 10044 1992 10084
rect 2113 10081 2125 10084
rect 2159 10081 2171 10115
rect 2113 10075 2171 10081
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10081 3387 10115
rect 3329 10075 3387 10081
rect 3421 10115 3479 10121
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 3786 10112 3792 10124
rect 3467 10084 3792 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 3786 10072 3792 10084
rect 3844 10112 3850 10124
rect 3881 10115 3939 10121
rect 3881 10112 3893 10115
rect 3844 10084 3893 10112
rect 3844 10072 3850 10084
rect 3881 10081 3893 10084
rect 3927 10081 3939 10115
rect 3881 10075 3939 10081
rect 1596 10016 1992 10044
rect 3988 10044 4016 10152
rect 4246 10140 4252 10192
rect 4304 10180 4310 10192
rect 4525 10183 4583 10189
rect 4525 10180 4537 10183
rect 4304 10152 4537 10180
rect 4304 10140 4310 10152
rect 4525 10149 4537 10152
rect 4571 10180 4583 10183
rect 4801 10183 4859 10189
rect 4801 10180 4813 10183
rect 4571 10152 4813 10180
rect 4571 10149 4583 10152
rect 4525 10143 4583 10149
rect 4801 10149 4813 10152
rect 4847 10149 4859 10183
rect 7466 10180 7472 10192
rect 4801 10143 4859 10149
rect 7208 10152 7472 10180
rect 4157 10115 4215 10121
rect 4157 10081 4169 10115
rect 4203 10112 4215 10115
rect 4264 10112 4292 10140
rect 4203 10084 4292 10112
rect 4433 10115 4491 10121
rect 4203 10081 4215 10084
rect 4157 10075 4215 10081
rect 4433 10081 4445 10115
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 4062 10044 4068 10056
rect 3988 10016 4068 10044
rect 1596 9920 1624 10016
rect 4062 10004 4068 10016
rect 4120 10044 4126 10056
rect 4448 10044 4476 10075
rect 4706 10072 4712 10124
rect 4764 10072 4770 10124
rect 7208 10121 7236 10152
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 7834 10180 7840 10192
rect 7668 10152 7840 10180
rect 7668 10121 7696 10152
rect 7834 10140 7840 10152
rect 7892 10140 7898 10192
rect 9582 10189 9588 10192
rect 9576 10143 9588 10189
rect 9582 10140 9588 10143
rect 9640 10140 9646 10192
rect 13357 10183 13415 10189
rect 13357 10180 13369 10183
rect 10704 10152 13369 10180
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7653 10115 7711 10121
rect 7653 10081 7665 10115
rect 7699 10081 7711 10115
rect 7653 10075 7711 10081
rect 7742 10072 7748 10124
rect 7800 10112 7806 10124
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 7800 10084 9321 10112
rect 7800 10072 7806 10084
rect 9309 10081 9321 10084
rect 9355 10081 9367 10115
rect 9309 10075 9367 10081
rect 8662 10044 8668 10056
rect 4120 10016 4476 10044
rect 5092 10016 8668 10044
rect 4120 10004 4126 10016
rect 3973 9979 4031 9985
rect 3973 9945 3985 9979
rect 4019 9976 4031 9979
rect 4154 9976 4160 9988
rect 4019 9948 4160 9976
rect 4019 9945 4031 9948
rect 3973 9939 4031 9945
rect 4154 9936 4160 9948
rect 4212 9936 4218 9988
rect 4249 9979 4307 9985
rect 4249 9945 4261 9979
rect 4295 9976 4307 9979
rect 4982 9976 4988 9988
rect 4295 9948 4988 9976
rect 4295 9945 4307 9948
rect 4249 9939 4307 9945
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 1210 9868 1216 9920
rect 1268 9908 1274 9920
rect 1305 9911 1363 9917
rect 1305 9908 1317 9911
rect 1268 9880 1317 9908
rect 1268 9868 1274 9880
rect 1305 9877 1317 9880
rect 1351 9877 1363 9911
rect 1305 9871 1363 9877
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 3237 9911 3295 9917
rect 3237 9877 3249 9911
rect 3283 9908 3295 9911
rect 5092 9908 5120 10016
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 10704 9985 10732 10152
rect 13357 10149 13369 10152
rect 13403 10149 13415 10183
rect 13357 10143 13415 10149
rect 13573 10183 13631 10189
rect 13573 10149 13585 10183
rect 13619 10180 13631 10183
rect 13906 10180 13912 10192
rect 13619 10152 13912 10180
rect 13619 10149 13631 10152
rect 13573 10143 13631 10149
rect 13906 10140 13912 10152
rect 13964 10140 13970 10192
rect 16132 10189 16160 10220
rect 17328 10220 19625 10248
rect 16117 10183 16175 10189
rect 14568 10152 15884 10180
rect 11790 10072 11796 10124
rect 11848 10112 11854 10124
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11848 10084 11897 10112
rect 11848 10072 11854 10084
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 11974 10072 11980 10124
rect 12032 10112 12038 10124
rect 12141 10115 12199 10121
rect 12141 10112 12153 10115
rect 12032 10084 12153 10112
rect 12032 10072 12038 10084
rect 12141 10081 12153 10084
rect 12187 10081 12199 10115
rect 12141 10075 12199 10081
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 14001 10115 14059 10121
rect 14001 10112 14013 10115
rect 13780 10084 14013 10112
rect 13780 10072 13786 10084
rect 14001 10081 14013 10084
rect 14047 10081 14059 10115
rect 14001 10075 14059 10081
rect 14182 10072 14188 10124
rect 14240 10072 14246 10124
rect 14274 10072 14280 10124
rect 14332 10072 14338 10124
rect 10689 9979 10747 9985
rect 10689 9945 10701 9979
rect 10735 9945 10747 9979
rect 10689 9939 10747 9945
rect 13262 9936 13268 9988
rect 13320 9936 13326 9988
rect 14568 9920 14596 10152
rect 15381 10115 15439 10121
rect 15381 10081 15393 10115
rect 15427 10081 15439 10115
rect 15381 10075 15439 10081
rect 14734 10004 14740 10056
rect 14792 10044 14798 10056
rect 15105 10047 15163 10053
rect 15105 10044 15117 10047
rect 14792 10016 15117 10044
rect 14792 10004 14798 10016
rect 15105 10013 15117 10016
rect 15151 10013 15163 10047
rect 15105 10007 15163 10013
rect 15197 10047 15255 10053
rect 15197 10013 15209 10047
rect 15243 10044 15255 10047
rect 15286 10044 15292 10056
rect 15243 10016 15292 10044
rect 15243 10013 15255 10016
rect 15197 10007 15255 10013
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 15396 10044 15424 10075
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 15746 10112 15752 10124
rect 15620 10084 15752 10112
rect 15620 10072 15626 10084
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 15856 10112 15884 10152
rect 16117 10149 16129 10183
rect 16163 10149 16175 10183
rect 16117 10143 16175 10149
rect 16942 10112 16948 10124
rect 15856 10084 16948 10112
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 17328 10044 17356 10220
rect 19613 10217 19625 10220
rect 19659 10217 19671 10251
rect 19613 10211 19671 10217
rect 21266 10208 21272 10260
rect 21324 10248 21330 10260
rect 21545 10251 21603 10257
rect 21545 10248 21557 10251
rect 21324 10220 21557 10248
rect 21324 10208 21330 10220
rect 21545 10217 21557 10220
rect 21591 10217 21603 10251
rect 21545 10211 21603 10217
rect 21821 10251 21879 10257
rect 21821 10217 21833 10251
rect 21867 10248 21879 10251
rect 22002 10248 22008 10260
rect 21867 10220 22008 10248
rect 21867 10217 21879 10220
rect 21821 10211 21879 10217
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 22094 10208 22100 10260
rect 22152 10248 22158 10260
rect 22738 10248 22744 10260
rect 22152 10220 22744 10248
rect 22152 10208 22158 10220
rect 22738 10208 22744 10220
rect 22796 10208 22802 10260
rect 22830 10208 22836 10260
rect 22888 10248 22894 10260
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 22888 10220 22937 10248
rect 22888 10208 22894 10220
rect 22925 10217 22937 10220
rect 22971 10217 22983 10251
rect 22925 10211 22983 10217
rect 23842 10208 23848 10260
rect 23900 10208 23906 10260
rect 25682 10208 25688 10260
rect 25740 10208 25746 10260
rect 26878 10208 26884 10260
rect 26936 10208 26942 10260
rect 29270 10208 29276 10260
rect 29328 10208 29334 10260
rect 30374 10208 30380 10260
rect 30432 10248 30438 10260
rect 30929 10251 30987 10257
rect 30929 10248 30941 10251
rect 30432 10220 30941 10248
rect 30432 10208 30438 10220
rect 30929 10217 30941 10220
rect 30975 10217 30987 10251
rect 30929 10211 30987 10217
rect 20438 10180 20444 10192
rect 15396 10016 17356 10044
rect 17420 10152 20444 10180
rect 17420 9985 17448 10152
rect 20438 10140 20444 10152
rect 20496 10180 20502 10192
rect 21910 10180 21916 10192
rect 20496 10152 21916 10180
rect 20496 10140 20502 10152
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 22373 10183 22431 10189
rect 22373 10180 22385 10183
rect 22020 10152 22385 10180
rect 17954 10072 17960 10124
rect 18012 10072 18018 10124
rect 18141 10115 18199 10121
rect 18141 10081 18153 10115
rect 18187 10081 18199 10115
rect 18141 10075 18199 10081
rect 17405 9979 17463 9985
rect 17405 9976 17417 9979
rect 14660 9948 17417 9976
rect 14660 9920 14688 9948
rect 17405 9945 17417 9948
rect 17451 9945 17463 9979
rect 17405 9939 17463 9945
rect 3283 9880 5120 9908
rect 7285 9911 7343 9917
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 7285 9877 7297 9911
rect 7331 9908 7343 9911
rect 7558 9908 7564 9920
rect 7331 9880 7564 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 13538 9868 13544 9920
rect 13596 9868 13602 9920
rect 13722 9868 13728 9920
rect 13780 9868 13786 9920
rect 14090 9868 14096 9920
rect 14148 9908 14154 9920
rect 14369 9911 14427 9917
rect 14369 9908 14381 9911
rect 14148 9880 14381 9908
rect 14148 9868 14154 9880
rect 14369 9877 14381 9880
rect 14415 9877 14427 9911
rect 14369 9871 14427 9877
rect 14461 9911 14519 9917
rect 14461 9877 14473 9911
rect 14507 9908 14519 9911
rect 14550 9908 14556 9920
rect 14507 9880 14556 9908
rect 14507 9877 14519 9880
rect 14461 9871 14519 9877
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 14642 9868 14648 9920
rect 14700 9868 14706 9920
rect 14734 9868 14740 9920
rect 14792 9868 14798 9920
rect 14826 9868 14832 9920
rect 14884 9868 14890 9920
rect 15289 9911 15347 9917
rect 15289 9877 15301 9911
rect 15335 9908 15347 9911
rect 15378 9908 15384 9920
rect 15335 9880 15384 9908
rect 15335 9877 15347 9880
rect 15289 9871 15347 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 18156 9908 18184 10075
rect 18322 10072 18328 10124
rect 18380 10072 18386 10124
rect 18693 10115 18751 10121
rect 18693 10081 18705 10115
rect 18739 10081 18751 10115
rect 18693 10075 18751 10081
rect 18946 10115 19004 10121
rect 18946 10081 18958 10115
rect 18992 10112 19004 10115
rect 19521 10115 19579 10121
rect 18992 10084 19334 10112
rect 18992 10081 19004 10084
rect 18946 10075 19004 10081
rect 18230 10004 18236 10056
rect 18288 10044 18294 10056
rect 18708 10044 18736 10075
rect 18288 10016 18920 10044
rect 18288 10004 18294 10016
rect 18892 9988 18920 10016
rect 18874 9936 18880 9988
rect 18932 9936 18938 9988
rect 16632 9880 18184 9908
rect 19306 9908 19334 10084
rect 19521 10081 19533 10115
rect 19567 10112 19579 10115
rect 19978 10112 19984 10124
rect 19567 10084 19984 10112
rect 19567 10081 19579 10084
rect 19521 10075 19579 10081
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 20737 10115 20795 10121
rect 20737 10081 20749 10115
rect 20783 10112 20795 10115
rect 20783 10084 20944 10112
rect 20783 10081 20795 10084
rect 20737 10075 20795 10081
rect 20916 10044 20944 10084
rect 20990 10072 20996 10124
rect 21048 10072 21054 10124
rect 21634 10072 21640 10124
rect 21692 10072 21698 10124
rect 21726 10072 21732 10124
rect 21784 10112 21790 10124
rect 22020 10112 22048 10152
rect 22373 10149 22385 10152
rect 22419 10149 22431 10183
rect 22373 10143 22431 10149
rect 21784 10084 22048 10112
rect 21784 10072 21790 10084
rect 22186 10072 22192 10124
rect 22244 10072 22250 10124
rect 22278 10072 22284 10124
rect 22336 10072 22342 10124
rect 22554 10072 22560 10124
rect 22612 10072 22618 10124
rect 22756 10112 22784 10208
rect 23584 10152 24532 10180
rect 23584 10121 23612 10152
rect 24504 10124 24532 10152
rect 25498 10140 25504 10192
rect 25556 10140 25562 10192
rect 22833 10115 22891 10121
rect 22833 10112 22845 10115
rect 22756 10084 22845 10112
rect 22833 10081 22845 10084
rect 22879 10081 22891 10115
rect 22833 10075 22891 10081
rect 23569 10115 23627 10121
rect 23569 10081 23581 10115
rect 23615 10081 23627 10115
rect 23569 10075 23627 10081
rect 23937 10115 23995 10121
rect 23937 10081 23949 10115
rect 23983 10081 23995 10115
rect 23937 10075 23995 10081
rect 20916 10016 21680 10044
rect 21542 9936 21548 9988
rect 21600 9936 21606 9988
rect 21560 9908 21588 9936
rect 19306 9880 21588 9908
rect 21652 9908 21680 10016
rect 22204 9908 22232 10072
rect 23382 10004 23388 10056
rect 23440 10044 23446 10056
rect 23952 10044 23980 10075
rect 24486 10072 24492 10124
rect 24544 10072 24550 10124
rect 25406 10072 25412 10124
rect 25464 10072 25470 10124
rect 25700 10112 25728 10208
rect 27982 10140 27988 10192
rect 28040 10189 28046 10192
rect 28040 10180 28052 10189
rect 28902 10180 28908 10192
rect 28040 10152 28085 10180
rect 28736 10152 28908 10180
rect 28040 10143 28052 10152
rect 28040 10140 28046 10143
rect 28736 10121 28764 10152
rect 28902 10140 28908 10152
rect 28960 10140 28966 10192
rect 25777 10115 25835 10121
rect 25777 10112 25789 10115
rect 25700 10084 25789 10112
rect 25777 10081 25789 10084
rect 25823 10081 25835 10115
rect 25777 10075 25835 10081
rect 28721 10115 28779 10121
rect 28721 10081 28733 10115
rect 28767 10081 28779 10115
rect 28721 10075 28779 10081
rect 28810 10072 28816 10124
rect 28868 10072 28874 10124
rect 29288 10121 29316 10208
rect 29632 10183 29690 10189
rect 29632 10149 29644 10183
rect 29678 10180 29690 10183
rect 30282 10180 30288 10192
rect 29678 10152 30288 10180
rect 29678 10149 29690 10152
rect 29632 10143 29690 10149
rect 30282 10140 30288 10152
rect 30340 10140 30346 10192
rect 29273 10115 29331 10121
rect 29273 10081 29285 10115
rect 29319 10081 29331 10115
rect 29273 10075 29331 10081
rect 29914 10072 29920 10124
rect 29972 10112 29978 10124
rect 30837 10115 30895 10121
rect 30837 10112 30849 10115
rect 29972 10084 30849 10112
rect 29972 10072 29978 10084
rect 30837 10081 30849 10084
rect 30883 10081 30895 10115
rect 30837 10075 30895 10081
rect 23440 10016 23980 10044
rect 23440 10004 23446 10016
rect 25590 10004 25596 10056
rect 25648 10044 25654 10056
rect 25685 10047 25743 10053
rect 25685 10044 25697 10047
rect 25648 10016 25697 10044
rect 25648 10004 25654 10016
rect 25685 10013 25697 10016
rect 25731 10013 25743 10047
rect 25685 10007 25743 10013
rect 28261 10047 28319 10053
rect 28261 10013 28273 10047
rect 28307 10044 28319 10047
rect 29362 10044 29368 10056
rect 28307 10016 29368 10044
rect 28307 10013 28319 10016
rect 28261 10007 28319 10013
rect 29362 10004 29368 10016
rect 29420 10004 29426 10056
rect 23198 9936 23204 9988
rect 23256 9936 23262 9988
rect 23477 9979 23535 9985
rect 23477 9945 23489 9979
rect 23523 9976 23535 9979
rect 24026 9976 24032 9988
rect 23523 9948 24032 9976
rect 23523 9945 23535 9948
rect 23477 9939 23535 9945
rect 24026 9936 24032 9948
rect 24084 9936 24090 9988
rect 24826 9948 25820 9976
rect 22649 9911 22707 9917
rect 22649 9908 22661 9911
rect 21652 9880 22661 9908
rect 16632 9868 16638 9880
rect 22649 9877 22661 9880
rect 22695 9877 22707 9911
rect 22649 9871 22707 9877
rect 23661 9911 23719 9917
rect 23661 9877 23673 9911
rect 23707 9908 23719 9911
rect 23842 9908 23848 9920
rect 23707 9880 23848 9908
rect 23707 9877 23719 9880
rect 23661 9871 23719 9877
rect 23842 9868 23848 9880
rect 23900 9868 23906 9920
rect 24394 9868 24400 9920
rect 24452 9908 24458 9920
rect 24826 9908 24854 9948
rect 24452 9880 24854 9908
rect 25792 9908 25820 9948
rect 28276 9948 29316 9976
rect 28276 9908 28304 9948
rect 25792 9880 28304 9908
rect 28629 9911 28687 9917
rect 24452 9868 24458 9880
rect 28629 9877 28641 9911
rect 28675 9908 28687 9911
rect 29178 9908 29184 9920
rect 28675 9880 29184 9908
rect 28675 9877 28687 9880
rect 28629 9871 28687 9877
rect 29178 9868 29184 9880
rect 29236 9868 29242 9920
rect 29288 9908 29316 9948
rect 30745 9911 30803 9917
rect 30745 9908 30757 9911
rect 29288 9880 30757 9908
rect 30745 9877 30757 9880
rect 30791 9877 30803 9911
rect 30745 9871 30803 9877
rect 552 9818 31372 9840
rect 552 9766 4250 9818
rect 4302 9766 4314 9818
rect 4366 9766 4378 9818
rect 4430 9766 4442 9818
rect 4494 9766 4506 9818
rect 4558 9766 11955 9818
rect 12007 9766 12019 9818
rect 12071 9766 12083 9818
rect 12135 9766 12147 9818
rect 12199 9766 12211 9818
rect 12263 9766 19660 9818
rect 19712 9766 19724 9818
rect 19776 9766 19788 9818
rect 19840 9766 19852 9818
rect 19904 9766 19916 9818
rect 19968 9766 27365 9818
rect 27417 9766 27429 9818
rect 27481 9766 27493 9818
rect 27545 9766 27557 9818
rect 27609 9766 27621 9818
rect 27673 9766 31372 9818
rect 552 9744 31372 9766
rect 1578 9664 1584 9716
rect 1636 9704 1642 9716
rect 1857 9707 1915 9713
rect 1857 9704 1869 9707
rect 1636 9676 1869 9704
rect 1636 9664 1642 9676
rect 1857 9673 1869 9676
rect 1903 9673 1915 9707
rect 1857 9667 1915 9673
rect 1762 9596 1768 9648
rect 1820 9596 1826 9648
rect 1872 9636 1900 9667
rect 3786 9664 3792 9716
rect 3844 9664 3850 9716
rect 4062 9664 4068 9716
rect 4120 9664 4126 9716
rect 4341 9707 4399 9713
rect 4341 9673 4353 9707
rect 4387 9704 4399 9707
rect 4706 9704 4712 9716
rect 4387 9676 4712 9704
rect 4387 9673 4399 9676
rect 4341 9667 4399 9673
rect 1872 9608 2360 9636
rect 1210 9528 1216 9580
rect 1268 9528 1274 9580
rect 1780 9568 1808 9596
rect 1688 9540 1900 9568
rect 1228 9500 1256 9528
rect 1688 9509 1716 9540
rect 1397 9503 1455 9509
rect 1397 9500 1409 9503
rect 1228 9472 1409 9500
rect 1397 9469 1409 9472
rect 1443 9500 1455 9503
rect 1581 9503 1639 9509
rect 1581 9500 1593 9503
rect 1443 9472 1593 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1581 9469 1593 9472
rect 1627 9469 1639 9503
rect 1581 9463 1639 9469
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9469 1731 9503
rect 1673 9463 1731 9469
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9469 1823 9503
rect 1872 9500 1900 9540
rect 2332 9509 2360 9608
rect 4356 9568 4384 9667
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 8754 9664 8760 9716
rect 8812 9704 8818 9716
rect 12526 9704 12532 9716
rect 8812 9676 12532 9704
rect 8812 9664 8818 9676
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 13722 9664 13728 9716
rect 13780 9664 13786 9716
rect 13817 9707 13875 9713
rect 13817 9673 13829 9707
rect 13863 9704 13875 9707
rect 13906 9704 13912 9716
rect 13863 9676 13912 9704
rect 13863 9673 13875 9676
rect 13817 9667 13875 9673
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 14642 9664 14648 9716
rect 14700 9664 14706 9716
rect 14826 9704 14832 9716
rect 14768 9676 14832 9704
rect 7561 9639 7619 9645
rect 7561 9636 7573 9639
rect 3896 9540 4384 9568
rect 7116 9608 7573 9636
rect 2041 9503 2099 9509
rect 2041 9500 2053 9503
rect 1872 9472 2053 9500
rect 1765 9463 1823 9469
rect 2041 9469 2053 9472
rect 2087 9469 2099 9503
rect 2041 9463 2099 9469
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9469 2375 9503
rect 2317 9463 2375 9469
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9500 3571 9503
rect 3602 9500 3608 9512
rect 3559 9472 3608 9500
rect 3559 9469 3571 9472
rect 3513 9463 3571 9469
rect 1596 9432 1624 9463
rect 1780 9432 1808 9463
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 3896 9509 3924 9540
rect 7116 9512 7144 9608
rect 7561 9605 7573 9608
rect 7607 9605 7619 9639
rect 12805 9639 12863 9645
rect 12805 9636 12817 9639
rect 7561 9599 7619 9605
rect 11880 9608 12817 9636
rect 7852 9540 8524 9568
rect 7852 9512 7880 9540
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3844 9472 3893 9500
rect 3844 9460 3850 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 3881 9463 3939 9469
rect 3988 9472 4169 9500
rect 3988 9432 4016 9472
rect 4157 9469 4169 9472
rect 4203 9500 4215 9503
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 4203 9472 4261 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 4908 9432 4936 9463
rect 4982 9460 4988 9512
rect 5040 9500 5046 9512
rect 5149 9503 5207 9509
rect 5149 9500 5161 9503
rect 5040 9472 5161 9500
rect 5040 9460 5046 9472
rect 5149 9469 5161 9472
rect 5195 9469 5207 9503
rect 5149 9463 5207 9469
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6871 9472 6929 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 6917 9469 6929 9472
rect 6963 9500 6975 9503
rect 7098 9500 7104 9512
rect 6963 9472 7104 9500
rect 6963 9469 6975 9472
rect 6917 9463 6975 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7377 9503 7435 9509
rect 7377 9469 7389 9503
rect 7423 9500 7435 9503
rect 7466 9500 7472 9512
rect 7423 9472 7472 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7558 9460 7564 9512
rect 7616 9500 7622 9512
rect 7653 9503 7711 9509
rect 7653 9500 7665 9503
rect 7616 9472 7665 9500
rect 7616 9460 7622 9472
rect 7653 9469 7665 9472
rect 7699 9500 7711 9503
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7699 9472 7757 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 7834 9460 7840 9512
rect 7892 9460 7898 9512
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9469 8447 9503
rect 8496 9500 8524 9540
rect 8645 9503 8703 9509
rect 8645 9500 8657 9503
rect 8496 9472 8657 9500
rect 8389 9463 8447 9469
rect 8645 9469 8657 9472
rect 8691 9469 8703 9503
rect 8645 9463 8703 9469
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9500 10931 9503
rect 10962 9500 10968 9512
rect 10919 9472 10968 9500
rect 10919 9469 10931 9472
rect 10873 9463 10931 9469
rect 8036 9432 8064 9463
rect 1596 9404 1808 9432
rect 3436 9404 4016 9432
rect 4172 9404 4936 9432
rect 7300 9404 8064 9432
rect 8404 9432 8432 9463
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 11140 9503 11198 9509
rect 11140 9469 11152 9503
rect 11186 9500 11198 9503
rect 11606 9500 11612 9512
rect 11186 9472 11612 9500
rect 11186 9469 11198 9472
rect 11140 9463 11198 9469
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 11698 9460 11704 9512
rect 11756 9500 11762 9512
rect 11880 9500 11908 9608
rect 12805 9605 12817 9608
rect 12851 9605 12863 9639
rect 13740 9636 13768 9664
rect 14001 9639 14059 9645
rect 14001 9636 14013 9639
rect 13740 9608 14013 9636
rect 12805 9599 12863 9605
rect 14001 9605 14013 9608
rect 14047 9605 14059 9639
rect 14001 9599 14059 9605
rect 12250 9528 12256 9580
rect 12308 9568 12314 9580
rect 12621 9571 12679 9577
rect 12621 9568 12633 9571
rect 12308 9540 12633 9568
rect 12308 9528 12314 9540
rect 12621 9537 12633 9540
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 14768 9577 14796 9676
rect 14826 9664 14832 9676
rect 14884 9664 14890 9716
rect 14918 9664 14924 9716
rect 14976 9664 14982 9716
rect 15102 9664 15108 9716
rect 15160 9664 15166 9716
rect 16574 9664 16580 9716
rect 16632 9664 16638 9716
rect 16669 9707 16727 9713
rect 16669 9673 16681 9707
rect 16715 9704 16727 9707
rect 16850 9704 16856 9716
rect 16715 9676 16856 9704
rect 16715 9673 16727 9676
rect 16669 9667 16727 9673
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 16945 9707 17003 9713
rect 16945 9673 16957 9707
rect 16991 9704 17003 9707
rect 17034 9704 17040 9716
rect 16991 9676 17040 9704
rect 16991 9673 17003 9676
rect 16945 9667 17003 9673
rect 17034 9664 17040 9676
rect 17092 9664 17098 9716
rect 17126 9664 17132 9716
rect 17184 9664 17190 9716
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 17497 9707 17555 9713
rect 17497 9704 17509 9707
rect 17276 9676 17509 9704
rect 17276 9664 17282 9676
rect 17497 9673 17509 9676
rect 17543 9673 17555 9707
rect 17497 9667 17555 9673
rect 17586 9664 17592 9716
rect 17644 9704 17650 9716
rect 19153 9707 19211 9713
rect 19153 9704 19165 9707
rect 17644 9676 19165 9704
rect 17644 9664 17650 9676
rect 19153 9673 19165 9676
rect 19199 9673 19211 9707
rect 20530 9704 20536 9716
rect 19153 9667 19211 9673
rect 20180 9676 20536 9704
rect 14936 9636 14964 9664
rect 15565 9639 15623 9645
rect 14936 9608 15516 9636
rect 13909 9571 13967 9577
rect 13909 9568 13921 9571
rect 13228 9540 13921 9568
rect 13228 9528 13234 9540
rect 13909 9537 13921 9540
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 14737 9571 14796 9577
rect 14737 9537 14749 9571
rect 14783 9540 14796 9571
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 15102 9528 15108 9580
rect 15160 9568 15166 9580
rect 15197 9571 15255 9577
rect 15197 9568 15209 9571
rect 15160 9540 15209 9568
rect 15160 9528 15166 9540
rect 15197 9537 15209 9540
rect 15243 9537 15255 9571
rect 15488 9568 15516 9608
rect 15565 9605 15577 9639
rect 15611 9636 15623 9639
rect 18230 9636 18236 9648
rect 15611 9608 17540 9636
rect 15611 9605 15623 9608
rect 15565 9599 15623 9605
rect 15488 9540 16160 9568
rect 15197 9531 15255 9537
rect 12342 9500 12348 9512
rect 11756 9472 11908 9500
rect 11992 9472 12348 9500
rect 11756 9460 11762 9472
rect 11882 9432 11888 9444
rect 8404 9404 8524 9432
rect 1305 9367 1363 9373
rect 1305 9333 1317 9367
rect 1351 9364 1363 9367
rect 1394 9364 1400 9376
rect 1351 9336 1400 9364
rect 1351 9333 1363 9336
rect 1305 9327 1363 9333
rect 1394 9324 1400 9336
rect 1452 9324 1458 9376
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 2409 9367 2467 9373
rect 2409 9364 2421 9367
rect 2188 9336 2421 9364
rect 2188 9324 2194 9336
rect 2409 9333 2421 9336
rect 2455 9333 2467 9367
rect 2409 9327 2467 9333
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 3436 9373 3464 9404
rect 4172 9376 4200 9404
rect 3421 9367 3479 9373
rect 3421 9364 3433 9367
rect 3292 9336 3433 9364
rect 3292 9324 3298 9336
rect 3421 9333 3433 9336
rect 3467 9333 3479 9367
rect 3421 9327 3479 9333
rect 4154 9324 4160 9376
rect 4212 9324 4218 9376
rect 6270 9324 6276 9376
rect 6328 9324 6334 9376
rect 6730 9324 6736 9376
rect 6788 9324 6794 9376
rect 7300 9373 7328 9404
rect 7668 9376 7696 9404
rect 8496 9376 8524 9404
rect 9784 9404 11888 9432
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9364 7067 9367
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 7055 9336 7297 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7285 9327 7343 9333
rect 7650 9324 7656 9376
rect 7708 9324 7714 9376
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 8113 9367 8171 9373
rect 8113 9364 8125 9367
rect 7892 9336 8125 9364
rect 7892 9324 7898 9336
rect 8113 9333 8125 9336
rect 8159 9333 8171 9367
rect 8113 9327 8171 9333
rect 8478 9324 8484 9376
rect 8536 9324 8542 9376
rect 9784 9373 9812 9404
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9333 9827 9367
rect 9769 9327 9827 9333
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 11992 9364 12020 9472
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 12710 9460 12716 9512
rect 12768 9460 12774 9512
rect 13446 9460 13452 9512
rect 13504 9500 13510 9512
rect 13541 9503 13599 9509
rect 13541 9500 13553 9503
rect 13504 9472 13553 9500
rect 13504 9460 13510 9472
rect 13541 9469 13553 9472
rect 13587 9500 13599 9503
rect 13587 9472 14796 9500
rect 13587 9469 13599 9472
rect 13541 9463 13599 9469
rect 12066 9392 12072 9444
rect 12124 9432 12130 9444
rect 13081 9435 13139 9441
rect 12124 9404 12572 9432
rect 12124 9392 12130 9404
rect 11388 9336 12020 9364
rect 12253 9367 12311 9373
rect 11388 9324 11394 9336
rect 12253 9333 12265 9367
rect 12299 9364 12311 9367
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 12299 9336 12449 9364
rect 12299 9333 12311 9336
rect 12253 9327 12311 9333
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12544 9364 12572 9404
rect 13081 9401 13093 9435
rect 13127 9432 13139 9435
rect 14553 9435 14611 9441
rect 14553 9432 14565 9435
rect 13127 9404 14565 9432
rect 13127 9401 13139 9404
rect 13081 9395 13139 9401
rect 14553 9401 14565 9404
rect 14599 9401 14611 9435
rect 14768 9432 14796 9472
rect 14826 9460 14832 9512
rect 14884 9460 14890 9512
rect 14927 9472 15332 9500
rect 14927 9432 14955 9472
rect 14768 9404 14955 9432
rect 15105 9435 15163 9441
rect 14553 9395 14611 9401
rect 15105 9401 15117 9435
rect 15151 9432 15163 9435
rect 15194 9432 15200 9444
rect 15151 9404 15200 9432
rect 15151 9401 15163 9404
rect 15105 9395 15163 9401
rect 15194 9392 15200 9404
rect 15252 9392 15258 9444
rect 15304 9432 15332 9472
rect 15378 9460 15384 9512
rect 15436 9460 15442 9512
rect 15654 9460 15660 9512
rect 15712 9500 15718 9512
rect 15940 9503 15998 9509
rect 15940 9502 15952 9503
rect 15856 9500 15952 9502
rect 15712 9474 15952 9500
rect 15712 9472 15884 9474
rect 15712 9460 15718 9472
rect 15940 9469 15952 9474
rect 15986 9469 15998 9503
rect 15940 9463 15998 9469
rect 16026 9503 16084 9509
rect 16026 9469 16038 9503
rect 16072 9469 16084 9503
rect 16132 9500 16160 9540
rect 16868 9540 17264 9568
rect 16298 9503 16356 9509
rect 16298 9500 16310 9503
rect 16132 9472 16310 9500
rect 16026 9463 16084 9469
rect 16298 9469 16310 9472
rect 16344 9469 16356 9503
rect 16298 9463 16356 9469
rect 15746 9432 15752 9444
rect 15304 9404 15752 9432
rect 15746 9392 15752 9404
rect 15804 9392 15810 9444
rect 16041 9432 16069 9463
rect 16390 9460 16396 9512
rect 16448 9509 16454 9512
rect 16448 9503 16475 9509
rect 16463 9469 16475 9503
rect 16448 9463 16475 9469
rect 16448 9460 16454 9463
rect 16114 9432 16120 9444
rect 16041 9404 16120 9432
rect 16114 9392 16120 9404
rect 16172 9392 16178 9444
rect 16209 9435 16267 9441
rect 16209 9401 16221 9435
rect 16255 9401 16267 9435
rect 16209 9395 16267 9401
rect 13633 9367 13691 9373
rect 13633 9364 13645 9367
rect 12544 9336 13645 9364
rect 12437 9327 12495 9333
rect 13633 9333 13645 9336
rect 13679 9333 13691 9367
rect 13633 9327 13691 9333
rect 14277 9367 14335 9373
rect 14277 9333 14289 9367
rect 14323 9364 14335 9367
rect 14734 9364 14740 9376
rect 14323 9336 14740 9364
rect 14323 9333 14335 9336
rect 14277 9327 14335 9333
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 14826 9324 14832 9376
rect 14884 9364 14890 9376
rect 15013 9367 15071 9373
rect 15013 9364 15025 9367
rect 14884 9336 15025 9364
rect 14884 9324 14890 9336
rect 15013 9333 15025 9336
rect 15059 9333 15071 9367
rect 16224 9364 16252 9395
rect 16868 9376 16896 9540
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 17037 9503 17095 9509
rect 17037 9500 17049 9503
rect 17000 9472 17049 9500
rect 17000 9460 17006 9472
rect 17037 9469 17049 9472
rect 17083 9500 17095 9503
rect 17126 9500 17132 9512
rect 17083 9472 17132 9500
rect 17083 9469 17095 9472
rect 17037 9463 17095 9469
rect 17126 9460 17132 9472
rect 17184 9460 17190 9512
rect 17236 9494 17264 9540
rect 17405 9503 17463 9509
rect 17405 9494 17417 9503
rect 17236 9469 17417 9494
rect 17451 9469 17463 9503
rect 17236 9466 17463 9469
rect 17405 9463 17463 9466
rect 16850 9364 16856 9376
rect 16224 9336 16856 9364
rect 15013 9327 15071 9333
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 17310 9373 17316 9376
rect 17267 9367 17316 9373
rect 17267 9333 17279 9367
rect 17313 9333 17316 9367
rect 17267 9327 17316 9333
rect 17310 9324 17316 9327
rect 17368 9324 17374 9376
rect 17512 9364 17540 9608
rect 17696 9608 18236 9636
rect 17696 9509 17724 9608
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 18506 9596 18512 9648
rect 18564 9596 18570 9648
rect 19518 9596 19524 9648
rect 19576 9636 19582 9648
rect 19613 9639 19671 9645
rect 19613 9636 19625 9639
rect 19576 9608 19625 9636
rect 19576 9596 19582 9608
rect 19613 9605 19625 9608
rect 19659 9605 19671 9639
rect 19613 9599 19671 9605
rect 19702 9596 19708 9648
rect 19760 9636 19766 9648
rect 20180 9636 20208 9676
rect 20530 9664 20536 9676
rect 20588 9704 20594 9716
rect 20588 9676 20944 9704
rect 20588 9664 20594 9676
rect 20806 9636 20812 9648
rect 19760 9608 20208 9636
rect 20272 9608 20812 9636
rect 19760 9596 19766 9608
rect 18524 9568 18552 9596
rect 20165 9571 20223 9577
rect 20165 9568 20177 9571
rect 18524 9540 20177 9568
rect 20165 9537 20177 9540
rect 20211 9537 20223 9571
rect 20165 9531 20223 9537
rect 17681 9503 17739 9509
rect 17773 9506 17831 9509
rect 17681 9469 17693 9503
rect 17727 9469 17739 9503
rect 17681 9463 17739 9469
rect 17770 9454 17776 9506
rect 17828 9500 17834 9506
rect 17828 9472 17867 9500
rect 17828 9454 17834 9472
rect 19334 9460 19340 9512
rect 19392 9460 19398 9512
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 19705 9503 19763 9509
rect 19705 9500 19717 9503
rect 19475 9472 19717 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 19705 9469 19717 9472
rect 19751 9469 19763 9503
rect 19705 9463 19763 9469
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9469 20039 9503
rect 19981 9463 20039 9469
rect 18322 9392 18328 9444
rect 18380 9392 18386 9444
rect 19153 9435 19211 9441
rect 19153 9401 19165 9435
rect 19199 9401 19211 9435
rect 19153 9395 19211 9401
rect 18340 9364 18368 9392
rect 17512 9336 18368 9364
rect 19168 9364 19196 9395
rect 19518 9392 19524 9444
rect 19576 9432 19582 9444
rect 19996 9432 20024 9463
rect 20070 9460 20076 9512
rect 20128 9460 20134 9512
rect 20272 9509 20300 9608
rect 20806 9596 20812 9608
rect 20864 9596 20870 9648
rect 20916 9568 20944 9676
rect 21266 9664 21272 9716
rect 21324 9664 21330 9716
rect 21634 9664 21640 9716
rect 21692 9704 21698 9716
rect 22097 9707 22155 9713
rect 22097 9704 22109 9707
rect 21692 9676 22109 9704
rect 21692 9664 21698 9676
rect 22097 9673 22109 9676
rect 22143 9704 22155 9707
rect 22554 9704 22560 9716
rect 22143 9676 22560 9704
rect 22143 9673 22155 9676
rect 22097 9667 22155 9673
rect 22554 9664 22560 9676
rect 22612 9704 22618 9716
rect 22649 9707 22707 9713
rect 22649 9704 22661 9707
rect 22612 9676 22661 9704
rect 22612 9664 22618 9676
rect 22649 9673 22661 9676
rect 22695 9673 22707 9707
rect 22649 9667 22707 9673
rect 28902 9664 28908 9716
rect 28960 9704 28966 9716
rect 30009 9707 30067 9713
rect 30009 9704 30021 9707
rect 28960 9676 30021 9704
rect 28960 9664 28966 9676
rect 21177 9639 21235 9645
rect 21177 9605 21189 9639
rect 21223 9605 21235 9639
rect 21284 9636 21312 9664
rect 21821 9639 21879 9645
rect 21821 9636 21833 9639
rect 21284 9608 21833 9636
rect 21177 9599 21235 9605
rect 21821 9605 21833 9608
rect 21867 9605 21879 9639
rect 21821 9599 21879 9605
rect 21192 9568 21220 9599
rect 29086 9596 29092 9648
rect 29144 9636 29150 9648
rect 29641 9639 29699 9645
rect 29641 9636 29653 9639
rect 29144 9608 29653 9636
rect 29144 9596 29150 9608
rect 29641 9605 29653 9608
rect 29687 9605 29699 9639
rect 29641 9599 29699 9605
rect 20916 9540 21036 9568
rect 21192 9540 24348 9568
rect 20257 9503 20315 9509
rect 20257 9469 20269 9503
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 20438 9460 20444 9512
rect 20496 9460 20502 9512
rect 20530 9460 20536 9512
rect 20588 9460 20594 9512
rect 20626 9503 20684 9509
rect 20626 9469 20638 9503
rect 20672 9469 20684 9503
rect 20626 9463 20684 9469
rect 19576 9404 20024 9432
rect 19576 9392 19582 9404
rect 20346 9392 20352 9444
rect 20404 9432 20410 9444
rect 20631 9432 20659 9463
rect 20898 9460 20904 9512
rect 20956 9460 20962 9512
rect 21008 9509 21036 9540
rect 20998 9503 21056 9509
rect 20998 9469 21010 9503
rect 21044 9469 21056 9503
rect 20998 9463 21056 9469
rect 21913 9503 21971 9509
rect 21913 9469 21925 9503
rect 21959 9500 21971 9503
rect 21959 9472 22094 9500
rect 21959 9469 21971 9472
rect 21913 9463 21971 9469
rect 22066 9444 22094 9472
rect 22186 9460 22192 9512
rect 22244 9460 22250 9512
rect 22281 9503 22339 9509
rect 22281 9469 22293 9503
rect 22327 9469 22339 9503
rect 22281 9463 22339 9469
rect 20404 9404 20659 9432
rect 20809 9435 20867 9441
rect 20404 9392 20410 9404
rect 20809 9401 20821 9435
rect 20855 9432 20867 9435
rect 21082 9432 21088 9444
rect 20855 9404 21088 9432
rect 20855 9401 20867 9404
rect 20809 9395 20867 9401
rect 21082 9392 21088 9404
rect 21140 9392 21146 9444
rect 21744 9404 21956 9432
rect 22066 9404 22100 9444
rect 21744 9364 21772 9404
rect 19168 9336 21772 9364
rect 21928 9364 21956 9404
rect 22094 9392 22100 9404
rect 22152 9432 22158 9444
rect 22296 9432 22324 9463
rect 22462 9460 22468 9512
rect 22520 9460 22526 9512
rect 22554 9460 22560 9512
rect 22612 9460 22618 9512
rect 24118 9460 24124 9512
rect 24176 9460 24182 9512
rect 24320 9509 24348 9540
rect 25682 9528 25688 9580
rect 25740 9528 25746 9580
rect 24305 9503 24363 9509
rect 24305 9469 24317 9503
rect 24351 9469 24363 9503
rect 24305 9463 24363 9469
rect 24486 9460 24492 9512
rect 24544 9460 24550 9512
rect 24670 9460 24676 9512
rect 24728 9500 24734 9512
rect 24857 9503 24915 9509
rect 24857 9500 24869 9503
rect 24728 9472 24869 9500
rect 24728 9460 24734 9472
rect 24857 9469 24869 9472
rect 24903 9469 24915 9503
rect 24857 9463 24915 9469
rect 25110 9503 25168 9509
rect 25110 9469 25122 9503
rect 25156 9500 25168 9503
rect 27157 9503 27215 9509
rect 25156 9472 25820 9500
rect 25156 9469 25168 9472
rect 25110 9463 25168 9469
rect 22152 9404 22324 9432
rect 22480 9432 22508 9460
rect 24578 9432 24584 9444
rect 22480 9404 24584 9432
rect 22152 9392 22158 9404
rect 24578 9392 24584 9404
rect 24636 9392 24642 9444
rect 22278 9364 22284 9376
rect 21928 9336 22284 9364
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 22370 9324 22376 9376
rect 22428 9324 22434 9376
rect 25792 9373 25820 9472
rect 27157 9469 27169 9503
rect 27203 9500 27215 9503
rect 27890 9500 27896 9512
rect 27203 9472 27896 9500
rect 27203 9469 27215 9472
rect 27157 9463 27215 9469
rect 27890 9460 27896 9472
rect 27948 9460 27954 9512
rect 29181 9503 29239 9509
rect 29181 9469 29193 9503
rect 29227 9500 29239 9503
rect 29227 9472 29408 9500
rect 29227 9469 29239 9472
rect 29181 9463 29239 9469
rect 26786 9392 26792 9444
rect 26844 9432 26850 9444
rect 29380 9441 29408 9472
rect 29454 9460 29460 9512
rect 29512 9460 29518 9512
rect 29733 9503 29791 9509
rect 29733 9469 29745 9503
rect 29779 9500 29791 9503
rect 29932 9500 29960 9676
rect 30009 9673 30021 9676
rect 30055 9673 30067 9707
rect 30009 9667 30067 9673
rect 30282 9664 30288 9716
rect 30340 9664 30346 9716
rect 30561 9571 30619 9577
rect 30561 9568 30573 9571
rect 29779 9472 29960 9500
rect 30024 9540 30573 9568
rect 29779 9469 29791 9472
rect 29733 9463 29791 9469
rect 26890 9435 26948 9441
rect 26890 9432 26902 9435
rect 26844 9404 26902 9432
rect 26844 9392 26850 9404
rect 26890 9401 26902 9404
rect 26936 9401 26948 9435
rect 26890 9395 26948 9401
rect 29365 9435 29423 9441
rect 29365 9401 29377 9435
rect 29411 9432 29423 9435
rect 30024 9432 30052 9540
rect 30101 9503 30159 9509
rect 30101 9469 30113 9503
rect 30147 9500 30159 9503
rect 30282 9500 30288 9512
rect 30147 9472 30288 9500
rect 30147 9469 30159 9472
rect 30101 9463 30159 9469
rect 30282 9460 30288 9472
rect 30340 9460 30346 9512
rect 30392 9509 30420 9540
rect 30561 9537 30573 9540
rect 30607 9537 30619 9571
rect 30561 9531 30619 9537
rect 30377 9503 30435 9509
rect 30377 9469 30389 9503
rect 30423 9469 30435 9503
rect 30377 9463 30435 9469
rect 30469 9503 30527 9509
rect 30469 9469 30481 9503
rect 30515 9469 30527 9503
rect 30469 9463 30527 9469
rect 30484 9432 30512 9463
rect 29411 9404 30052 9432
rect 30208 9404 30512 9432
rect 29411 9401 29423 9404
rect 29365 9395 29423 9401
rect 25777 9367 25835 9373
rect 25777 9333 25789 9367
rect 25823 9333 25835 9367
rect 25777 9327 25835 9333
rect 29178 9324 29184 9376
rect 29236 9364 29242 9376
rect 30208 9364 30236 9404
rect 29236 9336 30236 9364
rect 29236 9324 29242 9336
rect 552 9274 31531 9296
rect 552 9222 8102 9274
rect 8154 9222 8166 9274
rect 8218 9222 8230 9274
rect 8282 9222 8294 9274
rect 8346 9222 8358 9274
rect 8410 9222 15807 9274
rect 15859 9222 15871 9274
rect 15923 9222 15935 9274
rect 15987 9222 15999 9274
rect 16051 9222 16063 9274
rect 16115 9222 23512 9274
rect 23564 9222 23576 9274
rect 23628 9222 23640 9274
rect 23692 9222 23704 9274
rect 23756 9222 23768 9274
rect 23820 9222 31217 9274
rect 31269 9222 31281 9274
rect 31333 9222 31345 9274
rect 31397 9222 31409 9274
rect 31461 9222 31473 9274
rect 31525 9222 31531 9274
rect 552 9200 31531 9222
rect 1305 9163 1363 9169
rect 1305 9129 1317 9163
rect 1351 9160 1363 9163
rect 1394 9160 1400 9172
rect 1351 9132 1400 9160
rect 1351 9129 1363 9132
rect 1305 9123 1363 9129
rect 1394 9120 1400 9132
rect 1452 9120 1458 9172
rect 2130 9120 2136 9172
rect 2188 9120 2194 9172
rect 3234 9120 3240 9172
rect 3292 9120 3298 9172
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 3789 9163 3847 9169
rect 3789 9160 3801 9163
rect 3660 9132 3801 9160
rect 3660 9120 3666 9132
rect 3789 9129 3801 9132
rect 3835 9129 3847 9163
rect 3789 9123 3847 9129
rect 5629 9163 5687 9169
rect 5629 9129 5641 9163
rect 5675 9129 5687 9163
rect 5629 9123 5687 9129
rect 2148 9092 2176 9120
rect 1412 9064 2176 9092
rect 2685 9095 2743 9101
rect 1412 9033 1440 9064
rect 1121 9027 1179 9033
rect 1121 8993 1133 9027
rect 1167 8993 1179 9027
rect 1121 8987 1179 8993
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 1136 8956 1164 8987
rect 1670 8984 1676 9036
rect 1728 8984 1734 9036
rect 1964 9033 1992 9064
rect 2685 9061 2697 9095
rect 2731 9092 2743 9095
rect 3620 9092 3648 9120
rect 2731 9064 3648 9092
rect 5644 9092 5672 9123
rect 6270 9120 6276 9172
rect 6328 9160 6334 9172
rect 10229 9163 10287 9169
rect 6328 9132 9352 9160
rect 6328 9120 6334 9132
rect 6638 9092 6644 9104
rect 5644 9064 6644 9092
rect 2731 9061 2743 9064
rect 2685 9055 2743 9061
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 7285 9095 7343 9101
rect 7285 9092 7297 9095
rect 6788 9064 7297 9092
rect 6788 9052 6794 9064
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 8993 2007 9027
rect 1949 8987 2007 8993
rect 2133 9027 2191 9033
rect 2133 8993 2145 9027
rect 2179 8993 2191 9027
rect 2133 8987 2191 8993
rect 2225 9027 2283 9033
rect 2225 8993 2237 9027
rect 2271 9024 2283 9027
rect 2590 9024 2596 9036
rect 2271 8996 2596 9024
rect 2271 8993 2283 8996
rect 2225 8987 2283 8993
rect 1578 8956 1584 8968
rect 1136 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 2148 8956 2176 8987
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 2869 9027 2927 9033
rect 2869 8993 2881 9027
rect 2915 9024 2927 9027
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 2915 8996 3157 9024
rect 2915 8993 2927 8996
rect 2869 8987 2927 8993
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 3421 9027 3479 9033
rect 3421 8993 3433 9027
rect 3467 9024 3479 9027
rect 3881 9027 3939 9033
rect 3881 9024 3893 9027
rect 3467 8996 3893 9024
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 3881 8993 3893 8996
rect 3927 9024 3939 9027
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3927 8996 4077 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 4065 8993 4077 8996
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 4157 9027 4215 9033
rect 4157 8993 4169 9027
rect 4203 9024 4215 9027
rect 4505 9027 4563 9033
rect 4505 9024 4517 9027
rect 4203 8996 4517 9024
rect 4203 8993 4215 8996
rect 4157 8987 4215 8993
rect 4505 8993 4517 8996
rect 4551 8993 4563 9027
rect 4505 8987 4563 8993
rect 1872 8928 2176 8956
rect 1872 8897 1900 8928
rect 1029 8891 1087 8897
rect 1029 8857 1041 8891
rect 1075 8888 1087 8891
rect 1857 8891 1915 8897
rect 1857 8888 1869 8891
rect 1075 8860 1869 8888
rect 1075 8857 1087 8860
rect 1029 8851 1087 8857
rect 1857 8857 1869 8860
rect 1903 8857 1915 8891
rect 2148 8888 2176 8928
rect 2406 8916 2412 8968
rect 2464 8956 2470 8968
rect 2884 8956 2912 8987
rect 2464 8928 2912 8956
rect 2961 8959 3019 8965
rect 2464 8916 2470 8928
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3436 8956 3464 8987
rect 3007 8928 3464 8956
rect 3513 8959 3571 8965
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3513 8925 3525 8959
rect 3559 8956 3571 8959
rect 3786 8956 3792 8968
rect 3559 8928 3792 8956
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4172 8956 4200 8987
rect 4080 8928 4200 8956
rect 4249 8959 4307 8965
rect 4080 8888 4108 8928
rect 4249 8925 4261 8959
rect 4295 8925 4307 8959
rect 7024 8956 7052 9064
rect 7285 9061 7297 9064
rect 7331 9061 7343 9095
rect 7834 9092 7840 9104
rect 7285 9055 7343 9061
rect 7392 9064 7840 9092
rect 7392 9033 7420 9064
rect 7834 9052 7840 9064
rect 7892 9092 7898 9104
rect 9094 9095 9152 9101
rect 9094 9092 9106 9095
rect 7892 9064 9106 9092
rect 7892 9052 7898 9064
rect 9094 9061 9106 9064
rect 9140 9061 9152 9095
rect 9094 9055 9152 9061
rect 7101 9027 7159 9033
rect 7101 8993 7113 9027
rect 7147 9024 7159 9027
rect 7377 9027 7435 9033
rect 7377 9024 7389 9027
rect 7147 8996 7389 9024
rect 7147 8993 7159 8996
rect 7101 8987 7159 8993
rect 7377 8993 7389 8996
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 7650 8984 7656 9036
rect 7708 8984 7714 9036
rect 7745 9027 7803 9033
rect 7745 8993 7757 9027
rect 7791 8993 7803 9027
rect 9324 9024 9352 9132
rect 10229 9129 10241 9163
rect 10275 9160 10287 9163
rect 11517 9163 11575 9169
rect 10275 9132 11192 9160
rect 10275 9129 10287 9132
rect 10229 9123 10287 9129
rect 11164 9101 11192 9132
rect 11517 9129 11529 9163
rect 11563 9160 11575 9163
rect 12710 9160 12716 9172
rect 11563 9132 12716 9160
rect 11563 9129 11575 9132
rect 11517 9123 11575 9129
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 14182 9120 14188 9172
rect 14240 9160 14246 9172
rect 14550 9160 14556 9172
rect 14240 9132 14556 9160
rect 14240 9120 14246 9132
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 14918 9120 14924 9172
rect 14976 9160 14982 9172
rect 15013 9163 15071 9169
rect 15013 9160 15025 9163
rect 14976 9132 15025 9160
rect 14976 9120 14982 9132
rect 15013 9129 15025 9132
rect 15059 9129 15071 9163
rect 15013 9123 15071 9129
rect 15378 9120 15384 9172
rect 15436 9120 15442 9172
rect 16114 9120 16120 9172
rect 16172 9160 16178 9172
rect 16172 9132 16344 9160
rect 16172 9120 16178 9132
rect 11149 9095 11207 9101
rect 11149 9061 11161 9095
rect 11195 9061 11207 9095
rect 11149 9055 11207 9061
rect 11365 9095 11423 9101
rect 11365 9061 11377 9095
rect 11411 9092 11423 9095
rect 14369 9095 14427 9101
rect 11411 9064 11652 9092
rect 11411 9061 11423 9064
rect 11365 9055 11423 9061
rect 11624 9036 11652 9064
rect 11880 9064 13400 9092
rect 9324 8996 11284 9024
rect 7745 8987 7803 8993
rect 7466 8956 7472 8968
rect 7024 8928 7472 8956
rect 4249 8919 4307 8925
rect 4264 8888 4292 8919
rect 7466 8916 7472 8928
rect 7524 8956 7530 8968
rect 7760 8956 7788 8987
rect 8849 8959 8907 8965
rect 8849 8956 8861 8959
rect 7524 8928 7788 8956
rect 8404 8928 8861 8956
rect 7524 8916 7530 8928
rect 2148 8860 4108 8888
rect 4172 8860 4292 8888
rect 1857 8851 1915 8857
rect 4172 8832 4200 8860
rect 8404 8832 8432 8928
rect 8849 8925 8861 8928
rect 8895 8925 8907 8959
rect 11256 8956 11284 8996
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 11793 9027 11851 9033
rect 11793 9024 11805 9027
rect 11664 8996 11805 9024
rect 11664 8984 11670 8996
rect 11793 8993 11805 8996
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 11880 8956 11908 9064
rect 12986 8984 12992 9036
rect 13044 8984 13050 9036
rect 13078 8984 13084 9036
rect 13136 9024 13142 9036
rect 13173 9027 13231 9033
rect 13173 9024 13185 9027
rect 13136 8996 13185 9024
rect 13136 8984 13142 8996
rect 13173 8993 13185 8996
rect 13219 8993 13231 9027
rect 13173 8987 13231 8993
rect 13262 8984 13268 9036
rect 13320 8984 13326 9036
rect 13372 9024 13400 9064
rect 14369 9061 14381 9095
rect 14415 9092 14427 9095
rect 15396 9092 15424 9120
rect 14415 9064 15424 9092
rect 14415 9061 14427 9064
rect 14369 9055 14427 9061
rect 13372 8996 14412 9024
rect 11256 8928 11908 8956
rect 11977 8959 12035 8965
rect 8849 8919 8907 8925
rect 11977 8925 11989 8959
rect 12023 8925 12035 8959
rect 14384 8956 14412 8996
rect 14550 8984 14556 9036
rect 14608 9024 14614 9036
rect 14645 9027 14703 9033
rect 14645 9024 14657 9027
rect 14608 8996 14657 9024
rect 14608 8984 14614 8996
rect 14645 8993 14657 8996
rect 14691 8993 14703 9027
rect 14645 8987 14703 8993
rect 15105 9027 15163 9033
rect 15105 8993 15117 9027
rect 15151 9024 15163 9027
rect 16114 9024 16120 9036
rect 15151 8996 16120 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 16316 9033 16344 9132
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 19702 9160 19708 9172
rect 16868 9132 19708 9160
rect 16393 9095 16451 9101
rect 16393 9061 16405 9095
rect 16439 9061 16451 9095
rect 16684 9092 16712 9120
rect 16684 9064 16804 9092
rect 16393 9055 16451 9061
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 8993 16359 9027
rect 16301 8987 16359 8993
rect 15470 8956 15476 8968
rect 14384 8928 15476 8956
rect 11977 8919 12035 8925
rect 11609 8891 11667 8897
rect 11609 8888 11621 8891
rect 9784 8860 11621 8888
rect 4154 8780 4160 8832
rect 4212 8780 4218 8832
rect 7006 8780 7012 8832
rect 7064 8780 7070 8832
rect 7561 8823 7619 8829
rect 7561 8789 7573 8823
rect 7607 8820 7619 8823
rect 7834 8820 7840 8832
rect 7607 8792 7840 8820
rect 7607 8789 7619 8792
rect 7561 8783 7619 8789
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8386 8780 8392 8832
rect 8444 8780 8450 8832
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 9784 8820 9812 8860
rect 11609 8857 11621 8860
rect 11655 8857 11667 8891
rect 11609 8851 11667 8857
rect 8628 8792 9812 8820
rect 11333 8823 11391 8829
rect 8628 8780 8634 8792
rect 11333 8789 11345 8823
rect 11379 8820 11391 8823
rect 11514 8820 11520 8832
rect 11379 8792 11520 8820
rect 11379 8789 11391 8792
rect 11333 8783 11391 8789
rect 11514 8780 11520 8792
rect 11572 8820 11578 8832
rect 11992 8820 12020 8919
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 15654 8916 15660 8968
rect 15712 8956 15718 8968
rect 15712 8928 16160 8956
rect 15712 8916 15718 8928
rect 13446 8848 13452 8900
rect 13504 8848 13510 8900
rect 13538 8848 13544 8900
rect 13596 8888 13602 8900
rect 14737 8891 14795 8897
rect 14737 8888 14749 8891
rect 13596 8860 14749 8888
rect 13596 8848 13602 8860
rect 14737 8857 14749 8860
rect 14783 8857 14795 8891
rect 14737 8851 14795 8857
rect 14829 8891 14887 8897
rect 14829 8857 14841 8891
rect 14875 8888 14887 8891
rect 15194 8888 15200 8900
rect 14875 8860 15200 8888
rect 14875 8857 14887 8860
rect 14829 8851 14887 8857
rect 15194 8848 15200 8860
rect 15252 8848 15258 8900
rect 16132 8897 16160 8928
rect 16117 8891 16175 8897
rect 16117 8857 16129 8891
rect 16163 8857 16175 8891
rect 16117 8851 16175 8857
rect 16298 8848 16304 8900
rect 16356 8888 16362 8900
rect 16408 8888 16436 9055
rect 16776 9033 16804 9064
rect 16485 9027 16543 9033
rect 16485 8993 16497 9027
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 16623 9027 16681 9033
rect 16623 8993 16635 9027
rect 16669 8993 16681 9027
rect 16623 8987 16681 8993
rect 16761 9027 16819 9033
rect 16761 8993 16773 9027
rect 16807 8993 16819 9027
rect 16761 8987 16819 8993
rect 16356 8860 16436 8888
rect 16500 8888 16528 8987
rect 16638 8956 16666 8987
rect 16868 8956 16896 9132
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 20530 9120 20536 9172
rect 20588 9120 20594 9172
rect 21913 9163 21971 9169
rect 21913 9129 21925 9163
rect 21959 9160 21971 9163
rect 22094 9160 22100 9172
rect 21959 9132 22100 9160
rect 21959 9129 21971 9132
rect 21913 9123 21971 9129
rect 22094 9120 22100 9132
rect 22152 9160 22158 9172
rect 22189 9163 22247 9169
rect 22189 9160 22201 9163
rect 22152 9132 22201 9160
rect 22152 9120 22158 9132
rect 22189 9129 22201 9132
rect 22235 9129 22247 9163
rect 22189 9123 22247 9129
rect 23845 9163 23903 9169
rect 23845 9129 23857 9163
rect 23891 9160 23903 9163
rect 24581 9163 24639 9169
rect 24581 9160 24593 9163
rect 23891 9132 24593 9160
rect 23891 9129 23903 9132
rect 23845 9123 23903 9129
rect 24581 9129 24593 9132
rect 24627 9129 24639 9163
rect 24581 9123 24639 9129
rect 24854 9120 24860 9172
rect 24912 9160 24918 9172
rect 25015 9163 25073 9169
rect 25015 9160 25027 9163
rect 24912 9132 25027 9160
rect 24912 9120 24918 9132
rect 25015 9129 25027 9132
rect 25061 9160 25073 9163
rect 25475 9163 25533 9169
rect 25475 9160 25487 9163
rect 25061 9132 25487 9160
rect 25061 9129 25073 9132
rect 25015 9123 25073 9129
rect 25475 9129 25487 9132
rect 25521 9129 25533 9163
rect 25475 9123 25533 9129
rect 26513 9163 26571 9169
rect 26513 9129 26525 9163
rect 26559 9129 26571 9163
rect 26513 9123 26571 9129
rect 17586 9092 17592 9104
rect 17144 9064 17592 9092
rect 16942 8984 16948 9036
rect 17000 9024 17006 9036
rect 17144 9033 17172 9064
rect 17586 9052 17592 9064
rect 17644 9052 17650 9104
rect 17972 9064 18276 9092
rect 17129 9027 17187 9033
rect 17129 9024 17141 9027
rect 17000 8996 17141 9024
rect 17000 8984 17006 8996
rect 17129 8993 17141 8996
rect 17175 8993 17187 9027
rect 17972 9024 18000 9064
rect 17129 8987 17187 8993
rect 17236 8996 18000 9024
rect 16638 8928 16896 8956
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17236 8956 17264 8996
rect 18046 8984 18052 9036
rect 18104 8984 18110 9036
rect 18138 8984 18144 9036
rect 18196 8984 18202 9036
rect 18248 9033 18276 9064
rect 18322 9052 18328 9104
rect 18380 9092 18386 9104
rect 18506 9101 18512 9104
rect 18493 9095 18512 9101
rect 18493 9092 18505 9095
rect 18380 9064 18505 9092
rect 18380 9052 18386 9064
rect 18493 9061 18505 9064
rect 18493 9055 18512 9061
rect 18506 9052 18512 9055
rect 18564 9052 18570 9104
rect 18690 9052 18696 9104
rect 18748 9052 18754 9104
rect 19978 9052 19984 9104
rect 20036 9101 20042 9104
rect 20036 9095 20085 9101
rect 20036 9061 20039 9095
rect 20073 9061 20085 9095
rect 20036 9055 20085 9061
rect 20165 9095 20223 9101
rect 20165 9061 20177 9095
rect 20211 9092 20223 9095
rect 24118 9092 24124 9104
rect 20211 9064 24124 9092
rect 20211 9061 20223 9064
rect 20165 9055 20223 9061
rect 20036 9052 20042 9055
rect 24118 9052 24124 9064
rect 24176 9052 24182 9104
rect 25225 9095 25283 9101
rect 25225 9061 25237 9095
rect 25271 9061 25283 9095
rect 25225 9055 25283 9061
rect 25685 9095 25743 9101
rect 25685 9061 25697 9095
rect 25731 9092 25743 9095
rect 26528 9092 26556 9123
rect 29362 9120 29368 9172
rect 29420 9120 29426 9172
rect 30926 9120 30932 9172
rect 30984 9120 30990 9172
rect 29380 9092 29408 9120
rect 25731 9064 26556 9092
rect 27908 9064 29592 9092
rect 25731 9061 25743 9064
rect 25685 9055 25743 9061
rect 18233 9027 18291 9033
rect 18233 8993 18245 9027
rect 18279 8993 18291 9027
rect 20257 9027 20315 9033
rect 20257 9024 20269 9027
rect 18233 8987 18291 8993
rect 18616 8996 20269 9024
rect 17092 8928 17264 8956
rect 17497 8959 17555 8965
rect 17092 8916 17098 8928
rect 17497 8925 17509 8959
rect 17543 8956 17555 8959
rect 17954 8956 17960 8968
rect 17543 8928 17960 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 18156 8956 18184 8984
rect 18322 8956 18328 8968
rect 18156 8928 18328 8956
rect 18322 8916 18328 8928
rect 18380 8956 18386 8968
rect 18616 8956 18644 8996
rect 20257 8993 20269 8996
rect 20303 8993 20315 9027
rect 20257 8987 20315 8993
rect 20349 9027 20407 9033
rect 20349 8993 20361 9027
rect 20395 9024 20407 9027
rect 20622 9024 20628 9036
rect 20395 8996 20628 9024
rect 20395 8993 20407 8996
rect 20349 8987 20407 8993
rect 18380 8928 18644 8956
rect 18380 8916 18386 8928
rect 18690 8916 18696 8968
rect 18748 8956 18754 8968
rect 19889 8959 19947 8965
rect 19889 8956 19901 8959
rect 18748 8928 19901 8956
rect 18748 8916 18754 8928
rect 19889 8925 19901 8928
rect 19935 8925 19947 8959
rect 19889 8919 19947 8925
rect 16574 8888 16580 8900
rect 16500 8860 16580 8888
rect 16356 8848 16362 8860
rect 16574 8848 16580 8860
rect 16632 8848 16638 8900
rect 20272 8888 20300 8987
rect 20456 8968 20484 8996
rect 20622 8984 20628 8996
rect 20680 8984 20686 9036
rect 22005 9027 22063 9033
rect 22005 8993 22017 9027
rect 22051 8993 22063 9027
rect 22005 8987 22063 8993
rect 20438 8916 20444 8968
rect 20496 8916 20502 8968
rect 22020 8956 22048 8987
rect 22094 8984 22100 9036
rect 22152 8984 22158 9036
rect 22554 9024 22560 9036
rect 22388 8996 22560 9024
rect 22020 8928 22232 8956
rect 22002 8888 22008 8900
rect 16960 8860 19334 8888
rect 20272 8860 22008 8888
rect 12710 8820 12716 8832
rect 11572 8792 12716 8820
rect 11572 8780 11578 8792
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 13265 8823 13323 8829
rect 13265 8789 13277 8823
rect 13311 8820 13323 8823
rect 14274 8820 14280 8832
rect 13311 8792 14280 8820
rect 13311 8789 13323 8792
rect 13265 8783 13323 8789
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 14918 8780 14924 8832
rect 14976 8820 14982 8832
rect 16960 8820 16988 8860
rect 14976 8792 16988 8820
rect 14976 8780 14982 8792
rect 17034 8780 17040 8832
rect 17092 8820 17098 8832
rect 17313 8823 17371 8829
rect 17313 8820 17325 8823
rect 17092 8792 17325 8820
rect 17092 8780 17098 8792
rect 17313 8789 17325 8792
rect 17359 8789 17371 8823
rect 17313 8783 17371 8789
rect 17402 8780 17408 8832
rect 17460 8820 17466 8832
rect 17586 8820 17592 8832
rect 17460 8792 17592 8820
rect 17460 8780 17466 8792
rect 17586 8780 17592 8792
rect 17644 8820 17650 8832
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 17644 8792 17785 8820
rect 17644 8780 17650 8792
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 17773 8783 17831 8789
rect 17862 8780 17868 8832
rect 17920 8780 17926 8832
rect 17957 8823 18015 8829
rect 17957 8789 17969 8823
rect 18003 8820 18015 8823
rect 18325 8823 18383 8829
rect 18325 8820 18337 8823
rect 18003 8792 18337 8820
rect 18003 8789 18015 8792
rect 17957 8783 18015 8789
rect 18325 8789 18337 8792
rect 18371 8789 18383 8823
rect 18325 8783 18383 8789
rect 18506 8780 18512 8832
rect 18564 8820 18570 8832
rect 19058 8820 19064 8832
rect 18564 8792 19064 8820
rect 18564 8780 18570 8792
rect 19058 8780 19064 8792
rect 19116 8780 19122 8832
rect 19306 8820 19334 8860
rect 22002 8848 22008 8860
rect 22060 8848 22066 8900
rect 22204 8888 22232 8928
rect 22388 8888 22416 8996
rect 22554 8984 22560 8996
rect 22612 9024 22618 9036
rect 22721 9027 22779 9033
rect 22721 9024 22733 9027
rect 22612 8996 22733 9024
rect 22612 8984 22618 8996
rect 22721 8993 22733 8996
rect 22767 8993 22779 9027
rect 22721 8987 22779 8993
rect 23474 8984 23480 9036
rect 23532 9024 23538 9036
rect 23934 9024 23940 9036
rect 23532 8996 23940 9024
rect 23532 8984 23538 8996
rect 23934 8984 23940 8996
rect 23992 8984 23998 9036
rect 24394 8984 24400 9036
rect 24452 9024 24458 9036
rect 24673 9027 24731 9033
rect 24673 9024 24685 9027
rect 24452 8996 24685 9024
rect 24452 8984 24458 8996
rect 24673 8993 24685 8996
rect 24719 8993 24731 9027
rect 25240 9024 25268 9055
rect 27908 9036 27936 9064
rect 26510 9024 26516 9036
rect 25240 8996 26516 9024
rect 24673 8987 24731 8993
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 27637 9027 27695 9033
rect 27637 8993 27649 9027
rect 27683 9024 27695 9027
rect 27683 8996 27844 9024
rect 27683 8993 27695 8996
rect 27637 8987 27695 8993
rect 22462 8916 22468 8968
rect 22520 8916 22526 8968
rect 23952 8956 23980 8984
rect 27816 8956 27844 8996
rect 27890 8984 27896 9036
rect 27948 8984 27954 9036
rect 28353 9027 28411 9033
rect 28353 8993 28365 9027
rect 28399 9024 28411 9027
rect 28718 9024 28724 9036
rect 28399 8996 28724 9024
rect 28399 8993 28411 8996
rect 28353 8987 28411 8993
rect 28368 8956 28396 8987
rect 28718 8984 28724 8996
rect 28776 8984 28782 9036
rect 28813 9030 28871 9033
rect 28813 9027 29040 9030
rect 28813 8993 28825 9027
rect 28859 9002 29040 9027
rect 28859 8993 28871 9002
rect 28813 8987 28871 8993
rect 23952 8928 24854 8956
rect 27816 8928 28396 8956
rect 22204 8860 22416 8888
rect 23658 8848 23664 8900
rect 23716 8888 23722 8900
rect 24213 8891 24271 8897
rect 24213 8888 24225 8891
rect 23716 8860 24225 8888
rect 23716 8848 23722 8860
rect 24213 8857 24225 8860
rect 24259 8857 24271 8891
rect 24826 8888 24854 8928
rect 24826 8860 25544 8888
rect 24213 8851 24271 8857
rect 19886 8820 19892 8832
rect 19306 8792 19892 8820
rect 19886 8780 19892 8792
rect 19944 8780 19950 8832
rect 22278 8780 22284 8832
rect 22336 8820 22342 8832
rect 23937 8823 23995 8829
rect 23937 8820 23949 8823
rect 22336 8792 23949 8820
rect 22336 8780 22342 8792
rect 23937 8789 23949 8792
rect 23983 8789 23995 8823
rect 23937 8783 23995 8789
rect 24118 8780 24124 8832
rect 24176 8820 24182 8832
rect 25056 8829 25084 8860
rect 24305 8823 24363 8829
rect 24305 8820 24317 8823
rect 24176 8792 24317 8820
rect 24176 8780 24182 8792
rect 24305 8789 24317 8792
rect 24351 8789 24363 8823
rect 24305 8783 24363 8789
rect 24397 8823 24455 8829
rect 24397 8789 24409 8823
rect 24443 8820 24455 8823
rect 24857 8823 24915 8829
rect 24857 8820 24869 8823
rect 24443 8792 24869 8820
rect 24443 8789 24455 8792
rect 24397 8783 24455 8789
rect 24857 8789 24869 8792
rect 24903 8789 24915 8823
rect 24857 8783 24915 8789
rect 25041 8823 25099 8829
rect 25041 8789 25053 8823
rect 25087 8789 25099 8823
rect 25041 8783 25099 8789
rect 25314 8780 25320 8832
rect 25372 8780 25378 8832
rect 25516 8829 25544 8860
rect 25501 8823 25559 8829
rect 25501 8789 25513 8823
rect 25547 8789 25559 8823
rect 25501 8783 25559 8789
rect 28442 8780 28448 8832
rect 28500 8780 28506 8832
rect 28718 8780 28724 8832
rect 28776 8780 28782 8832
rect 29012 8829 29040 9002
rect 29086 8984 29092 9036
rect 29144 8984 29150 9036
rect 29178 8984 29184 9036
rect 29236 9024 29242 9036
rect 29564 9033 29592 9064
rect 29365 9027 29423 9033
rect 29365 9024 29377 9027
rect 29236 8996 29377 9024
rect 29236 8984 29242 8996
rect 29365 8993 29377 8996
rect 29411 8993 29423 9027
rect 29365 8987 29423 8993
rect 29549 9027 29607 9033
rect 29549 8993 29561 9027
rect 29595 8993 29607 9027
rect 29805 9027 29863 9033
rect 29805 9024 29817 9027
rect 29549 8987 29607 8993
rect 29656 8996 29817 9024
rect 29380 8956 29408 8987
rect 29656 8956 29684 8996
rect 29805 8993 29817 8996
rect 29851 8993 29863 9027
rect 29805 8987 29863 8993
rect 29380 8928 29684 8956
rect 28997 8823 29055 8829
rect 28997 8789 29009 8823
rect 29043 8820 29055 8823
rect 29178 8820 29184 8832
rect 29043 8792 29184 8820
rect 29043 8789 29055 8792
rect 28997 8783 29055 8789
rect 29178 8780 29184 8792
rect 29236 8820 29242 8832
rect 29273 8823 29331 8829
rect 29273 8820 29285 8823
rect 29236 8792 29285 8820
rect 29236 8780 29242 8792
rect 29273 8789 29285 8792
rect 29319 8789 29331 8823
rect 29273 8783 29331 8789
rect 552 8730 31372 8752
rect 552 8678 4250 8730
rect 4302 8678 4314 8730
rect 4366 8678 4378 8730
rect 4430 8678 4442 8730
rect 4494 8678 4506 8730
rect 4558 8678 11955 8730
rect 12007 8678 12019 8730
rect 12071 8678 12083 8730
rect 12135 8678 12147 8730
rect 12199 8678 12211 8730
rect 12263 8678 19660 8730
rect 19712 8678 19724 8730
rect 19776 8678 19788 8730
rect 19840 8678 19852 8730
rect 19904 8678 19916 8730
rect 19968 8678 27365 8730
rect 27417 8678 27429 8730
rect 27481 8678 27493 8730
rect 27545 8678 27557 8730
rect 27609 8678 27621 8730
rect 27673 8678 31372 8730
rect 552 8656 31372 8678
rect 1578 8576 1584 8628
rect 1636 8616 1642 8628
rect 1673 8619 1731 8625
rect 1673 8616 1685 8619
rect 1636 8588 1685 8616
rect 1636 8576 1642 8588
rect 1673 8585 1685 8588
rect 1719 8585 1731 8619
rect 1673 8579 1731 8585
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 2406 8616 2412 8628
rect 2179 8588 2412 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 1452 8452 1624 8480
rect 1452 8440 1458 8452
rect 1596 8421 1624 8452
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8381 1639 8415
rect 1688 8412 1716 8579
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 2648 8588 2697 8616
rect 2648 8576 2654 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 5776 8588 5825 8616
rect 5776 8576 5782 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 5813 8579 5871 8585
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7101 8619 7159 8625
rect 7101 8616 7113 8619
rect 7064 8588 7113 8616
rect 7064 8576 7070 8588
rect 7101 8585 7113 8588
rect 7147 8585 7159 8619
rect 12529 8619 12587 8625
rect 7101 8579 7159 8585
rect 9784 8588 11468 8616
rect 2608 8480 2636 8576
rect 7024 8480 7052 8576
rect 9784 8557 9812 8588
rect 9769 8551 9827 8557
rect 9769 8517 9781 8551
rect 9815 8517 9827 8551
rect 9769 8511 9827 8517
rect 7834 8480 7840 8492
rect 2516 8452 2636 8480
rect 6932 8452 7604 8480
rect 2516 8421 2544 8452
rect 2041 8415 2099 8421
rect 2041 8412 2053 8415
rect 1688 8384 2053 8412
rect 1581 8375 1639 8381
rect 2041 8381 2053 8384
rect 2087 8381 2099 8415
rect 2041 8375 2099 8381
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8381 2651 8415
rect 2593 8375 2651 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 1596 8344 1624 8375
rect 2608 8344 2636 8375
rect 1596 8316 2636 8344
rect 3694 8236 3700 8288
rect 3752 8276 3758 8288
rect 4154 8276 4160 8288
rect 3752 8248 4160 8276
rect 3752 8236 3758 8248
rect 4154 8236 4160 8248
rect 4212 8276 4218 8288
rect 4448 8276 4476 8375
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 6932 8421 6960 8452
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 6420 8384 6561 8412
rect 6420 8372 6426 8384
rect 6549 8381 6561 8384
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8381 7067 8415
rect 7009 8375 7067 8381
rect 4700 8347 4758 8353
rect 4700 8313 4712 8347
rect 4746 8344 4758 8347
rect 5718 8344 5724 8356
rect 4746 8316 5724 8344
rect 4746 8313 4758 8316
rect 4700 8307 4758 8313
rect 5718 8304 5724 8316
rect 5776 8344 5782 8356
rect 6273 8347 6331 8353
rect 6273 8344 6285 8347
rect 5776 8316 6285 8344
rect 5776 8304 5782 8316
rect 6273 8313 6285 8316
rect 6319 8313 6331 8347
rect 6656 8344 6684 8375
rect 7024 8344 7052 8375
rect 7466 8372 7472 8424
rect 7524 8372 7530 8424
rect 7576 8421 7604 8452
rect 7668 8452 7840 8480
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8381 7619 8415
rect 7561 8375 7619 8381
rect 7668 8344 7696 8452
rect 7834 8440 7840 8452
rect 7892 8480 7898 8492
rect 7892 8452 8524 8480
rect 7892 8440 7898 8452
rect 8386 8412 8392 8424
rect 6656 8316 7696 8344
rect 7852 8384 8392 8412
rect 6273 8307 6331 8313
rect 4212 8248 4476 8276
rect 6288 8276 6316 8307
rect 7852 8288 7880 8384
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8496 8412 8524 8452
rect 8645 8415 8703 8421
rect 8645 8412 8657 8415
rect 8496 8384 8657 8412
rect 8645 8381 8657 8384
rect 8691 8381 8703 8415
rect 8645 8375 8703 8381
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8412 10471 8415
rect 10962 8412 10968 8424
rect 10459 8384 10968 8412
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 10226 8304 10232 8356
rect 10284 8344 10290 8356
rect 10658 8347 10716 8353
rect 10658 8344 10670 8347
rect 10284 8316 10670 8344
rect 10284 8304 10290 8316
rect 10658 8313 10670 8316
rect 10704 8313 10716 8347
rect 11440 8344 11468 8588
rect 12529 8585 12541 8619
rect 12575 8616 12587 8619
rect 12894 8616 12900 8628
rect 12575 8588 12900 8616
rect 12575 8585 12587 8588
rect 12529 8579 12587 8585
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 12986 8576 12992 8628
rect 13044 8576 13050 8628
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 13320 8588 14289 8616
rect 13320 8576 13326 8588
rect 14277 8585 14289 8588
rect 14323 8585 14335 8619
rect 14277 8579 14335 8585
rect 14550 8576 14556 8628
rect 14608 8576 14614 8628
rect 15010 8576 15016 8628
rect 15068 8616 15074 8628
rect 15197 8619 15255 8625
rect 15197 8616 15209 8619
rect 15068 8588 15209 8616
rect 15068 8576 15074 8588
rect 15197 8585 15209 8588
rect 15243 8585 15255 8619
rect 15197 8579 15255 8585
rect 15838 8576 15844 8628
rect 15896 8616 15902 8628
rect 16390 8616 16396 8628
rect 15896 8588 16396 8616
rect 15896 8576 15902 8588
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 16758 8576 16764 8628
rect 16816 8576 16822 8628
rect 17037 8619 17095 8625
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 17126 8616 17132 8628
rect 17083 8588 17132 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 17221 8619 17279 8625
rect 17221 8585 17233 8619
rect 17267 8585 17279 8619
rect 17221 8579 17279 8585
rect 17681 8619 17739 8625
rect 17681 8585 17693 8619
rect 17727 8616 17739 8619
rect 17770 8616 17776 8628
rect 17727 8588 17776 8616
rect 17727 8585 17739 8588
rect 17681 8579 17739 8585
rect 11793 8551 11851 8557
rect 11793 8517 11805 8551
rect 11839 8517 11851 8551
rect 11793 8511 11851 8517
rect 11808 8480 11836 8511
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 12621 8551 12679 8557
rect 12621 8548 12633 8551
rect 11940 8520 12633 8548
rect 11940 8508 11946 8520
rect 12621 8517 12633 8520
rect 12667 8517 12679 8551
rect 12621 8511 12679 8517
rect 13354 8508 13360 8560
rect 13412 8548 13418 8560
rect 13909 8551 13967 8557
rect 13909 8548 13921 8551
rect 13412 8520 13921 8548
rect 13412 8508 13418 8520
rect 13909 8517 13921 8520
rect 13955 8517 13967 8551
rect 13909 8511 13967 8517
rect 14001 8551 14059 8557
rect 14001 8517 14013 8551
rect 14047 8548 14059 8551
rect 14182 8548 14188 8560
rect 14047 8520 14188 8548
rect 14047 8517 14059 8520
rect 14001 8511 14059 8517
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 14737 8551 14795 8557
rect 14737 8517 14749 8551
rect 14783 8548 14795 8551
rect 15289 8551 15347 8557
rect 15289 8548 15301 8551
rect 14783 8520 15301 8548
rect 14783 8517 14795 8520
rect 14737 8511 14795 8517
rect 15289 8517 15301 8520
rect 15335 8517 15347 8551
rect 15289 8511 15347 8517
rect 16114 8508 16120 8560
rect 16172 8548 16178 8560
rect 16776 8548 16804 8576
rect 16172 8520 16804 8548
rect 16172 8508 16178 8520
rect 14921 8483 14979 8489
rect 11808 8452 12480 8480
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12342 8412 12348 8424
rect 12299 8384 12348 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 12452 8421 12480 8452
rect 12544 8452 13584 8480
rect 12544 8424 12572 8452
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 12526 8372 12532 8424
rect 12584 8372 12590 8424
rect 12710 8372 12716 8424
rect 12768 8372 12774 8424
rect 13354 8372 13360 8424
rect 13412 8412 13418 8424
rect 13556 8421 13584 8452
rect 14921 8449 14933 8483
rect 14967 8480 14979 8483
rect 17236 8480 17264 8579
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 19705 8619 19763 8625
rect 19705 8616 19717 8619
rect 18288 8588 19717 8616
rect 18288 8576 18294 8588
rect 19705 8585 19717 8588
rect 19751 8585 19763 8619
rect 19705 8579 19763 8585
rect 19978 8576 19984 8628
rect 20036 8576 20042 8628
rect 21082 8576 21088 8628
rect 21140 8616 21146 8628
rect 21726 8616 21732 8628
rect 21140 8588 21732 8616
rect 21140 8576 21146 8588
rect 21726 8576 21732 8588
rect 21784 8576 21790 8628
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 23474 8616 23480 8628
rect 22060 8588 23480 8616
rect 22060 8576 22066 8588
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 23658 8576 23664 8628
rect 23716 8576 23722 8628
rect 24305 8619 24363 8625
rect 24305 8585 24317 8619
rect 24351 8616 24363 8619
rect 25314 8616 25320 8628
rect 24351 8588 25320 8616
rect 24351 8585 24363 8588
rect 24305 8579 24363 8585
rect 25314 8576 25320 8588
rect 25372 8576 25378 8628
rect 26510 8576 26516 8628
rect 26568 8576 26574 8628
rect 28442 8576 28448 8628
rect 28500 8616 28506 8628
rect 29365 8619 29423 8625
rect 29365 8616 29377 8619
rect 28500 8588 29377 8616
rect 28500 8576 28506 8588
rect 29365 8585 29377 8588
rect 29411 8616 29423 8619
rect 29730 8616 29736 8628
rect 29411 8588 29736 8616
rect 29411 8585 29423 8588
rect 29365 8579 29423 8585
rect 29730 8576 29736 8588
rect 29788 8616 29794 8628
rect 29788 8588 30144 8616
rect 29788 8576 29794 8588
rect 19337 8551 19395 8557
rect 19337 8517 19349 8551
rect 19383 8548 19395 8551
rect 19797 8551 19855 8557
rect 19797 8548 19809 8551
rect 19383 8520 19809 8548
rect 19383 8517 19395 8520
rect 19337 8511 19395 8517
rect 19797 8517 19809 8520
rect 19843 8517 19855 8551
rect 19797 8511 19855 8517
rect 22646 8508 22652 8560
rect 22704 8548 22710 8560
rect 22704 8520 24256 8548
rect 22704 8508 22710 8520
rect 14967 8452 17264 8480
rect 14967 8449 14979 8452
rect 14921 8443 14979 8449
rect 17586 8440 17592 8492
rect 17644 8480 17650 8492
rect 19518 8480 19524 8492
rect 17644 8452 19524 8480
rect 17644 8440 17650 8452
rect 19518 8440 19524 8452
rect 19576 8440 19582 8492
rect 19610 8440 19616 8492
rect 19668 8480 19674 8492
rect 19886 8480 19892 8492
rect 19668 8452 19892 8480
rect 19668 8440 19674 8452
rect 19886 8440 19892 8452
rect 19944 8480 19950 8492
rect 20162 8480 20168 8492
rect 19944 8452 20168 8480
rect 19944 8440 19950 8452
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 24228 8489 24256 8520
rect 30006 8508 30012 8560
rect 30064 8508 30070 8560
rect 24213 8483 24271 8489
rect 22296 8452 23888 8480
rect 13541 8415 13599 8421
rect 13541 8412 13553 8415
rect 13412 8384 13553 8412
rect 13412 8372 13418 8384
rect 13541 8381 13553 8384
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 13814 8372 13820 8424
rect 13872 8372 13878 8424
rect 14182 8372 14188 8424
rect 14240 8412 14246 8424
rect 14550 8412 14556 8424
rect 14240 8384 14556 8412
rect 14240 8372 14246 8384
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 15378 8372 15384 8424
rect 15436 8372 15442 8424
rect 15470 8372 15476 8424
rect 15528 8372 15534 8424
rect 15660 8415 15718 8421
rect 15660 8381 15672 8415
rect 15706 8412 15718 8415
rect 15838 8412 15844 8424
rect 15706 8384 15844 8412
rect 15706 8381 15718 8384
rect 15660 8375 15718 8381
rect 15838 8372 15844 8384
rect 15896 8372 15902 8424
rect 16025 8415 16083 8421
rect 16025 8381 16037 8415
rect 16071 8381 16083 8415
rect 16025 8375 16083 8381
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8381 16267 8415
rect 16209 8375 16267 8381
rect 14369 8347 14427 8353
rect 14369 8344 14381 8347
rect 11440 8316 14381 8344
rect 10658 8307 10716 8313
rect 14369 8313 14381 8316
rect 14415 8313 14427 8347
rect 16040 8344 16068 8375
rect 14369 8307 14427 8313
rect 15672 8316 16068 8344
rect 16224 8344 16252 8375
rect 16666 8372 16672 8424
rect 16724 8372 16730 8424
rect 16853 8415 16911 8421
rect 16853 8381 16865 8415
rect 16899 8412 16911 8415
rect 16942 8412 16948 8424
rect 16899 8384 16948 8412
rect 16899 8381 16911 8384
rect 16853 8375 16911 8381
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 17310 8412 17316 8424
rect 17052 8384 17316 8412
rect 16390 8344 16396 8356
rect 16224 8316 16396 8344
rect 15672 8288 15700 8316
rect 16390 8304 16396 8316
rect 16448 8344 16454 8356
rect 17052 8344 17080 8384
rect 17310 8372 17316 8384
rect 17368 8372 17374 8424
rect 17402 8372 17408 8424
rect 17460 8372 17466 8424
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8412 17555 8415
rect 17954 8412 17960 8424
rect 17543 8384 17960 8412
rect 17543 8381 17555 8384
rect 17497 8375 17555 8381
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 18969 8415 19027 8421
rect 18969 8381 18981 8415
rect 19015 8412 19027 8415
rect 19058 8412 19064 8424
rect 19015 8384 19064 8412
rect 19015 8381 19027 8384
rect 18969 8375 19027 8381
rect 19058 8372 19064 8384
rect 19116 8372 19122 8424
rect 19150 8372 19156 8424
rect 19208 8372 19214 8424
rect 19242 8372 19248 8424
rect 19300 8372 19306 8424
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8412 19487 8415
rect 19794 8412 19800 8424
rect 19475 8384 19800 8412
rect 19475 8381 19487 8384
rect 19429 8375 19487 8381
rect 19794 8372 19800 8384
rect 19852 8372 19858 8424
rect 22296 8412 22324 8452
rect 20104 8384 22324 8412
rect 22373 8415 22431 8421
rect 16448 8316 17080 8344
rect 17221 8347 17279 8353
rect 16448 8304 16454 8316
rect 17221 8313 17233 8347
rect 17267 8344 17279 8347
rect 20104 8344 20132 8384
rect 22373 8381 22385 8415
rect 22419 8412 22431 8415
rect 22462 8412 22468 8424
rect 22419 8384 22468 8412
rect 22419 8381 22431 8384
rect 22373 8375 22431 8381
rect 22462 8372 22468 8384
rect 22520 8412 22526 8424
rect 22922 8412 22928 8424
rect 22520 8384 22928 8412
rect 22520 8372 22526 8384
rect 22922 8372 22928 8384
rect 22980 8372 22986 8424
rect 23106 8372 23112 8424
rect 23164 8372 23170 8424
rect 23860 8421 23888 8452
rect 24213 8449 24225 8483
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 27890 8440 27896 8492
rect 27948 8440 27954 8492
rect 28718 8440 28724 8492
rect 28776 8480 28782 8492
rect 30024 8480 30052 8508
rect 28776 8452 29316 8480
rect 28776 8440 28782 8452
rect 23845 8415 23903 8421
rect 23845 8381 23857 8415
rect 23891 8381 23903 8415
rect 23845 8375 23903 8381
rect 24118 8372 24124 8424
rect 24176 8372 24182 8424
rect 24394 8372 24400 8424
rect 24452 8412 24458 8424
rect 24581 8415 24639 8421
rect 24581 8412 24593 8415
rect 24452 8384 24593 8412
rect 24452 8372 24458 8384
rect 24581 8381 24593 8384
rect 24627 8381 24639 8415
rect 24581 8375 24639 8381
rect 26237 8415 26295 8421
rect 26237 8381 26249 8415
rect 26283 8412 26295 8415
rect 27908 8412 27936 8440
rect 28813 8415 28871 8421
rect 28813 8412 28825 8415
rect 26283 8384 27936 8412
rect 28644 8384 28825 8412
rect 26283 8381 26295 8384
rect 26237 8375 26295 8381
rect 17267 8316 20132 8344
rect 20165 8347 20223 8353
rect 17267 8313 17279 8316
rect 17221 8307 17279 8313
rect 20165 8313 20177 8347
rect 20211 8344 20223 8347
rect 20211 8316 21036 8344
rect 20211 8313 20223 8316
rect 20165 8307 20223 8313
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6288 8248 6837 8276
rect 4212 8236 4218 8248
rect 6825 8245 6837 8248
rect 6871 8245 6883 8279
rect 6825 8239 6883 8245
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 7653 8279 7711 8285
rect 7653 8276 7665 8279
rect 7432 8248 7665 8276
rect 7432 8236 7438 8248
rect 7653 8245 7665 8248
rect 7699 8245 7711 8279
rect 7653 8239 7711 8245
rect 7834 8236 7840 8288
rect 7892 8236 7898 8288
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 13633 8279 13691 8285
rect 13633 8276 13645 8279
rect 13044 8248 13645 8276
rect 13044 8236 13050 8248
rect 13633 8245 13645 8248
rect 13679 8245 13691 8279
rect 13633 8239 13691 8245
rect 14550 8236 14556 8288
rect 14608 8285 14614 8288
rect 14608 8279 14627 8285
rect 14615 8245 14627 8279
rect 14608 8239 14627 8245
rect 14608 8236 14614 8239
rect 15654 8236 15660 8288
rect 15712 8236 15718 8288
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 16758 8276 16764 8288
rect 16080 8248 16764 8276
rect 16080 8236 16086 8248
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 17034 8236 17040 8288
rect 17092 8276 17098 8288
rect 18966 8276 18972 8288
rect 17092 8248 18972 8276
rect 17092 8236 17098 8248
rect 18966 8236 18972 8248
rect 19024 8276 19030 8288
rect 21008 8285 21036 8316
rect 22094 8304 22100 8356
rect 22152 8353 22158 8356
rect 22152 8344 22164 8353
rect 23124 8344 23152 8372
rect 23293 8347 23351 8353
rect 22152 8316 22197 8344
rect 23124 8316 23244 8344
rect 22152 8307 22164 8316
rect 22152 8304 22158 8307
rect 19955 8279 20013 8285
rect 19955 8276 19967 8279
rect 19024 8248 19967 8276
rect 19024 8236 19030 8248
rect 19955 8245 19967 8248
rect 20001 8245 20013 8279
rect 19955 8239 20013 8245
rect 20993 8279 21051 8285
rect 20993 8245 21005 8279
rect 21039 8245 21051 8279
rect 23216 8276 23244 8316
rect 23293 8313 23305 8347
rect 23339 8344 23351 8347
rect 23339 8316 24900 8344
rect 23339 8313 23351 8316
rect 23293 8307 23351 8313
rect 23493 8279 23551 8285
rect 23493 8276 23505 8279
rect 23216 8248 23505 8276
rect 20993 8239 21051 8245
rect 23493 8245 23505 8248
rect 23539 8245 23551 8279
rect 23493 8239 23551 8245
rect 24486 8236 24492 8288
rect 24544 8236 24550 8288
rect 24872 8285 24900 8316
rect 25774 8304 25780 8356
rect 25832 8344 25838 8356
rect 25970 8347 26028 8353
rect 25970 8344 25982 8347
rect 25832 8316 25982 8344
rect 25832 8304 25838 8316
rect 25970 8313 25982 8316
rect 26016 8313 26028 8347
rect 25970 8307 26028 8313
rect 27648 8347 27706 8353
rect 27648 8313 27660 8347
rect 27694 8344 27706 8347
rect 28534 8344 28540 8356
rect 27694 8316 28540 8344
rect 27694 8313 27706 8316
rect 27648 8307 27706 8313
rect 28534 8304 28540 8316
rect 28592 8304 28598 8356
rect 24857 8279 24915 8285
rect 24857 8245 24869 8279
rect 24903 8245 24915 8279
rect 28644 8276 28672 8384
rect 28813 8381 28825 8384
rect 28859 8381 28871 8415
rect 28813 8375 28871 8381
rect 29178 8372 29184 8424
rect 29236 8372 29242 8424
rect 29288 8412 29316 8452
rect 29656 8452 30052 8480
rect 29457 8415 29515 8421
rect 29457 8412 29469 8415
rect 29288 8384 29469 8412
rect 29457 8381 29469 8384
rect 29503 8412 29515 8415
rect 29656 8412 29684 8452
rect 29503 8384 29684 8412
rect 29503 8381 29515 8384
rect 29457 8375 29515 8381
rect 29730 8372 29736 8424
rect 29788 8372 29794 8424
rect 30024 8421 30052 8452
rect 30116 8421 30144 8588
rect 30009 8415 30067 8421
rect 30009 8381 30021 8415
rect 30055 8381 30067 8415
rect 30009 8375 30067 8381
rect 30101 8415 30159 8421
rect 30101 8381 30113 8415
rect 30147 8381 30159 8415
rect 30101 8375 30159 8381
rect 30466 8372 30472 8424
rect 30524 8412 30530 8424
rect 30561 8415 30619 8421
rect 30561 8412 30573 8415
rect 30524 8384 30573 8412
rect 30524 8372 30530 8384
rect 30561 8381 30573 8384
rect 30607 8381 30619 8415
rect 30561 8375 30619 8381
rect 30653 8415 30711 8421
rect 30653 8381 30665 8415
rect 30699 8381 30711 8415
rect 30653 8375 30711 8381
rect 28721 8347 28779 8353
rect 28721 8313 28733 8347
rect 28767 8344 28779 8347
rect 28994 8344 29000 8356
rect 28767 8316 29000 8344
rect 28767 8313 28779 8316
rect 28721 8307 28779 8313
rect 28994 8304 29000 8316
rect 29052 8344 29058 8356
rect 29917 8347 29975 8353
rect 29917 8344 29929 8347
rect 29052 8316 29929 8344
rect 29052 8304 29058 8316
rect 29917 8313 29929 8316
rect 29963 8313 29975 8347
rect 30668 8344 30696 8375
rect 29917 8307 29975 8313
rect 30208 8316 30696 8344
rect 30208 8288 30236 8316
rect 29089 8279 29147 8285
rect 29089 8276 29101 8279
rect 28644 8248 29101 8276
rect 24857 8239 24915 8245
rect 29089 8245 29101 8248
rect 29135 8276 29147 8279
rect 29641 8279 29699 8285
rect 29641 8276 29653 8279
rect 29135 8248 29653 8276
rect 29135 8245 29147 8248
rect 29089 8239 29147 8245
rect 29641 8245 29653 8248
rect 29687 8276 29699 8279
rect 29730 8276 29736 8288
rect 29687 8248 29736 8276
rect 29687 8245 29699 8248
rect 29641 8239 29699 8245
rect 29730 8236 29736 8248
rect 29788 8236 29794 8288
rect 30190 8236 30196 8288
rect 30248 8236 30254 8288
rect 30374 8236 30380 8288
rect 30432 8276 30438 8288
rect 30469 8279 30527 8285
rect 30469 8276 30481 8279
rect 30432 8248 30481 8276
rect 30432 8236 30438 8248
rect 30469 8245 30481 8248
rect 30515 8245 30527 8279
rect 30469 8239 30527 8245
rect 30742 8236 30748 8288
rect 30800 8236 30806 8288
rect 552 8186 31531 8208
rect 552 8134 8102 8186
rect 8154 8134 8166 8186
rect 8218 8134 8230 8186
rect 8282 8134 8294 8186
rect 8346 8134 8358 8186
rect 8410 8134 15807 8186
rect 15859 8134 15871 8186
rect 15923 8134 15935 8186
rect 15987 8134 15999 8186
rect 16051 8134 16063 8186
rect 16115 8134 23512 8186
rect 23564 8134 23576 8186
rect 23628 8134 23640 8186
rect 23692 8134 23704 8186
rect 23756 8134 23768 8186
rect 23820 8134 31217 8186
rect 31269 8134 31281 8186
rect 31333 8134 31345 8186
rect 31397 8134 31409 8186
rect 31461 8134 31473 8186
rect 31525 8134 31531 8186
rect 552 8112 31531 8134
rect 3605 8075 3663 8081
rect 3605 8041 3617 8075
rect 3651 8072 3663 8075
rect 6181 8075 6239 8081
rect 3651 8044 6132 8072
rect 3651 8041 3663 8044
rect 3605 8035 3663 8041
rect 2240 7976 2774 8004
rect 1946 7828 1952 7880
rect 2004 7868 2010 7880
rect 2240 7877 2268 7976
rect 2498 7945 2504 7948
rect 2492 7936 2504 7945
rect 2459 7908 2504 7936
rect 2492 7899 2504 7908
rect 2498 7896 2504 7899
rect 2556 7896 2562 7948
rect 2746 7936 2774 7976
rect 3786 7964 3792 8016
rect 3844 8004 3850 8016
rect 3942 8007 4000 8013
rect 3942 8004 3954 8007
rect 3844 7976 3954 8004
rect 3844 7964 3850 7976
rect 3942 7973 3954 7976
rect 3988 7973 4000 8007
rect 3942 7967 4000 7973
rect 5718 7964 5724 8016
rect 5776 8004 5782 8016
rect 6104 8004 6132 8044
rect 6181 8041 6193 8075
rect 6227 8072 6239 8075
rect 6362 8072 6368 8084
rect 6227 8044 6368 8072
rect 6227 8041 6239 8044
rect 6181 8035 6239 8041
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 7116 8044 8800 8072
rect 7116 8004 7144 8044
rect 7374 8004 7380 8016
rect 5776 7976 5856 8004
rect 6104 7976 7144 8004
rect 7208 7976 7380 8004
rect 5776 7964 5782 7976
rect 3694 7936 3700 7948
rect 2746 7908 3700 7936
rect 3694 7896 3700 7908
rect 3752 7896 3758 7948
rect 5828 7945 5856 7976
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 5813 7939 5871 7945
rect 5675 7908 5764 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 5736 7880 5764 7908
rect 5813 7905 5825 7939
rect 5859 7936 5871 7939
rect 6086 7936 6092 7948
rect 5859 7908 6092 7936
rect 5859 7905 5871 7908
rect 5813 7899 5871 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7936 6331 7939
rect 7208 7936 7236 7976
rect 7374 7964 7380 7976
rect 7432 8004 7438 8016
rect 8082 8007 8140 8013
rect 8082 8004 8094 8007
rect 7432 7976 8094 8004
rect 7432 7964 7438 7976
rect 6319 7908 7236 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 7282 7896 7288 7948
rect 7340 7896 7346 7948
rect 7576 7945 7604 7976
rect 8082 7973 8094 7976
rect 8128 7973 8140 8007
rect 8772 8004 8800 8044
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 12986 8072 12992 8084
rect 8904 8044 12992 8072
rect 8904 8032 8910 8044
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 13173 8075 13231 8081
rect 13173 8041 13185 8075
rect 13219 8072 13231 8075
rect 13633 8075 13691 8081
rect 13219 8044 13584 8072
rect 13219 8041 13231 8044
rect 13173 8035 13231 8041
rect 8772 7976 12664 8004
rect 8082 7967 8140 7973
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 10318 7896 10324 7948
rect 10376 7936 10382 7948
rect 11221 7939 11279 7945
rect 11221 7936 11233 7939
rect 10376 7908 11233 7936
rect 10376 7896 10382 7908
rect 11221 7905 11233 7908
rect 11267 7905 11279 7939
rect 11221 7899 11279 7905
rect 12437 7939 12495 7945
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 12526 7936 12532 7948
rect 12483 7908 12532 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 12636 7945 12664 7976
rect 13262 7964 13268 8016
rect 13320 7964 13326 8016
rect 13354 7964 13360 8016
rect 13412 7964 13418 8016
rect 13446 7964 13452 8016
rect 13504 8013 13510 8016
rect 13504 8007 13523 8013
rect 13511 7973 13523 8007
rect 13556 8004 13584 8044
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13814 8072 13820 8084
rect 13679 8044 13820 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 15102 8032 15108 8084
rect 15160 8032 15166 8084
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 16117 8075 16175 8081
rect 15252 8044 16068 8072
rect 15252 8032 15258 8044
rect 15120 8004 15148 8032
rect 13556 7976 15148 8004
rect 13504 7967 13523 7973
rect 13504 7964 13510 7967
rect 15286 7964 15292 8016
rect 15344 7964 15350 8016
rect 16040 8004 16068 8044
rect 16117 8041 16129 8075
rect 16163 8072 16175 8075
rect 16390 8072 16396 8084
rect 16163 8044 16396 8072
rect 16163 8041 16175 8044
rect 16117 8035 16175 8041
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 16666 8032 16672 8084
rect 16724 8032 16730 8084
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 17034 8072 17040 8084
rect 16816 8044 17040 8072
rect 16816 8032 16822 8044
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 17678 8032 17684 8084
rect 17736 8072 17742 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17736 8044 17785 8072
rect 17736 8032 17742 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 17773 8035 17831 8041
rect 17862 8032 17868 8084
rect 17920 8072 17926 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 17920 8044 18613 8072
rect 17920 8032 17926 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 18769 8075 18827 8081
rect 18769 8041 18781 8075
rect 18815 8072 18827 8075
rect 18815 8044 18920 8072
rect 18815 8041 18827 8044
rect 18769 8035 18827 8041
rect 16040 7976 18276 8004
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7905 12679 7939
rect 13372 7936 13400 7964
rect 14001 7939 14059 7945
rect 14001 7936 14013 7939
rect 13372 7908 14013 7936
rect 12621 7899 12679 7905
rect 14001 7905 14013 7908
rect 14047 7905 14059 7939
rect 14001 7899 14059 7905
rect 14185 7939 14243 7945
rect 14185 7905 14197 7939
rect 14231 7936 14243 7939
rect 14231 7908 14320 7936
rect 15304 7935 15332 7964
rect 15473 7939 15531 7945
rect 14231 7905 14243 7908
rect 14185 7899 14243 7905
rect 14292 7880 14320 7908
rect 15289 7929 15347 7935
rect 15289 7895 15301 7929
rect 15335 7895 15347 7929
rect 15473 7905 15485 7939
rect 15519 7936 15531 7939
rect 15562 7936 15568 7948
rect 15519 7908 15568 7936
rect 15519 7905 15531 7908
rect 15473 7899 15531 7905
rect 15562 7896 15568 7908
rect 15620 7936 15626 7948
rect 16390 7936 16396 7948
rect 15620 7908 16396 7936
rect 15620 7896 15626 7908
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 16516 7908 16865 7936
rect 15289 7889 15347 7895
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 2004 7840 2237 7868
rect 2004 7828 2010 7840
rect 2225 7837 2237 7840
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 5718 7828 5724 7880
rect 5776 7828 5782 7880
rect 6546 7828 6552 7880
rect 6604 7868 6610 7880
rect 7834 7868 7840 7880
rect 6604 7840 7840 7868
rect 6604 7828 6610 7840
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 8846 7828 8852 7880
rect 8904 7828 8910 7880
rect 10962 7828 10968 7880
rect 11020 7828 11026 7880
rect 12360 7840 14228 7868
rect 5077 7803 5135 7809
rect 5077 7769 5089 7803
rect 5123 7800 5135 7803
rect 5123 7772 7604 7800
rect 5123 7769 5135 7772
rect 5077 7763 5135 7769
rect 5537 7735 5595 7741
rect 5537 7701 5549 7735
rect 5583 7732 5595 7735
rect 5626 7732 5632 7744
rect 5583 7704 5632 7732
rect 5583 7701 5595 7704
rect 5537 7695 5595 7701
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 5718 7692 5724 7744
rect 5776 7732 5782 7744
rect 5905 7735 5963 7741
rect 5905 7732 5917 7735
rect 5776 7704 5917 7732
rect 5776 7692 5782 7704
rect 5905 7701 5917 7704
rect 5951 7732 5963 7735
rect 6270 7732 6276 7744
rect 5951 7704 6276 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 6270 7692 6276 7704
rect 6328 7732 6334 7744
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 6328 7704 7481 7732
rect 6328 7692 6334 7704
rect 7469 7701 7481 7704
rect 7515 7701 7527 7735
rect 7576 7732 7604 7772
rect 8864 7732 8892 7828
rect 12360 7809 12388 7840
rect 12345 7803 12403 7809
rect 12345 7769 12357 7803
rect 12391 7769 12403 7803
rect 14090 7800 14096 7812
rect 12345 7763 12403 7769
rect 13004 7772 14096 7800
rect 13004 7744 13032 7772
rect 7576 7704 8892 7732
rect 9217 7735 9275 7741
rect 7469 7695 7527 7701
rect 9217 7701 9229 7735
rect 9263 7732 9275 7735
rect 11238 7732 11244 7744
rect 9263 7704 11244 7732
rect 9263 7701 9275 7704
rect 9217 7695 9275 7701
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 12618 7692 12624 7744
rect 12676 7732 12682 7744
rect 12713 7735 12771 7741
rect 12713 7732 12725 7735
rect 12676 7704 12725 7732
rect 12676 7692 12682 7704
rect 12713 7701 12725 7704
rect 12759 7701 12771 7735
rect 12713 7695 12771 7701
rect 12802 7692 12808 7744
rect 12860 7692 12866 7744
rect 12894 7692 12900 7744
rect 12952 7692 12958 7744
rect 12986 7692 12992 7744
rect 13044 7692 13050 7744
rect 13464 7741 13492 7772
rect 14090 7760 14096 7772
rect 14148 7760 14154 7812
rect 14200 7800 14228 7840
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7868 14427 7871
rect 14734 7868 14740 7880
rect 14415 7840 14740 7868
rect 14415 7837 14427 7840
rect 14369 7831 14427 7837
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 16301 7803 16359 7809
rect 14200 7772 15884 7800
rect 13449 7735 13507 7741
rect 13449 7701 13461 7735
rect 13495 7701 13507 7735
rect 13449 7695 13507 7701
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 15105 7735 15163 7741
rect 15105 7732 15117 7735
rect 13872 7704 15117 7732
rect 13872 7692 13878 7704
rect 15105 7701 15117 7704
rect 15151 7701 15163 7735
rect 15856 7732 15884 7772
rect 16301 7769 16313 7803
rect 16347 7800 16359 7803
rect 16516 7800 16544 7908
rect 16853 7905 16865 7908
rect 16899 7936 16911 7939
rect 16899 7908 17356 7936
rect 16899 7905 16911 7908
rect 16853 7899 16911 7905
rect 17328 7877 17356 7908
rect 18138 7896 18144 7948
rect 18196 7896 18202 7948
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 16623 7840 17049 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 17037 7837 17049 7840
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 17313 7871 17371 7877
rect 17313 7837 17325 7871
rect 17359 7868 17371 7871
rect 17678 7868 17684 7880
rect 17359 7840 17684 7868
rect 17359 7837 17371 7840
rect 17313 7831 17371 7837
rect 16347 7772 16544 7800
rect 17052 7800 17080 7831
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 17218 7800 17224 7812
rect 17052 7772 17224 7800
rect 16347 7769 16359 7772
rect 16301 7763 16359 7769
rect 17218 7760 17224 7772
rect 17276 7800 17282 7812
rect 17589 7803 17647 7809
rect 17589 7800 17601 7803
rect 17276 7772 17601 7800
rect 17276 7760 17282 7772
rect 17589 7769 17601 7772
rect 17635 7769 17647 7803
rect 18248 7800 18276 7976
rect 18506 7896 18512 7948
rect 18564 7936 18570 7948
rect 18782 7936 18788 7948
rect 18564 7908 18788 7936
rect 18564 7896 18570 7908
rect 18782 7896 18788 7908
rect 18840 7896 18846 7948
rect 18892 7936 18920 8044
rect 19242 8032 19248 8084
rect 19300 8072 19306 8084
rect 19337 8075 19395 8081
rect 19337 8072 19349 8075
rect 19300 8044 19349 8072
rect 19300 8032 19306 8044
rect 19337 8041 19349 8044
rect 19383 8041 19395 8075
rect 19337 8035 19395 8041
rect 19505 8075 19563 8081
rect 19505 8041 19517 8075
rect 19551 8072 19563 8075
rect 19610 8072 19616 8084
rect 19551 8044 19616 8072
rect 19551 8041 19563 8044
rect 19505 8035 19563 8041
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 19794 8032 19800 8084
rect 19852 8072 19858 8084
rect 20257 8075 20315 8081
rect 20257 8072 20269 8075
rect 19852 8044 20269 8072
rect 19852 8032 19858 8044
rect 20257 8041 20269 8044
rect 20303 8041 20315 8075
rect 20257 8035 20315 8041
rect 20425 8075 20483 8081
rect 20425 8041 20437 8075
rect 20471 8072 20483 8075
rect 20530 8072 20536 8084
rect 20471 8044 20536 8072
rect 20471 8041 20483 8044
rect 20425 8035 20483 8041
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 21634 8072 21640 8084
rect 21560 8044 21640 8072
rect 18966 7964 18972 8016
rect 19024 7964 19030 8016
rect 19702 7964 19708 8016
rect 19760 7964 19766 8016
rect 20165 8007 20223 8013
rect 19935 7973 19993 7979
rect 19935 7939 19947 7973
rect 19981 7939 19993 7973
rect 20165 7973 20177 8007
rect 20211 8004 20223 8007
rect 20625 8007 20683 8013
rect 20211 7976 20576 8004
rect 20211 7973 20223 7976
rect 20165 7967 20223 7973
rect 19935 7936 19993 7939
rect 18892 7933 19993 7936
rect 18892 7908 19992 7933
rect 19260 7880 19288 7908
rect 19242 7828 19248 7880
rect 19300 7828 19306 7880
rect 19978 7828 19984 7880
rect 20036 7828 20042 7880
rect 19797 7803 19855 7809
rect 19797 7800 19809 7803
rect 18248 7772 19809 7800
rect 17589 7763 17647 7769
rect 19797 7769 19809 7772
rect 19843 7769 19855 7803
rect 19797 7763 19855 7769
rect 18690 7732 18696 7744
rect 15856 7704 18696 7732
rect 15105 7695 15163 7701
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 18782 7692 18788 7744
rect 18840 7732 18846 7744
rect 19996 7741 20024 7828
rect 20548 7800 20576 7976
rect 20625 7973 20637 8007
rect 20671 7973 20683 8007
rect 20625 7967 20683 7973
rect 20640 7868 20668 7967
rect 21560 7945 21588 8044
rect 21634 8032 21640 8044
rect 21692 8032 21698 8084
rect 21726 8032 21732 8084
rect 21784 8072 21790 8084
rect 22005 8075 22063 8081
rect 22005 8072 22017 8075
rect 21784 8044 22017 8072
rect 21784 8032 21790 8044
rect 22005 8041 22017 8044
rect 22051 8072 22063 8075
rect 22094 8072 22100 8084
rect 22051 8044 22100 8072
rect 22051 8041 22063 8044
rect 22005 8035 22063 8041
rect 22094 8032 22100 8044
rect 22152 8032 22158 8084
rect 22281 8075 22339 8081
rect 22281 8041 22293 8075
rect 22327 8072 22339 8075
rect 22554 8072 22560 8084
rect 22327 8044 22560 8072
rect 22327 8041 22339 8044
rect 22281 8035 22339 8041
rect 22554 8032 22560 8044
rect 22612 8032 22618 8084
rect 24397 8075 24455 8081
rect 24397 8041 24409 8075
rect 24443 8072 24455 8075
rect 24486 8072 24492 8084
rect 24443 8044 24492 8072
rect 24443 8041 24455 8044
rect 24397 8035 24455 8041
rect 24486 8032 24492 8044
rect 24544 8032 24550 8084
rect 27890 8032 27896 8084
rect 27948 8032 27954 8084
rect 28534 8032 28540 8084
rect 28592 8072 28598 8084
rect 30282 8072 30288 8084
rect 28592 8044 30288 8072
rect 28592 8032 28598 8044
rect 30282 8032 30288 8044
rect 30340 8032 30346 8084
rect 30926 8032 30932 8084
rect 30984 8032 30990 8084
rect 21545 7939 21603 7945
rect 21545 7905 21557 7939
rect 21591 7905 21603 7939
rect 21545 7899 21603 7905
rect 21637 7939 21695 7945
rect 21637 7905 21649 7939
rect 21683 7934 21695 7939
rect 21744 7934 21772 8032
rect 21818 7964 21824 8016
rect 21876 8004 21882 8016
rect 21876 7976 22508 8004
rect 21876 7964 21882 7976
rect 21683 7906 21772 7934
rect 22097 7939 22155 7945
rect 21683 7905 21695 7906
rect 21637 7899 21695 7905
rect 22097 7905 22109 7939
rect 22143 7936 22155 7939
rect 22186 7936 22192 7948
rect 22143 7908 22192 7936
rect 22143 7905 22155 7908
rect 22097 7899 22155 7905
rect 22186 7896 22192 7908
rect 22244 7936 22250 7948
rect 22480 7945 22508 7976
rect 22373 7939 22431 7945
rect 22373 7936 22385 7939
rect 22244 7908 22385 7936
rect 22244 7896 22250 7908
rect 22373 7905 22385 7908
rect 22419 7905 22431 7939
rect 22373 7899 22431 7905
rect 22465 7939 22523 7945
rect 22465 7905 22477 7939
rect 22511 7905 22523 7939
rect 22465 7899 22523 7905
rect 22646 7896 22652 7948
rect 22704 7936 22710 7948
rect 23273 7939 23331 7945
rect 23273 7936 23285 7939
rect 22704 7908 23285 7936
rect 22704 7896 22710 7908
rect 23273 7905 23285 7908
rect 23319 7905 23331 7939
rect 23273 7899 23331 7905
rect 25958 7896 25964 7948
rect 26016 7936 26022 7948
rect 26237 7939 26295 7945
rect 26237 7936 26249 7939
rect 26016 7908 26249 7936
rect 26016 7896 26022 7908
rect 26237 7905 26249 7908
rect 26283 7905 26295 7939
rect 26237 7899 26295 7905
rect 27798 7896 27804 7948
rect 27856 7945 27862 7948
rect 27856 7899 27868 7945
rect 27908 7936 27936 8032
rect 28905 8007 28963 8013
rect 28905 7973 28917 8007
rect 28951 8004 28963 8007
rect 29794 8007 29852 8013
rect 29794 8004 29806 8007
rect 28951 7976 29806 8004
rect 28951 7973 28963 7976
rect 28905 7967 28963 7973
rect 29794 7973 29806 7976
rect 29840 8004 29852 8007
rect 30190 8004 30196 8016
rect 29840 7976 30196 8004
rect 29840 7973 29852 7976
rect 29794 7967 29852 7973
rect 30190 7964 30196 7976
rect 30248 8004 30254 8016
rect 30558 8004 30564 8016
rect 30248 7976 30564 8004
rect 30248 7964 30254 7976
rect 30558 7964 30564 7976
rect 30616 7964 30622 8016
rect 28077 7939 28135 7945
rect 28077 7936 28089 7939
rect 27908 7908 28089 7936
rect 28077 7905 28089 7908
rect 28123 7905 28135 7939
rect 28077 7899 28135 7905
rect 28721 7939 28779 7945
rect 28721 7905 28733 7939
rect 28767 7905 28779 7939
rect 28721 7899 28779 7905
rect 28813 7939 28871 7945
rect 28813 7905 28825 7939
rect 28859 7936 28871 7939
rect 28994 7936 29000 7948
rect 28859 7908 29000 7936
rect 28859 7905 28871 7908
rect 28813 7899 28871 7905
rect 27856 7896 27862 7899
rect 20640 7840 21956 7868
rect 21266 7800 21272 7812
rect 20548 7772 21272 7800
rect 21266 7760 21272 7772
rect 21324 7760 21330 7812
rect 21928 7800 21956 7840
rect 22922 7828 22928 7880
rect 22980 7868 22986 7880
rect 23017 7871 23075 7877
rect 23017 7868 23029 7871
rect 22980 7840 23029 7868
rect 22980 7828 22986 7840
rect 23017 7837 23029 7840
rect 23063 7837 23075 7871
rect 23017 7831 23075 7837
rect 25406 7828 25412 7880
rect 25464 7828 25470 7880
rect 21468 7772 21864 7800
rect 21928 7772 23060 7800
rect 19521 7735 19579 7741
rect 19521 7732 19533 7735
rect 18840 7704 19533 7732
rect 18840 7692 18846 7704
rect 19521 7701 19533 7704
rect 19567 7732 19579 7735
rect 19981 7735 20039 7741
rect 19981 7732 19993 7735
rect 19567 7704 19993 7732
rect 19567 7701 19579 7704
rect 19521 7695 19579 7701
rect 19981 7701 19993 7704
rect 20027 7701 20039 7735
rect 19981 7695 20039 7701
rect 20162 7692 20168 7744
rect 20220 7732 20226 7744
rect 21468 7741 21496 7772
rect 20441 7735 20499 7741
rect 20441 7732 20453 7735
rect 20220 7704 20453 7732
rect 20220 7692 20226 7704
rect 20441 7701 20453 7704
rect 20487 7701 20499 7735
rect 20441 7695 20499 7701
rect 21453 7735 21511 7741
rect 21453 7701 21465 7735
rect 21499 7701 21511 7735
rect 21453 7695 21511 7701
rect 21634 7692 21640 7744
rect 21692 7732 21698 7744
rect 21729 7735 21787 7741
rect 21729 7732 21741 7735
rect 21692 7704 21741 7732
rect 21692 7692 21698 7704
rect 21729 7701 21741 7704
rect 21775 7701 21787 7735
rect 21836 7732 21864 7772
rect 22278 7732 22284 7744
rect 21836 7704 22284 7732
rect 21729 7695 21787 7701
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 23032 7732 23060 7772
rect 26694 7760 26700 7812
rect 26752 7760 26758 7812
rect 28442 7760 28448 7812
rect 28500 7800 28506 7812
rect 28736 7800 28764 7899
rect 28994 7896 29000 7908
rect 29052 7936 29058 7948
rect 29089 7939 29147 7945
rect 29089 7936 29101 7939
rect 29052 7908 29101 7936
rect 29052 7896 29058 7908
rect 29089 7905 29101 7908
rect 29135 7905 29147 7939
rect 29089 7899 29147 7905
rect 29362 7896 29368 7948
rect 29420 7896 29426 7948
rect 29380 7868 29408 7896
rect 29549 7871 29607 7877
rect 29549 7868 29561 7871
rect 29380 7840 29561 7868
rect 29549 7837 29561 7840
rect 29595 7837 29607 7871
rect 29549 7831 29607 7837
rect 28500 7772 29316 7800
rect 28500 7760 28506 7772
rect 24670 7732 24676 7744
rect 23032 7704 24676 7732
rect 24670 7692 24676 7704
rect 24728 7692 24734 7744
rect 28626 7692 28632 7744
rect 28684 7692 28690 7744
rect 29178 7692 29184 7744
rect 29236 7692 29242 7744
rect 29288 7732 29316 7772
rect 30742 7760 30748 7812
rect 30800 7760 30806 7812
rect 30760 7732 30788 7760
rect 29288 7704 30788 7732
rect 552 7642 31372 7664
rect 552 7590 4250 7642
rect 4302 7590 4314 7642
rect 4366 7590 4378 7642
rect 4430 7590 4442 7642
rect 4494 7590 4506 7642
rect 4558 7590 11955 7642
rect 12007 7590 12019 7642
rect 12071 7590 12083 7642
rect 12135 7590 12147 7642
rect 12199 7590 12211 7642
rect 12263 7590 19660 7642
rect 19712 7590 19724 7642
rect 19776 7590 19788 7642
rect 19840 7590 19852 7642
rect 19904 7590 19916 7642
rect 19968 7590 27365 7642
rect 27417 7590 27429 7642
rect 27481 7590 27493 7642
rect 27545 7590 27557 7642
rect 27609 7590 27621 7642
rect 27673 7590 31372 7642
rect 552 7568 31372 7590
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 2547 7500 11468 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 6178 7420 6184 7472
rect 6236 7460 6242 7472
rect 6273 7463 6331 7469
rect 6273 7460 6285 7463
rect 6236 7432 6285 7460
rect 6236 7420 6242 7432
rect 6273 7429 6285 7432
rect 6319 7460 6331 7463
rect 6319 7432 6684 7460
rect 6319 7429 6331 7432
rect 6273 7423 6331 7429
rect 6546 7392 6552 7404
rect 5736 7364 6552 7392
rect 5736 7336 5764 7364
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 1121 7327 1179 7333
rect 1121 7293 1133 7327
rect 1167 7324 1179 7327
rect 1946 7324 1952 7336
rect 1167 7296 1952 7324
rect 1167 7293 1179 7296
rect 1121 7287 1179 7293
rect 1946 7284 1952 7296
rect 2004 7324 2010 7336
rect 4157 7327 4215 7333
rect 4157 7324 4169 7327
rect 2004 7296 4169 7324
rect 2004 7284 2010 7296
rect 4157 7293 4169 7296
rect 4203 7324 4215 7327
rect 5718 7324 5724 7336
rect 4203 7296 5724 7324
rect 4203 7293 4215 7296
rect 4157 7287 4215 7293
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7324 5871 7327
rect 5994 7324 6000 7336
rect 5859 7296 6000 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 6086 7284 6092 7336
rect 6144 7284 6150 7336
rect 6270 7284 6276 7336
rect 6328 7324 6334 7336
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 6328 7296 6377 7324
rect 6328 7284 6334 7296
rect 6365 7293 6377 7296
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 6454 7284 6460 7336
rect 6512 7284 6518 7336
rect 6656 7324 6684 7432
rect 8018 7420 8024 7472
rect 8076 7460 8082 7472
rect 8113 7463 8171 7469
rect 8113 7460 8125 7463
rect 8076 7432 8125 7460
rect 8076 7420 8082 7432
rect 8113 7429 8125 7432
rect 8159 7429 8171 7463
rect 11440 7460 11468 7500
rect 11514 7488 11520 7540
rect 11572 7528 11578 7540
rect 11609 7531 11667 7537
rect 11609 7528 11621 7531
rect 11572 7500 11621 7528
rect 11572 7488 11578 7500
rect 11609 7497 11621 7500
rect 11655 7497 11667 7531
rect 11609 7491 11667 7497
rect 11793 7531 11851 7537
rect 11793 7497 11805 7531
rect 11839 7528 11851 7531
rect 12894 7528 12900 7540
rect 11839 7500 12900 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 12986 7488 12992 7540
rect 13044 7528 13050 7540
rect 13081 7531 13139 7537
rect 13081 7528 13093 7531
rect 13044 7500 13093 7528
rect 13044 7488 13050 7500
rect 13081 7497 13093 7500
rect 13127 7497 13139 7531
rect 13081 7491 13139 7497
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7528 13323 7531
rect 13906 7528 13912 7540
rect 13311 7500 13912 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 14553 7531 14611 7537
rect 14553 7497 14565 7531
rect 14599 7528 14611 7531
rect 14734 7528 14740 7540
rect 14599 7500 14740 7528
rect 14599 7497 14611 7500
rect 14553 7491 14611 7497
rect 14734 7488 14740 7500
rect 14792 7528 14798 7540
rect 15562 7528 15568 7540
rect 14792 7500 15568 7528
rect 14792 7488 14798 7500
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 16206 7488 16212 7540
rect 16264 7528 16270 7540
rect 19153 7531 19211 7537
rect 19153 7528 19165 7531
rect 16264 7500 19165 7528
rect 16264 7488 16270 7500
rect 19153 7497 19165 7500
rect 19199 7497 19211 7531
rect 21450 7528 21456 7540
rect 19153 7491 19211 7497
rect 21169 7500 21456 7528
rect 11440 7432 13584 7460
rect 8113 7423 8171 7429
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 8754 7352 8760 7404
rect 8812 7392 8818 7404
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 8812 7364 8953 7392
rect 8812 7352 8818 7364
rect 8941 7361 8953 7364
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 6656 7296 8861 7324
rect 8849 7293 8861 7296
rect 8895 7324 8907 7327
rect 10413 7327 10471 7333
rect 8895 7296 8984 7324
rect 8895 7293 8907 7296
rect 8849 7287 8907 7293
rect 1394 7265 1400 7268
rect 1388 7256 1400 7265
rect 1355 7228 1400 7256
rect 1388 7219 1400 7228
rect 1394 7216 1400 7219
rect 1452 7216 1458 7268
rect 4424 7259 4482 7265
rect 4424 7225 4436 7259
rect 4470 7256 4482 7259
rect 5626 7256 5632 7268
rect 4470 7228 5632 7256
rect 4470 7225 4482 7228
rect 4424 7219 4482 7225
rect 5626 7216 5632 7228
rect 5684 7216 5690 7268
rect 6978 7259 7036 7265
rect 6978 7256 6990 7259
rect 5736 7228 6990 7256
rect 5534 7148 5540 7200
rect 5592 7148 5598 7200
rect 5736 7197 5764 7228
rect 6978 7225 6990 7228
rect 7024 7256 7036 7259
rect 7190 7256 7196 7268
rect 7024 7228 7196 7256
rect 7024 7225 7036 7228
rect 6978 7219 7036 7225
rect 7190 7216 7196 7228
rect 7248 7216 7254 7268
rect 8018 7216 8024 7268
rect 8076 7256 8082 7268
rect 8956 7256 8984 7296
rect 10413 7293 10425 7327
rect 10459 7324 10471 7327
rect 12434 7324 12440 7336
rect 10459 7296 12440 7324
rect 10459 7293 10471 7296
rect 10413 7287 10471 7293
rect 9186 7259 9244 7265
rect 9186 7256 9198 7259
rect 8076 7228 8892 7256
rect 8956 7228 9198 7256
rect 8076 7216 8082 7228
rect 5721 7191 5779 7197
rect 5721 7157 5733 7191
rect 5767 7157 5779 7191
rect 5721 7151 5779 7157
rect 6546 7148 6552 7200
rect 6604 7148 6610 7200
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 8757 7191 8815 7197
rect 8757 7188 8769 7191
rect 8720 7160 8769 7188
rect 8720 7148 8726 7160
rect 8757 7157 8769 7160
rect 8803 7157 8815 7191
rect 8864 7188 8892 7228
rect 9186 7225 9198 7228
rect 9232 7225 9244 7259
rect 10428 7256 10456 7287
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 13446 7324 13452 7336
rect 13162 7299 13452 7324
rect 13127 7296 13452 7299
rect 13127 7293 13190 7296
rect 9186 7219 9244 7225
rect 9324 7228 10456 7256
rect 9324 7188 9352 7228
rect 10962 7216 10968 7268
rect 11020 7256 11026 7268
rect 11149 7259 11207 7265
rect 11149 7256 11161 7259
rect 11020 7228 11161 7256
rect 11020 7216 11026 7228
rect 11149 7225 11161 7228
rect 11195 7225 11207 7259
rect 11149 7219 11207 7225
rect 11238 7216 11244 7268
rect 11296 7256 11302 7268
rect 11425 7259 11483 7265
rect 11425 7256 11437 7259
rect 11296 7228 11437 7256
rect 11296 7216 11302 7228
rect 11425 7225 11437 7228
rect 11471 7225 11483 7259
rect 12897 7259 12955 7265
rect 12897 7256 12909 7259
rect 11425 7219 11483 7225
rect 11532 7228 12909 7256
rect 8864 7160 9352 7188
rect 10321 7191 10379 7197
rect 8757 7151 8815 7157
rect 10321 7157 10333 7191
rect 10367 7188 10379 7191
rect 11532 7188 11560 7228
rect 12897 7225 12909 7228
rect 12943 7225 12955 7259
rect 13127 7259 13139 7293
rect 13173 7262 13190 7293
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 13173 7259 13185 7262
rect 13127 7253 13185 7259
rect 13556 7256 13584 7432
rect 15194 7420 15200 7472
rect 15252 7460 15258 7472
rect 15289 7463 15347 7469
rect 15289 7460 15301 7463
rect 15252 7432 15301 7460
rect 15252 7420 15258 7432
rect 15289 7429 15301 7432
rect 15335 7460 15347 7463
rect 16298 7460 16304 7472
rect 15335 7432 16304 7460
rect 15335 7429 15347 7432
rect 15289 7423 15347 7429
rect 16298 7420 16304 7432
rect 16356 7420 16362 7472
rect 16390 7420 16396 7472
rect 16448 7460 16454 7472
rect 16485 7463 16543 7469
rect 16485 7460 16497 7463
rect 16448 7432 16497 7460
rect 16448 7420 16454 7432
rect 16485 7429 16497 7432
rect 16531 7429 16543 7463
rect 16485 7423 16543 7429
rect 18049 7463 18107 7469
rect 18049 7429 18061 7463
rect 18095 7460 18107 7463
rect 18322 7460 18328 7472
rect 18095 7432 18328 7460
rect 18095 7429 18107 7432
rect 18049 7423 18107 7429
rect 18322 7420 18328 7432
rect 18380 7420 18386 7472
rect 14550 7352 14556 7404
rect 14608 7392 14614 7404
rect 14921 7395 14979 7401
rect 14921 7392 14933 7395
rect 14608 7364 14933 7392
rect 14608 7352 14614 7364
rect 14921 7361 14933 7364
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7392 15899 7395
rect 21169 7392 21197 7500
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 21637 7531 21695 7537
rect 21637 7497 21649 7531
rect 21683 7528 21695 7531
rect 21726 7528 21732 7540
rect 21683 7500 21732 7528
rect 21683 7497 21695 7500
rect 21637 7491 21695 7497
rect 21726 7488 21732 7500
rect 21784 7488 21790 7540
rect 21818 7488 21824 7540
rect 21876 7528 21882 7540
rect 21913 7531 21971 7537
rect 21913 7528 21925 7531
rect 21876 7500 21925 7528
rect 21876 7488 21882 7500
rect 21913 7497 21925 7500
rect 21959 7497 21971 7531
rect 21913 7491 21971 7497
rect 22186 7488 22192 7540
rect 22244 7528 22250 7540
rect 22465 7531 22523 7537
rect 22465 7528 22477 7531
rect 22244 7500 22477 7528
rect 22244 7488 22250 7500
rect 22465 7497 22477 7500
rect 22511 7497 22523 7531
rect 26145 7531 26203 7537
rect 26145 7528 26157 7531
rect 22465 7491 22523 7497
rect 23190 7500 26157 7528
rect 21266 7420 21272 7472
rect 21324 7460 21330 7472
rect 23190 7460 23218 7500
rect 26145 7497 26157 7500
rect 26191 7497 26203 7531
rect 26145 7491 26203 7497
rect 27798 7488 27804 7540
rect 27856 7528 27862 7540
rect 28537 7531 28595 7537
rect 28537 7528 28549 7531
rect 27856 7500 28549 7528
rect 27856 7488 27862 7500
rect 28537 7497 28549 7500
rect 28583 7497 28595 7531
rect 28537 7491 28595 7497
rect 30282 7488 30288 7540
rect 30340 7488 30346 7540
rect 30742 7488 30748 7540
rect 30800 7528 30806 7540
rect 30929 7531 30987 7537
rect 30929 7528 30941 7531
rect 30800 7500 30941 7528
rect 30800 7488 30806 7500
rect 30929 7497 30941 7500
rect 30975 7497 30987 7531
rect 30929 7491 30987 7497
rect 21324 7432 23218 7460
rect 21324 7420 21330 7432
rect 24670 7420 24676 7472
rect 24728 7420 24734 7472
rect 15887 7364 17448 7392
rect 15887 7361 15899 7364
rect 15841 7355 15899 7361
rect 14274 7284 14280 7336
rect 14332 7284 14338 7336
rect 15933 7327 15991 7333
rect 15933 7293 15945 7327
rect 15979 7293 15991 7327
rect 15933 7287 15991 7293
rect 16025 7327 16083 7333
rect 16025 7293 16037 7327
rect 16071 7324 16083 7327
rect 16482 7324 16488 7336
rect 16071 7296 16488 7324
rect 16071 7293 16083 7296
rect 16025 7287 16083 7293
rect 14369 7259 14427 7265
rect 14369 7256 14381 7259
rect 13556 7228 14381 7256
rect 12897 7219 12955 7225
rect 14369 7225 14381 7228
rect 14415 7225 14427 7259
rect 15105 7259 15163 7265
rect 14369 7219 14427 7225
rect 14584 7228 15056 7256
rect 10367 7160 11560 7188
rect 10367 7157 10379 7160
rect 10321 7151 10379 7157
rect 11606 7148 11612 7200
rect 11664 7197 11670 7200
rect 11664 7191 11683 7197
rect 11671 7157 11683 7191
rect 11664 7151 11683 7157
rect 11664 7148 11670 7151
rect 12710 7148 12716 7200
rect 12768 7188 12774 7200
rect 14584 7197 14612 7228
rect 14093 7191 14151 7197
rect 14093 7188 14105 7191
rect 12768 7160 14105 7188
rect 12768 7148 12774 7160
rect 14093 7157 14105 7160
rect 14139 7188 14151 7191
rect 14569 7191 14627 7197
rect 14569 7188 14581 7191
rect 14139 7160 14581 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 14569 7157 14581 7160
rect 14615 7157 14627 7191
rect 14569 7151 14627 7157
rect 14734 7148 14740 7200
rect 14792 7148 14798 7200
rect 15028 7188 15056 7228
rect 15105 7225 15117 7259
rect 15151 7256 15163 7259
rect 15473 7259 15531 7265
rect 15473 7256 15485 7259
rect 15151 7228 15485 7256
rect 15151 7225 15163 7228
rect 15105 7219 15163 7225
rect 15473 7225 15485 7228
rect 15519 7256 15531 7259
rect 15657 7259 15715 7265
rect 15657 7256 15669 7259
rect 15519 7228 15669 7256
rect 15519 7225 15531 7228
rect 15473 7219 15531 7225
rect 15657 7225 15669 7228
rect 15703 7225 15715 7259
rect 15948 7256 15976 7287
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 16666 7284 16672 7336
rect 16724 7284 16730 7336
rect 17218 7284 17224 7336
rect 17276 7284 17282 7336
rect 17310 7284 17316 7336
rect 17368 7284 17374 7336
rect 17420 7333 17448 7364
rect 20456 7364 21197 7392
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7324 17463 7327
rect 17678 7324 17684 7336
rect 17451 7296 17684 7324
rect 17451 7293 17463 7296
rect 17405 7287 17463 7293
rect 17678 7284 17684 7296
rect 17736 7284 17742 7336
rect 20277 7327 20335 7333
rect 20277 7293 20289 7327
rect 20323 7324 20335 7327
rect 20456 7324 20484 7364
rect 21910 7352 21916 7404
rect 21968 7392 21974 7404
rect 27525 7395 27583 7401
rect 21968 7364 23704 7392
rect 21968 7352 21974 7364
rect 20323 7296 20484 7324
rect 20533 7327 20591 7333
rect 20323 7293 20335 7296
rect 20277 7287 20335 7293
rect 20533 7293 20545 7327
rect 20579 7324 20591 7327
rect 20579 7296 20852 7324
rect 20579 7293 20591 7296
rect 20533 7287 20591 7293
rect 17236 7256 17264 7284
rect 15948 7228 17264 7256
rect 17328 7256 17356 7284
rect 17773 7259 17831 7265
rect 17773 7256 17785 7259
rect 17328 7228 17785 7256
rect 15657 7219 15715 7225
rect 17773 7225 17785 7228
rect 17819 7225 17831 7259
rect 17773 7219 17831 7225
rect 20824 7256 20852 7296
rect 21174 7284 21180 7336
rect 21232 7284 21238 7336
rect 21450 7284 21456 7336
rect 21508 7284 21514 7336
rect 21542 7284 21548 7336
rect 21600 7284 21606 7336
rect 21818 7284 21824 7336
rect 21876 7324 21882 7336
rect 22005 7327 22063 7333
rect 22005 7324 22017 7327
rect 21876 7296 22017 7324
rect 21876 7284 21882 7296
rect 22005 7293 22017 7296
rect 22051 7324 22063 7327
rect 22281 7327 22339 7333
rect 22281 7324 22293 7327
rect 22051 7296 22293 7324
rect 22051 7293 22063 7296
rect 22005 7287 22063 7293
rect 22281 7293 22293 7296
rect 22327 7293 22339 7327
rect 22281 7287 22339 7293
rect 22370 7284 22376 7336
rect 22428 7284 22434 7336
rect 23676 7333 23704 7364
rect 27525 7361 27537 7395
rect 27571 7392 27583 7395
rect 27890 7392 27896 7404
rect 27571 7364 27896 7392
rect 27571 7361 27583 7364
rect 27525 7355 27583 7361
rect 23661 7327 23719 7333
rect 23661 7293 23673 7327
rect 23707 7324 23719 7327
rect 25958 7324 25964 7336
rect 23707 7296 25964 7324
rect 23707 7293 23719 7296
rect 23661 7287 23719 7293
rect 25958 7284 25964 7296
rect 26016 7284 26022 7336
rect 26053 7327 26111 7333
rect 26053 7293 26065 7327
rect 26099 7324 26111 7327
rect 27540 7324 27568 7355
rect 27890 7352 27896 7364
rect 27948 7352 27954 7404
rect 27985 7395 28043 7401
rect 27985 7361 27997 7395
rect 28031 7392 28043 7395
rect 28902 7392 28908 7404
rect 28031 7364 28908 7392
rect 28031 7361 28043 7364
rect 27985 7355 28043 7361
rect 28902 7352 28908 7364
rect 28960 7392 28966 7404
rect 29089 7395 29147 7401
rect 29089 7392 29101 7395
rect 28960 7364 29101 7392
rect 28960 7352 28966 7364
rect 29089 7361 29101 7364
rect 29135 7361 29147 7395
rect 29089 7355 29147 7361
rect 26099 7296 27568 7324
rect 28077 7327 28135 7333
rect 26099 7293 26111 7296
rect 26053 7287 26111 7293
rect 28077 7293 28089 7327
rect 28123 7324 28135 7327
rect 28442 7324 28448 7336
rect 28123 7296 28448 7324
rect 28123 7293 28135 7296
rect 28077 7287 28135 7293
rect 28442 7284 28448 7296
rect 28500 7284 28506 7336
rect 28721 7327 28779 7333
rect 28721 7324 28733 7327
rect 28552 7296 28733 7324
rect 22922 7256 22928 7268
rect 20824 7228 22928 7256
rect 20824 7200 20852 7228
rect 22922 7216 22928 7228
rect 22980 7216 22986 7268
rect 25808 7259 25866 7265
rect 25808 7225 25820 7259
rect 25854 7256 25866 7259
rect 27280 7259 27338 7265
rect 25854 7228 26096 7256
rect 25854 7225 25866 7228
rect 25808 7219 25866 7225
rect 26068 7200 26096 7228
rect 27280 7225 27292 7259
rect 27326 7256 27338 7259
rect 27522 7256 27528 7268
rect 27326 7228 27528 7256
rect 27326 7225 27338 7228
rect 27280 7219 27338 7225
rect 27522 7216 27528 7228
rect 27580 7216 27586 7268
rect 28552 7200 28580 7296
rect 28721 7293 28733 7296
rect 28767 7293 28779 7327
rect 28721 7287 28779 7293
rect 29181 7327 29239 7333
rect 29181 7293 29193 7327
rect 29227 7293 29239 7327
rect 29181 7287 29239 7293
rect 29457 7327 29515 7333
rect 29457 7293 29469 7327
rect 29503 7324 29515 7327
rect 29730 7324 29736 7336
rect 29503 7296 29736 7324
rect 29503 7293 29515 7296
rect 29457 7287 29515 7293
rect 29196 7256 29224 7287
rect 29730 7284 29736 7296
rect 29788 7284 29794 7336
rect 30466 7333 30472 7336
rect 30461 7324 30472 7333
rect 30427 7296 30472 7324
rect 30461 7287 30472 7296
rect 30466 7284 30472 7287
rect 30524 7284 30530 7336
rect 30558 7284 30564 7336
rect 30616 7284 30622 7336
rect 30837 7327 30895 7333
rect 30837 7293 30849 7327
rect 30883 7293 30895 7327
rect 30837 7287 30895 7293
rect 29196 7228 29868 7256
rect 29840 7200 29868 7228
rect 30742 7216 30748 7268
rect 30800 7256 30806 7268
rect 30852 7256 30880 7287
rect 30800 7228 30880 7256
rect 30800 7216 30806 7228
rect 19242 7188 19248 7200
rect 15028 7160 19248 7188
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 20806 7148 20812 7200
rect 20864 7148 20870 7200
rect 21085 7191 21143 7197
rect 21085 7157 21097 7191
rect 21131 7188 21143 7191
rect 21361 7191 21419 7197
rect 21361 7188 21373 7191
rect 21131 7160 21373 7188
rect 21131 7157 21143 7160
rect 21085 7151 21143 7157
rect 21361 7157 21373 7160
rect 21407 7188 21419 7191
rect 21542 7188 21548 7200
rect 21407 7160 21548 7188
rect 21407 7157 21419 7160
rect 21361 7151 21419 7157
rect 21542 7148 21548 7160
rect 21600 7148 21606 7200
rect 23198 7148 23204 7200
rect 23256 7188 23262 7200
rect 24394 7188 24400 7200
rect 23256 7160 24400 7188
rect 23256 7148 23262 7160
rect 24394 7148 24400 7160
rect 24452 7148 24458 7200
rect 26050 7148 26056 7200
rect 26108 7148 26114 7200
rect 28534 7148 28540 7200
rect 28592 7148 28598 7200
rect 29270 7148 29276 7200
rect 29328 7148 29334 7200
rect 29822 7148 29828 7200
rect 29880 7148 29886 7200
rect 30650 7148 30656 7200
rect 30708 7148 30714 7200
rect 552 7098 31531 7120
rect 552 7046 8102 7098
rect 8154 7046 8166 7098
rect 8218 7046 8230 7098
rect 8282 7046 8294 7098
rect 8346 7046 8358 7098
rect 8410 7046 15807 7098
rect 15859 7046 15871 7098
rect 15923 7046 15935 7098
rect 15987 7046 15999 7098
rect 16051 7046 16063 7098
rect 16115 7046 23512 7098
rect 23564 7046 23576 7098
rect 23628 7046 23640 7098
rect 23692 7046 23704 7098
rect 23756 7046 23768 7098
rect 23820 7046 31217 7098
rect 31269 7046 31281 7098
rect 31333 7046 31345 7098
rect 31397 7046 31409 7098
rect 31461 7046 31473 7098
rect 31525 7046 31531 7098
rect 552 7024 31531 7046
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 5592 6956 8616 6984
rect 5592 6944 5598 6956
rect 5626 6876 5632 6928
rect 5684 6916 5690 6928
rect 6546 6916 6552 6928
rect 5684 6888 6552 6916
rect 5684 6876 5690 6888
rect 1946 6808 1952 6860
rect 2004 6848 2010 6860
rect 2133 6851 2191 6857
rect 2133 6848 2145 6851
rect 2004 6820 2145 6848
rect 2004 6808 2010 6820
rect 2133 6817 2145 6820
rect 2179 6817 2191 6851
rect 2133 6811 2191 6817
rect 2222 6808 2228 6860
rect 2280 6848 2286 6860
rect 5828 6857 5856 6888
rect 6546 6876 6552 6888
rect 6604 6876 6610 6928
rect 7190 6876 7196 6928
rect 7248 6876 7254 6928
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 8018 6916 8024 6928
rect 7340 6888 8024 6916
rect 7340 6876 7346 6888
rect 8018 6876 8024 6888
rect 8076 6876 8082 6928
rect 8588 6916 8616 6956
rect 8662 6944 8668 6996
rect 8720 6944 8726 6996
rect 12739 6987 12797 6993
rect 9646 6956 12664 6984
rect 9646 6916 9674 6956
rect 8588 6888 9674 6916
rect 12526 6876 12532 6928
rect 12584 6876 12590 6928
rect 12636 6916 12664 6956
rect 12739 6953 12751 6987
rect 12785 6984 12797 6987
rect 13446 6984 13452 6996
rect 12785 6956 13452 6984
rect 12785 6953 12797 6956
rect 12739 6947 12797 6953
rect 13446 6944 13452 6956
rect 13504 6984 13510 6996
rect 13906 6984 13912 6996
rect 13504 6956 13912 6984
rect 13504 6944 13510 6956
rect 13906 6944 13912 6956
rect 13964 6944 13970 6996
rect 14642 6944 14648 6996
rect 14700 6984 14706 6996
rect 14737 6987 14795 6993
rect 14737 6984 14749 6987
rect 14700 6956 14749 6984
rect 14700 6944 14706 6956
rect 14737 6953 14749 6956
rect 14783 6953 14795 6987
rect 14737 6947 14795 6953
rect 15286 6944 15292 6996
rect 15344 6984 15350 6996
rect 15344 6956 16441 6984
rect 15344 6944 15350 6956
rect 13262 6916 13268 6928
rect 12636 6888 13268 6916
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 14274 6876 14280 6928
rect 14332 6916 14338 6928
rect 14553 6919 14611 6925
rect 14553 6916 14565 6919
rect 14332 6888 14565 6916
rect 14332 6876 14338 6888
rect 14553 6885 14565 6888
rect 14599 6916 14611 6919
rect 15654 6916 15660 6928
rect 14599 6888 15660 6916
rect 14599 6885 14611 6888
rect 14553 6879 14611 6885
rect 15654 6876 15660 6888
rect 15712 6916 15718 6928
rect 16413 6916 16441 6956
rect 16482 6944 16488 6996
rect 16540 6984 16546 6996
rect 16577 6987 16635 6993
rect 16577 6984 16589 6987
rect 16540 6956 16589 6984
rect 16540 6944 16546 6956
rect 16577 6953 16589 6956
rect 16623 6984 16635 6987
rect 16758 6984 16764 6996
rect 16623 6956 16764 6984
rect 16623 6953 16635 6956
rect 16577 6947 16635 6953
rect 16758 6944 16764 6956
rect 16816 6944 16822 6996
rect 17218 6944 17224 6996
rect 17276 6984 17282 6996
rect 17276 6956 17816 6984
rect 17276 6944 17282 6956
rect 17126 6916 17132 6928
rect 15712 6888 15976 6916
rect 16413 6888 17132 6916
rect 15712 6876 15718 6888
rect 2389 6851 2447 6857
rect 2389 6848 2401 6851
rect 2280 6820 2401 6848
rect 2280 6808 2286 6820
rect 2389 6817 2401 6820
rect 2435 6817 2447 6851
rect 2389 6811 2447 6817
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6817 5871 6851
rect 5813 6811 5871 6817
rect 6178 6808 6184 6860
rect 6236 6848 6242 6860
rect 6273 6851 6331 6857
rect 6273 6848 6285 6851
rect 6236 6820 6285 6848
rect 6236 6808 6242 6820
rect 6273 6817 6285 6820
rect 6319 6817 6331 6851
rect 7208 6848 7236 6876
rect 15948 6860 15976 6888
rect 17126 6876 17132 6888
rect 17184 6876 17190 6928
rect 7466 6848 7472 6860
rect 7208 6820 7472 6848
rect 6273 6811 6331 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7561 6851 7619 6857
rect 7561 6817 7573 6851
rect 7607 6848 7619 6851
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7607 6820 7665 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 6914 6780 6920 6792
rect 6595 6752 6920 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 5905 6715 5963 6721
rect 5905 6681 5917 6715
rect 5951 6712 5963 6715
rect 6181 6715 6239 6721
rect 6181 6712 6193 6715
rect 5951 6684 6193 6712
rect 5951 6681 5963 6684
rect 5905 6675 5963 6681
rect 6181 6681 6193 6684
rect 6227 6712 6239 6715
rect 7576 6712 7604 6811
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 7800 6820 8309 6848
rect 7800 6808 7806 6820
rect 8297 6817 8309 6820
rect 8343 6848 8355 6851
rect 8573 6851 8631 6857
rect 8573 6848 8585 6851
rect 8343 6820 8585 6848
rect 8343 6817 8355 6820
rect 8297 6811 8355 6817
rect 8573 6817 8585 6820
rect 8619 6817 8631 6851
rect 8573 6811 8631 6817
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 8720 6820 9045 6848
rect 8720 6808 8726 6820
rect 9033 6817 9045 6820
rect 9079 6848 9091 6851
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 9079 6820 9321 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 11221 6851 11279 6857
rect 11221 6848 11233 6851
rect 10560 6820 11233 6848
rect 10560 6808 10566 6820
rect 11221 6817 11233 6820
rect 11267 6817 11279 6851
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 11221 6811 11279 6817
rect 12636 6820 13645 6848
rect 6227 6684 7604 6712
rect 7668 6752 10916 6780
rect 6227 6681 6239 6684
rect 6181 6675 6239 6681
rect 3510 6604 3516 6656
rect 3568 6604 3574 6656
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 7668 6644 7696 6752
rect 7745 6715 7803 6721
rect 7745 6681 7757 6715
rect 7791 6712 7803 6715
rect 8846 6712 8852 6724
rect 7791 6684 8852 6712
rect 7791 6681 7803 6684
rect 7745 6675 7803 6681
rect 8846 6672 8852 6684
rect 8904 6712 8910 6724
rect 9401 6715 9459 6721
rect 9401 6712 9413 6715
rect 8904 6684 9413 6712
rect 8904 6672 8910 6684
rect 9401 6681 9413 6684
rect 9447 6681 9459 6715
rect 9401 6675 9459 6681
rect 3660 6616 7696 6644
rect 8389 6647 8447 6653
rect 3660 6604 3666 6616
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8478 6644 8484 6656
rect 8435 6616 8484 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8478 6604 8484 6616
rect 8536 6644 8542 6656
rect 8938 6644 8944 6656
rect 8536 6616 8944 6644
rect 8536 6604 8542 6616
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9125 6647 9183 6653
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 10318 6644 10324 6656
rect 9171 6616 10324 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 10888 6644 10916 6752
rect 10962 6740 10968 6792
rect 11020 6740 11026 6792
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 12345 6715 12403 6721
rect 12345 6712 12357 6715
rect 12308 6684 12357 6712
rect 12308 6672 12314 6684
rect 12345 6681 12357 6684
rect 12391 6681 12403 6715
rect 12345 6675 12403 6681
rect 12636 6644 12664 6820
rect 13633 6817 13645 6820
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 13814 6808 13820 6860
rect 13872 6808 13878 6860
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 14056 6820 14197 6848
rect 14056 6808 14062 6820
rect 14185 6817 14197 6820
rect 14231 6817 14243 6851
rect 14185 6811 14243 6817
rect 14734 6808 14740 6860
rect 14792 6848 14798 6860
rect 15197 6851 15255 6857
rect 15197 6848 15209 6851
rect 14792 6820 15209 6848
rect 14792 6808 14798 6820
rect 15197 6817 15209 6820
rect 15243 6817 15255 6851
rect 15197 6811 15255 6817
rect 15286 6808 15292 6860
rect 15344 6808 15350 6860
rect 15473 6851 15531 6857
rect 15473 6817 15485 6851
rect 15519 6817 15531 6851
rect 15473 6811 15531 6817
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 12768 6752 12940 6780
rect 12768 6740 12774 6752
rect 12912 6721 12940 6752
rect 13078 6740 13084 6792
rect 13136 6740 13142 6792
rect 14826 6780 14832 6792
rect 13280 6752 14832 6780
rect 12897 6715 12955 6721
rect 12897 6681 12909 6715
rect 12943 6681 12955 6715
rect 12897 6675 12955 6681
rect 10888 6616 12664 6644
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 13280 6644 13308 6752
rect 14826 6740 14832 6752
rect 14884 6780 14890 6792
rect 15488 6780 15516 6811
rect 15930 6808 15936 6860
rect 15988 6808 15994 6860
rect 16114 6808 16120 6860
rect 16172 6808 16178 6860
rect 16209 6851 16267 6857
rect 16209 6817 16221 6851
rect 16255 6848 16267 6851
rect 17236 6848 17264 6944
rect 17310 6876 17316 6928
rect 17368 6916 17374 6928
rect 17405 6919 17463 6925
rect 17405 6916 17417 6919
rect 17368 6888 17417 6916
rect 17368 6876 17374 6888
rect 17405 6885 17417 6888
rect 17451 6885 17463 6919
rect 17405 6879 17463 6885
rect 17788 6860 17816 6956
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 19505 6987 19563 6993
rect 18380 6956 19012 6984
rect 18380 6944 18386 6956
rect 16255 6820 17264 6848
rect 16255 6817 16267 6820
rect 16209 6811 16267 6817
rect 17494 6808 17500 6860
rect 17552 6848 17558 6860
rect 17681 6851 17739 6857
rect 17681 6848 17693 6851
rect 17552 6820 17693 6848
rect 17552 6808 17558 6820
rect 17681 6817 17693 6820
rect 17727 6817 17739 6851
rect 17681 6811 17739 6817
rect 17770 6808 17776 6860
rect 17828 6848 17834 6860
rect 18141 6851 18199 6857
rect 18141 6848 18153 6851
rect 17828 6820 18153 6848
rect 17828 6808 17834 6820
rect 18141 6817 18153 6820
rect 18187 6817 18199 6851
rect 18141 6811 18199 6817
rect 18506 6808 18512 6860
rect 18564 6808 18570 6860
rect 18984 6857 19012 6956
rect 19505 6953 19517 6987
rect 19551 6984 19563 6987
rect 20530 6984 20536 6996
rect 19551 6956 20536 6984
rect 19551 6953 19563 6956
rect 19505 6947 19563 6953
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 21542 6944 21548 6996
rect 21600 6944 21606 6996
rect 27522 6944 27528 6996
rect 27580 6984 27586 6996
rect 27706 6984 27712 6996
rect 27580 6956 27712 6984
rect 27580 6944 27586 6956
rect 27706 6944 27712 6956
rect 27764 6984 27770 6996
rect 27801 6987 27859 6993
rect 27801 6984 27813 6987
rect 27764 6956 27813 6984
rect 27764 6944 27770 6956
rect 27801 6953 27813 6956
rect 27847 6953 27859 6987
rect 27801 6947 27859 6953
rect 27890 6944 27896 6996
rect 27948 6944 27954 6996
rect 29178 6944 29184 6996
rect 29236 6984 29242 6996
rect 30101 6987 30159 6993
rect 30101 6984 30113 6987
rect 29236 6956 30113 6984
rect 29236 6944 29242 6956
rect 30101 6953 30113 6956
rect 30147 6984 30159 6987
rect 30558 6984 30564 6996
rect 30147 6956 30564 6984
rect 30147 6953 30159 6956
rect 30101 6947 30159 6953
rect 30558 6944 30564 6956
rect 30616 6944 30622 6996
rect 30650 6944 30656 6996
rect 30708 6944 30714 6996
rect 19702 6876 19708 6928
rect 19760 6876 19766 6928
rect 21560 6857 21588 6944
rect 23842 6876 23848 6928
rect 23900 6916 23906 6928
rect 24394 6916 24400 6928
rect 23900 6888 24400 6916
rect 23900 6876 23906 6888
rect 24394 6876 24400 6888
rect 24452 6876 24458 6928
rect 25958 6876 25964 6928
rect 26016 6916 26022 6928
rect 26421 6919 26479 6925
rect 26421 6916 26433 6919
rect 26016 6888 26433 6916
rect 26016 6876 26022 6888
rect 26421 6885 26433 6888
rect 26467 6885 26479 6919
rect 26421 6879 26479 6885
rect 27249 6919 27307 6925
rect 27249 6885 27261 6919
rect 27295 6916 27307 6919
rect 27908 6916 27936 6944
rect 27295 6888 27936 6916
rect 27295 6885 27307 6888
rect 27249 6879 27307 6885
rect 28626 6876 28632 6928
rect 28684 6916 28690 6928
rect 28684 6888 29132 6916
rect 28684 6876 28690 6888
rect 18969 6851 19027 6857
rect 18969 6817 18981 6851
rect 19015 6817 19027 6851
rect 18969 6811 19027 6817
rect 21545 6851 21603 6857
rect 21545 6817 21557 6851
rect 21591 6817 21603 6851
rect 21545 6811 21603 6817
rect 22005 6851 22063 6857
rect 22005 6817 22017 6851
rect 22051 6817 22063 6851
rect 22005 6811 22063 6817
rect 16132 6780 16160 6808
rect 14884 6752 15424 6780
rect 15488 6752 16160 6780
rect 14884 6740 14890 6752
rect 14550 6672 14556 6724
rect 14608 6712 14614 6724
rect 15013 6715 15071 6721
rect 15013 6712 15025 6715
rect 14608 6684 15025 6712
rect 14608 6672 14614 6684
rect 15013 6681 15025 6684
rect 15059 6681 15071 6715
rect 15013 6675 15071 6681
rect 12768 6616 13308 6644
rect 12768 6604 12774 6616
rect 13354 6604 13360 6656
rect 13412 6604 13418 6656
rect 13446 6604 13452 6656
rect 13504 6604 13510 6656
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 14182 6644 14188 6656
rect 13587 6616 14188 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 15102 6604 15108 6656
rect 15160 6604 15166 6656
rect 15396 6644 15424 6752
rect 16758 6740 16764 6792
rect 16816 6780 16822 6792
rect 17512 6780 17540 6808
rect 16816 6752 17540 6780
rect 16816 6740 16822 6752
rect 18874 6740 18880 6792
rect 18932 6740 18938 6792
rect 17589 6715 17647 6721
rect 16592 6684 16887 6712
rect 16298 6644 16304 6656
rect 15396 6616 16304 6644
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 16592 6653 16620 6684
rect 16577 6647 16635 6653
rect 16577 6613 16589 6647
rect 16623 6613 16635 6647
rect 16577 6607 16635 6613
rect 16758 6604 16764 6656
rect 16816 6604 16822 6656
rect 16859 6644 16887 6684
rect 17589 6681 17601 6715
rect 17635 6712 17647 6715
rect 18984 6712 19012 6811
rect 21450 6740 21456 6792
rect 21508 6780 21514 6792
rect 21913 6783 21971 6789
rect 21913 6780 21925 6783
rect 21508 6752 21925 6780
rect 21508 6740 21514 6752
rect 21913 6749 21925 6752
rect 21959 6749 21971 6783
rect 22020 6780 22048 6811
rect 22278 6808 22284 6860
rect 22336 6808 22342 6860
rect 22557 6851 22615 6857
rect 22557 6817 22569 6851
rect 22603 6817 22615 6851
rect 22557 6811 22615 6817
rect 22094 6780 22100 6792
rect 22020 6752 22100 6780
rect 21913 6743 21971 6749
rect 19058 6712 19064 6724
rect 17635 6684 17816 6712
rect 18984 6684 19064 6712
rect 17635 6681 17647 6684
rect 17589 6675 17647 6681
rect 17678 6644 17684 6656
rect 16859 6616 17684 6644
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 17788 6644 17816 6684
rect 19058 6672 19064 6684
rect 19116 6712 19122 6724
rect 20162 6712 20168 6724
rect 19116 6684 20168 6712
rect 19116 6672 19122 6684
rect 17862 6644 17868 6656
rect 17788 6616 17868 6644
rect 17862 6604 17868 6616
rect 17920 6604 17926 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 19536 6653 19564 6684
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 21174 6672 21180 6724
rect 21232 6712 21238 6724
rect 21928 6712 21956 6743
rect 22094 6740 22100 6752
rect 22152 6780 22158 6792
rect 22465 6783 22523 6789
rect 22465 6780 22477 6783
rect 22152 6752 22477 6780
rect 22152 6740 22158 6752
rect 22465 6749 22477 6752
rect 22511 6749 22523 6783
rect 22465 6743 22523 6749
rect 22189 6715 22247 6721
rect 22189 6712 22201 6715
rect 21232 6684 21864 6712
rect 21928 6684 22201 6712
rect 21232 6672 21238 6684
rect 19337 6647 19395 6653
rect 19337 6644 19349 6647
rect 18012 6616 19349 6644
rect 18012 6604 18018 6616
rect 19337 6613 19349 6616
rect 19383 6613 19395 6647
rect 19337 6607 19395 6613
rect 19521 6647 19579 6653
rect 19521 6613 19533 6647
rect 19567 6613 19579 6647
rect 19521 6607 19579 6613
rect 21634 6604 21640 6656
rect 21692 6604 21698 6656
rect 21836 6644 21864 6684
rect 22189 6681 22201 6684
rect 22235 6712 22247 6715
rect 22370 6712 22376 6724
rect 22235 6684 22376 6712
rect 22235 6681 22247 6684
rect 22189 6675 22247 6681
rect 22370 6672 22376 6684
rect 22428 6672 22434 6724
rect 22572 6644 22600 6811
rect 23934 6808 23940 6860
rect 23992 6857 23998 6860
rect 23992 6848 24004 6857
rect 23992 6820 24037 6848
rect 23992 6811 24004 6820
rect 23992 6808 23998 6811
rect 26234 6808 26240 6860
rect 26292 6808 26298 6860
rect 27617 6851 27675 6857
rect 27617 6817 27629 6851
rect 27663 6848 27675 6851
rect 27798 6848 27804 6860
rect 27663 6820 27804 6848
rect 27663 6817 27675 6820
rect 27617 6811 27675 6817
rect 27798 6808 27804 6820
rect 27856 6808 27862 6860
rect 27893 6851 27951 6857
rect 27893 6817 27905 6851
rect 27939 6848 27951 6851
rect 28261 6851 28319 6857
rect 28261 6848 28273 6851
rect 27939 6820 28273 6848
rect 27939 6817 27951 6820
rect 27893 6811 27951 6817
rect 28261 6817 28273 6820
rect 28307 6817 28319 6851
rect 28261 6811 28319 6817
rect 28445 6851 28503 6857
rect 28445 6817 28457 6851
rect 28491 6848 28503 6851
rect 28644 6848 28672 6876
rect 28491 6820 28672 6848
rect 28491 6817 28503 6820
rect 28445 6811 28503 6817
rect 24213 6783 24271 6789
rect 24213 6749 24225 6783
rect 24259 6749 24271 6783
rect 28276 6780 28304 6811
rect 28718 6808 28724 6860
rect 28776 6808 28782 6860
rect 28902 6808 28908 6860
rect 28960 6808 28966 6860
rect 29104 6857 29132 6888
rect 29089 6851 29147 6857
rect 29089 6817 29101 6851
rect 29135 6817 29147 6851
rect 29089 6811 29147 6817
rect 29730 6808 29736 6860
rect 29788 6808 29794 6860
rect 29822 6808 29828 6860
rect 29880 6848 29886 6860
rect 30193 6851 30251 6857
rect 30193 6848 30205 6851
rect 29880 6820 30205 6848
rect 29880 6808 29886 6820
rect 30193 6817 30205 6820
rect 30239 6848 30251 6851
rect 30668 6848 30696 6944
rect 30239 6820 30696 6848
rect 30837 6851 30895 6857
rect 30239 6817 30251 6820
rect 30193 6811 30251 6817
rect 30837 6817 30849 6851
rect 30883 6817 30895 6851
rect 30837 6811 30895 6817
rect 28920 6780 28948 6808
rect 30852 6780 30880 6811
rect 28276 6752 28580 6780
rect 28920 6752 30880 6780
rect 24213 6743 24271 6749
rect 22646 6644 22652 6656
rect 21836 6616 22652 6644
rect 22646 6604 22652 6616
rect 22704 6604 22710 6656
rect 22830 6604 22836 6656
rect 22888 6604 22894 6656
rect 22922 6604 22928 6656
rect 22980 6644 22986 6656
rect 24228 6644 24256 6743
rect 28552 6721 28580 6752
rect 28537 6715 28595 6721
rect 28537 6681 28549 6715
rect 28583 6712 28595 6715
rect 28583 6684 30972 6712
rect 28583 6681 28595 6684
rect 28537 6675 28595 6681
rect 30944 6656 30972 6684
rect 22980 6616 24256 6644
rect 26145 6647 26203 6653
rect 22980 6604 22986 6616
rect 26145 6613 26157 6647
rect 26191 6644 26203 6647
rect 27154 6644 27160 6656
rect 26191 6616 27160 6644
rect 26191 6613 26203 6616
rect 26145 6607 26203 6613
rect 27154 6604 27160 6616
rect 27212 6604 27218 6656
rect 28166 6604 28172 6656
rect 28224 6604 28230 6656
rect 28810 6604 28816 6656
rect 28868 6604 28874 6656
rect 29273 6647 29331 6653
rect 29273 6613 29285 6647
rect 29319 6644 29331 6647
rect 29730 6644 29736 6656
rect 29319 6616 29736 6644
rect 29319 6613 29331 6616
rect 29273 6607 29331 6613
rect 29730 6604 29736 6616
rect 29788 6604 29794 6656
rect 30650 6604 30656 6656
rect 30708 6604 30714 6656
rect 30926 6604 30932 6656
rect 30984 6604 30990 6656
rect 552 6554 31372 6576
rect 552 6502 4250 6554
rect 4302 6502 4314 6554
rect 4366 6502 4378 6554
rect 4430 6502 4442 6554
rect 4494 6502 4506 6554
rect 4558 6502 11955 6554
rect 12007 6502 12019 6554
rect 12071 6502 12083 6554
rect 12135 6502 12147 6554
rect 12199 6502 12211 6554
rect 12263 6502 19660 6554
rect 19712 6502 19724 6554
rect 19776 6502 19788 6554
rect 19840 6502 19852 6554
rect 19904 6502 19916 6554
rect 19968 6502 27365 6554
rect 27417 6502 27429 6554
rect 27481 6502 27493 6554
rect 27545 6502 27557 6554
rect 27609 6502 27621 6554
rect 27673 6502 31372 6554
rect 552 6480 31372 6502
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6181 6443 6239 6449
rect 6181 6440 6193 6443
rect 6052 6412 6193 6440
rect 6052 6400 6058 6412
rect 6181 6409 6193 6412
rect 6227 6409 6239 6443
rect 6181 6403 6239 6409
rect 2501 6375 2559 6381
rect 2501 6341 2513 6375
rect 2547 6372 2559 6375
rect 2547 6344 2774 6372
rect 2547 6341 2559 6344
rect 2501 6335 2559 6341
rect 937 6239 995 6245
rect 937 6205 949 6239
rect 983 6205 995 6239
rect 937 6199 995 6205
rect 952 6100 980 6199
rect 1026 6196 1032 6248
rect 1084 6236 1090 6248
rect 1193 6239 1251 6245
rect 1193 6236 1205 6239
rect 1084 6208 1205 6236
rect 1084 6196 1090 6208
rect 1193 6205 1205 6208
rect 1239 6205 1251 6239
rect 1193 6199 1251 6205
rect 2590 6196 2596 6248
rect 2648 6196 2654 6248
rect 2746 6236 2774 6344
rect 2958 6264 2964 6316
rect 3016 6304 3022 6316
rect 6196 6304 6224 6403
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6328 6412 6561 6440
rect 6328 6400 6334 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 6840 6412 8432 6440
rect 6840 6381 6868 6412
rect 6825 6375 6883 6381
rect 6825 6341 6837 6375
rect 6871 6341 6883 6375
rect 8404 6372 8432 6412
rect 8478 6400 8484 6452
rect 8536 6400 8542 6452
rect 9585 6443 9643 6449
rect 9585 6409 9597 6443
rect 9631 6440 9643 6443
rect 9766 6440 9772 6452
rect 9631 6412 9772 6440
rect 9631 6409 9643 6412
rect 9585 6403 9643 6409
rect 9766 6400 9772 6412
rect 9824 6440 9830 6452
rect 10502 6440 10508 6452
rect 9824 6412 10508 6440
rect 9824 6400 9830 6412
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 10980 6412 11928 6440
rect 10980 6372 11008 6412
rect 8404 6344 11008 6372
rect 11900 6372 11928 6412
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 12897 6443 12955 6449
rect 12897 6440 12909 6443
rect 12768 6412 12909 6440
rect 12768 6400 12774 6412
rect 12897 6409 12909 6412
rect 12943 6409 12955 6443
rect 12897 6403 12955 6409
rect 13081 6443 13139 6449
rect 13081 6409 13093 6443
rect 13127 6440 13139 6443
rect 13354 6440 13360 6452
rect 13127 6412 13360 6440
rect 13127 6409 13139 6412
rect 13081 6403 13139 6409
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 13998 6400 14004 6452
rect 14056 6400 14062 6452
rect 14277 6443 14335 6449
rect 14277 6409 14289 6443
rect 14323 6440 14335 6443
rect 14366 6440 14372 6452
rect 14323 6412 14372 6440
rect 14323 6409 14335 6412
rect 14277 6403 14335 6409
rect 14366 6400 14372 6412
rect 14424 6400 14430 6452
rect 14458 6400 14464 6452
rect 14516 6400 14522 6452
rect 14553 6443 14611 6449
rect 14553 6409 14565 6443
rect 14599 6440 14611 6443
rect 14826 6440 14832 6452
rect 14599 6412 14832 6440
rect 14599 6409 14611 6412
rect 14553 6403 14611 6409
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 15344 6412 19441 6440
rect 15344 6400 15350 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 21450 6440 21456 6452
rect 19429 6403 19487 6409
rect 19904 6412 21456 6440
rect 14476 6372 14504 6400
rect 14737 6375 14795 6381
rect 14737 6372 14749 6375
rect 11900 6344 13768 6372
rect 14476 6344 14749 6372
rect 6825 6335 6883 6341
rect 8205 6307 8263 6313
rect 3016 6276 3740 6304
rect 3016 6264 3022 6276
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2746 6208 2881 6236
rect 2869 6205 2881 6208
rect 2915 6236 2927 6239
rect 3050 6236 3056 6248
rect 2915 6208 3056 6236
rect 2915 6205 2927 6208
rect 2869 6199 2927 6205
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 3602 6196 3608 6248
rect 3660 6196 3666 6248
rect 3712 6245 3740 6276
rect 4356 6276 4568 6304
rect 6196 6276 6500 6304
rect 4356 6245 4384 6276
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 4341 6239 4399 6245
rect 4341 6236 4353 6239
rect 4111 6208 4353 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4341 6205 4353 6208
rect 4387 6205 4399 6239
rect 4341 6199 4399 6205
rect 3620 6168 3648 6196
rect 2332 6140 3648 6168
rect 3712 6168 3740 6199
rect 4430 6196 4436 6248
rect 4488 6196 4494 6248
rect 4540 6236 4568 6276
rect 5074 6236 5080 6248
rect 4540 6208 5080 6236
rect 5074 6196 5080 6208
rect 5132 6196 5138 6248
rect 6472 6245 6500 6276
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8754 6304 8760 6316
rect 8251 6276 8760 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8754 6264 8760 6276
rect 8812 6304 8818 6316
rect 10594 6304 10600 6316
rect 8812 6276 10600 6304
rect 8812 6264 8818 6276
rect 10594 6264 10600 6276
rect 10652 6304 10658 6316
rect 10962 6304 10968 6316
rect 10652 6276 10968 6304
rect 10652 6264 10658 6276
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 6273 6239 6331 6245
rect 6273 6205 6285 6239
rect 6319 6205 6331 6239
rect 6273 6199 6331 6205
rect 6457 6239 6515 6245
rect 6457 6205 6469 6239
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 4678 6171 4736 6177
rect 4678 6168 4690 6171
rect 3712 6140 4690 6168
rect 2332 6109 2360 6140
rect 4678 6137 4690 6140
rect 4724 6168 4736 6171
rect 4890 6168 4896 6180
rect 4724 6140 4896 6168
rect 4724 6137 4736 6140
rect 4678 6131 4736 6137
rect 4890 6128 4896 6140
rect 4948 6128 4954 6180
rect 6288 6168 6316 6199
rect 6546 6196 6552 6248
rect 6604 6196 6610 6248
rect 7949 6239 8007 6245
rect 7949 6205 7961 6239
rect 7995 6236 8007 6239
rect 8389 6239 8447 6245
rect 8389 6236 8401 6239
rect 7995 6208 8401 6236
rect 7995 6205 8007 6208
rect 7949 6199 8007 6205
rect 8389 6205 8401 6208
rect 8435 6236 8447 6239
rect 8665 6239 8723 6245
rect 8665 6236 8677 6239
rect 8435 6208 8677 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 8665 6205 8677 6208
rect 8711 6236 8723 6239
rect 8846 6236 8852 6248
rect 8711 6208 8852 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 8846 6196 8852 6208
rect 8904 6196 8910 6248
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 9217 6239 9275 6245
rect 9217 6236 9229 6239
rect 8996 6208 9229 6236
rect 8996 6196 9002 6208
rect 9217 6205 9229 6208
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6205 9551 6239
rect 9493 6199 9551 6205
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6236 10011 6239
rect 10137 6239 10195 6245
rect 10137 6236 10149 6239
rect 9999 6208 10149 6236
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 10137 6205 10149 6208
rect 10183 6236 10195 6239
rect 10318 6236 10324 6248
rect 10183 6208 10324 6236
rect 10183 6205 10195 6208
rect 10137 6199 10195 6205
rect 6564 6168 6592 6196
rect 6288 6140 6592 6168
rect 8757 6171 8815 6177
rect 8757 6137 8769 6171
rect 8803 6168 8815 6171
rect 9508 6168 9536 6199
rect 9674 6168 9680 6180
rect 8803 6140 9680 6168
rect 8803 6137 8815 6140
rect 8757 6131 8815 6137
rect 9674 6128 9680 6140
rect 9732 6168 9738 6180
rect 9861 6171 9919 6177
rect 9861 6168 9873 6171
rect 9732 6140 9873 6168
rect 9732 6128 9738 6140
rect 9861 6137 9873 6140
rect 9907 6137 9919 6171
rect 9861 6131 9919 6137
rect 492 6072 980 6100
rect 2317 6103 2375 6109
rect 492 5828 520 6072
rect 2317 6069 2329 6103
rect 2363 6069 2375 6103
rect 2317 6063 2375 6069
rect 2406 6060 2412 6112
rect 2464 6100 2470 6112
rect 2777 6103 2835 6109
rect 2777 6100 2789 6103
rect 2464 6072 2789 6100
rect 2464 6060 2470 6072
rect 2777 6069 2789 6072
rect 2823 6069 2835 6103
rect 2777 6063 2835 6069
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3200 6072 3617 6100
rect 3200 6060 3206 6072
rect 3605 6069 3617 6072
rect 3651 6100 3663 6103
rect 3973 6103 4031 6109
rect 3973 6100 3985 6103
rect 3651 6072 3985 6100
rect 3651 6069 3663 6072
rect 3605 6063 3663 6069
rect 3973 6069 3985 6072
rect 4019 6069 4031 6103
rect 3973 6063 4031 6069
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 4212 6072 4261 6100
rect 4212 6060 4218 6072
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 4249 6063 4307 6069
rect 5813 6103 5871 6109
rect 5813 6069 5825 6103
rect 5859 6100 5871 6103
rect 8938 6100 8944 6112
rect 5859 6072 8944 6100
rect 5859 6069 5871 6072
rect 5813 6063 5871 6069
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 9030 6060 9036 6112
rect 9088 6060 9094 6112
rect 9309 6103 9367 6109
rect 9309 6069 9321 6103
rect 9355 6100 9367 6103
rect 9968 6100 9996 6199
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 10410 6196 10416 6248
rect 10468 6236 10474 6248
rect 10468 6208 10548 6236
rect 10468 6196 10474 6208
rect 10229 6171 10287 6177
rect 10229 6137 10241 6171
rect 10275 6168 10287 6171
rect 10520 6168 10548 6208
rect 10686 6196 10692 6248
rect 10744 6196 10750 6248
rect 11606 6196 11612 6248
rect 11664 6236 11670 6248
rect 11664 6211 12956 6236
rect 11664 6208 13001 6211
rect 11664 6196 11670 6208
rect 12928 6205 13001 6208
rect 10781 6171 10839 6177
rect 10781 6168 10793 6171
rect 10275 6140 10793 6168
rect 10275 6137 10287 6140
rect 10229 6131 10287 6137
rect 10781 6137 10793 6140
rect 10827 6137 10839 6171
rect 11210 6171 11268 6177
rect 11210 6168 11222 6171
rect 10781 6131 10839 6137
rect 10888 6140 11222 6168
rect 9355 6072 9996 6100
rect 9355 6069 9367 6072
rect 9309 6063 9367 6069
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 10888 6100 10916 6140
rect 11210 6137 11222 6140
rect 11256 6137 11268 6171
rect 11210 6131 11268 6137
rect 12710 6128 12716 6180
rect 12768 6128 12774 6180
rect 12928 6171 12955 6205
rect 12989 6171 13001 6205
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13740 6245 13768 6344
rect 14737 6341 14749 6344
rect 14783 6341 14795 6375
rect 14737 6335 14795 6341
rect 15930 6332 15936 6384
rect 15988 6332 15994 6384
rect 16114 6332 16120 6384
rect 16172 6372 16178 6384
rect 16850 6372 16856 6384
rect 16172 6344 16856 6372
rect 16172 6332 16178 6344
rect 16850 6332 16856 6344
rect 16908 6372 16914 6384
rect 19061 6375 19119 6381
rect 19061 6372 19073 6375
rect 16908 6344 19073 6372
rect 16908 6332 16914 6344
rect 19061 6341 19073 6344
rect 19107 6372 19119 6375
rect 19904 6372 19932 6412
rect 21450 6400 21456 6412
rect 21508 6400 21514 6452
rect 22094 6400 22100 6452
rect 22152 6400 22158 6452
rect 22278 6400 22284 6452
rect 22336 6440 22342 6452
rect 22925 6443 22983 6449
rect 22925 6440 22937 6443
rect 22336 6412 22937 6440
rect 22336 6400 22342 6412
rect 19107 6344 19932 6372
rect 19107 6341 19119 6344
rect 19061 6335 19119 6341
rect 15657 6307 15715 6313
rect 15657 6304 15669 6307
rect 14936 6276 15669 6304
rect 14936 6248 14964 6276
rect 15657 6273 15669 6276
rect 15703 6273 15715 6307
rect 15657 6267 15715 6273
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6304 15807 6307
rect 17862 6304 17868 6316
rect 15795 6276 17448 6304
rect 15795 6273 15807 6276
rect 15749 6267 15807 6273
rect 13541 6239 13599 6245
rect 13541 6236 13553 6239
rect 13412 6208 13553 6236
rect 13412 6196 13418 6208
rect 13541 6205 13553 6208
rect 13587 6205 13599 6239
rect 13541 6199 13599 6205
rect 13725 6239 13783 6245
rect 13725 6205 13737 6239
rect 13771 6205 13783 6239
rect 13725 6199 13783 6205
rect 13814 6196 13820 6248
rect 13872 6196 13878 6248
rect 13906 6196 13912 6248
rect 13964 6196 13970 6248
rect 14918 6196 14924 6248
rect 14976 6196 14982 6248
rect 15194 6196 15200 6248
rect 15252 6196 15258 6248
rect 15562 6245 15568 6248
rect 15547 6239 15568 6245
rect 15547 6205 15559 6239
rect 15620 6238 15626 6248
rect 15547 6199 15568 6205
rect 15562 6196 15568 6199
rect 15620 6196 15634 6238
rect 15672 6236 15700 6267
rect 17420 6245 17448 6276
rect 17696 6276 17868 6304
rect 17696 6245 17724 6276
rect 17862 6264 17868 6276
rect 17920 6304 17926 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 17920 6276 18705 6304
rect 17920 6264 17926 6276
rect 18693 6273 18705 6276
rect 18739 6304 18751 6307
rect 18782 6304 18788 6316
rect 18739 6276 18788 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 19334 6264 19340 6316
rect 19392 6264 19398 6316
rect 20732 6276 22048 6304
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 15672 6208 17325 6236
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 17405 6239 17463 6245
rect 17405 6205 17417 6239
rect 17451 6236 17463 6239
rect 17681 6239 17739 6245
rect 17451 6208 17540 6236
rect 17451 6205 17463 6208
rect 17405 6199 17463 6205
rect 12928 6168 13001 6171
rect 12928 6140 13768 6168
rect 10376 6072 10916 6100
rect 12345 6103 12403 6109
rect 10376 6060 10382 6072
rect 12345 6069 12357 6103
rect 12391 6100 12403 6103
rect 13630 6100 13636 6112
rect 12391 6072 13636 6100
rect 12391 6069 12403 6072
rect 12345 6063 12403 6069
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 13740 6100 13768 6140
rect 14366 6128 14372 6180
rect 14424 6128 14430 6180
rect 14585 6171 14643 6177
rect 14585 6137 14597 6171
rect 14631 6168 14643 6171
rect 15212 6168 15240 6196
rect 14631 6140 15240 6168
rect 15606 6168 15634 6196
rect 17512 6180 17540 6208
rect 17681 6205 17693 6239
rect 17727 6205 17739 6239
rect 17957 6239 18015 6245
rect 17957 6236 17969 6239
rect 17681 6199 17739 6205
rect 17788 6208 17969 6236
rect 17788 6180 17816 6208
rect 17957 6205 17969 6208
rect 18003 6205 18015 6239
rect 17957 6199 18015 6205
rect 18101 6239 18159 6245
rect 18101 6205 18113 6239
rect 18147 6236 18159 6239
rect 18506 6236 18512 6248
rect 18147 6208 18512 6236
rect 18147 6205 18159 6208
rect 18101 6199 18159 6205
rect 18506 6196 18512 6208
rect 18564 6196 18570 6248
rect 18874 6196 18880 6248
rect 18932 6196 18938 6248
rect 19352 6236 19380 6264
rect 20162 6236 20168 6248
rect 19352 6208 20168 6236
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 20553 6239 20611 6245
rect 20553 6205 20565 6239
rect 20599 6236 20611 6239
rect 20732 6236 20760 6276
rect 20599 6208 20760 6236
rect 20599 6205 20611 6208
rect 20553 6199 20611 6205
rect 20806 6196 20812 6248
rect 20864 6236 20870 6248
rect 21358 6236 21364 6248
rect 20864 6208 21364 6236
rect 20864 6196 20870 6208
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 21910 6196 21916 6248
rect 21968 6196 21974 6248
rect 22020 6245 22048 6276
rect 22005 6239 22063 6245
rect 22005 6205 22017 6239
rect 22051 6205 22063 6239
rect 22112 6236 22140 6400
rect 22646 6332 22652 6384
rect 22704 6332 22710 6384
rect 22756 6245 22784 6412
rect 22925 6409 22937 6412
rect 22971 6440 22983 6443
rect 23201 6443 23259 6449
rect 23201 6440 23213 6443
rect 22971 6412 23213 6440
rect 22971 6409 22983 6412
rect 22925 6403 22983 6409
rect 23201 6409 23213 6412
rect 23247 6409 23259 6443
rect 23201 6403 23259 6409
rect 23477 6443 23535 6449
rect 23477 6409 23489 6443
rect 23523 6440 23535 6443
rect 24210 6440 24216 6452
rect 23523 6412 24216 6440
rect 23523 6409 23535 6412
rect 23477 6403 23535 6409
rect 24210 6400 24216 6412
rect 24268 6400 24274 6452
rect 28626 6400 28632 6452
rect 28684 6440 28690 6452
rect 28721 6443 28779 6449
rect 28721 6440 28733 6443
rect 28684 6412 28733 6440
rect 28684 6400 28690 6412
rect 28721 6409 28733 6412
rect 28767 6409 28779 6443
rect 28721 6403 28779 6409
rect 31018 6400 31024 6452
rect 31076 6400 31082 6452
rect 24489 6375 24547 6381
rect 24489 6372 24501 6375
rect 22848 6344 24501 6372
rect 22848 6245 22876 6344
rect 24489 6341 24501 6344
rect 24535 6372 24547 6375
rect 24765 6375 24823 6381
rect 24765 6372 24777 6375
rect 24535 6344 24777 6372
rect 24535 6341 24547 6344
rect 24489 6335 24547 6341
rect 24765 6341 24777 6344
rect 24811 6341 24823 6375
rect 24765 6335 24823 6341
rect 26234 6332 26240 6384
rect 26292 6372 26298 6384
rect 27801 6375 27859 6381
rect 27801 6372 27813 6375
rect 26292 6344 27813 6372
rect 26292 6332 26298 6344
rect 27801 6341 27813 6344
rect 27847 6372 27859 6375
rect 28077 6375 28135 6381
rect 28077 6372 28089 6375
rect 27847 6344 28089 6372
rect 27847 6341 27859 6344
rect 27801 6335 27859 6341
rect 28077 6341 28089 6344
rect 28123 6341 28135 6375
rect 28077 6335 28135 6341
rect 28810 6332 28816 6384
rect 28868 6332 28874 6384
rect 23934 6304 23940 6316
rect 23308 6276 23940 6304
rect 23308 6245 23336 6276
rect 23934 6264 23940 6276
rect 23992 6304 23998 6316
rect 26421 6307 26479 6313
rect 26421 6304 26433 6307
rect 23992 6276 25084 6304
rect 23992 6264 23998 6276
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 22112 6208 22477 6236
rect 22005 6199 22063 6205
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 22465 6199 22523 6205
rect 22741 6239 22799 6245
rect 22741 6205 22753 6239
rect 22787 6205 22799 6239
rect 22741 6199 22799 6205
rect 22833 6239 22891 6245
rect 22833 6205 22845 6239
rect 22879 6205 22891 6239
rect 22833 6199 22891 6205
rect 23293 6239 23351 6245
rect 23293 6205 23305 6239
rect 23339 6205 23351 6239
rect 23293 6199 23351 6205
rect 23569 6239 23627 6245
rect 23569 6205 23581 6239
rect 23615 6236 23627 6239
rect 23750 6236 23756 6248
rect 23615 6208 23756 6236
rect 23615 6205 23627 6208
rect 23569 6199 23627 6205
rect 16850 6168 16856 6180
rect 15606 6140 16856 6168
rect 14631 6137 14643 6140
rect 14585 6131 14643 6137
rect 14600 6100 14628 6131
rect 16850 6128 16856 6140
rect 16908 6168 16914 6180
rect 17129 6171 17187 6177
rect 17129 6168 17141 6171
rect 16908 6140 17141 6168
rect 16908 6128 16914 6140
rect 17129 6137 17141 6140
rect 17175 6137 17187 6171
rect 17129 6131 17187 6137
rect 17494 6128 17500 6180
rect 17552 6128 17558 6180
rect 17770 6128 17776 6180
rect 17828 6128 17834 6180
rect 17865 6171 17923 6177
rect 17865 6137 17877 6171
rect 17911 6137 17923 6171
rect 17865 6131 17923 6137
rect 13740 6072 14628 6100
rect 17405 6103 17463 6109
rect 17405 6069 17417 6103
rect 17451 6100 17463 6103
rect 17880 6100 17908 6131
rect 21174 6128 21180 6180
rect 21232 6128 21238 6180
rect 18138 6100 18144 6112
rect 17451 6072 18144 6100
rect 17451 6069 17463 6072
rect 17405 6063 17463 6069
rect 18138 6060 18144 6072
rect 18196 6060 18202 6112
rect 18250 6103 18308 6109
rect 18250 6069 18262 6103
rect 18296 6100 18308 6103
rect 19518 6100 19524 6112
rect 18296 6072 19524 6100
rect 18296 6069 18308 6072
rect 18250 6063 18308 6069
rect 19518 6060 19524 6072
rect 19576 6060 19582 6112
rect 22020 6100 22048 6199
rect 22848 6168 22876 6199
rect 23750 6196 23756 6208
rect 23808 6196 23814 6248
rect 24029 6239 24087 6245
rect 24029 6205 24041 6239
rect 24075 6236 24087 6239
rect 24210 6236 24216 6248
rect 24075 6208 24216 6236
rect 24075 6205 24087 6208
rect 24029 6199 24087 6205
rect 24210 6196 24216 6208
rect 24268 6196 24274 6248
rect 24320 6245 24348 6276
rect 24305 6239 24363 6245
rect 24305 6205 24317 6239
rect 24351 6205 24363 6239
rect 24305 6199 24363 6205
rect 24397 6239 24455 6245
rect 24397 6205 24409 6239
rect 24443 6205 24455 6239
rect 24857 6239 24915 6245
rect 24857 6236 24869 6239
rect 24397 6199 24455 6205
rect 24504 6208 24869 6236
rect 22296 6140 22876 6168
rect 24228 6168 24256 6196
rect 24412 6168 24440 6199
rect 24228 6140 24440 6168
rect 22296 6100 22324 6140
rect 24504 6112 24532 6208
rect 24857 6205 24869 6208
rect 24903 6236 24915 6239
rect 24949 6239 25007 6245
rect 24949 6236 24961 6239
rect 24903 6208 24961 6236
rect 24903 6205 24915 6208
rect 24857 6199 24915 6205
rect 24949 6205 24961 6208
rect 24995 6205 25007 6239
rect 24949 6199 25007 6205
rect 22020 6072 22324 6100
rect 22370 6060 22376 6112
rect 22428 6060 22434 6112
rect 22646 6060 22652 6112
rect 22704 6100 22710 6112
rect 23937 6103 23995 6109
rect 23937 6100 23949 6103
rect 22704 6072 23949 6100
rect 22704 6060 22710 6072
rect 23937 6069 23949 6072
rect 23983 6069 23995 6103
rect 23937 6063 23995 6069
rect 24486 6060 24492 6112
rect 24544 6060 24550 6112
rect 24872 6100 24900 6199
rect 25056 6177 25084 6276
rect 25976 6276 26433 6304
rect 25130 6196 25136 6248
rect 25188 6236 25194 6248
rect 25409 6239 25467 6245
rect 25409 6236 25421 6239
rect 25188 6208 25421 6236
rect 25188 6196 25194 6208
rect 25409 6205 25421 6208
rect 25455 6205 25467 6239
rect 25409 6199 25467 6205
rect 25685 6239 25743 6245
rect 25685 6205 25697 6239
rect 25731 6236 25743 6239
rect 25774 6236 25780 6248
rect 25731 6208 25780 6236
rect 25731 6205 25743 6208
rect 25685 6199 25743 6205
rect 25041 6171 25099 6177
rect 25041 6137 25053 6171
rect 25087 6168 25099 6171
rect 25317 6171 25375 6177
rect 25317 6168 25329 6171
rect 25087 6140 25329 6168
rect 25087 6137 25099 6140
rect 25041 6131 25099 6137
rect 25317 6137 25329 6140
rect 25363 6137 25375 6171
rect 25424 6168 25452 6199
rect 25774 6196 25780 6208
rect 25832 6236 25838 6248
rect 25976 6245 26004 6276
rect 26421 6273 26433 6276
rect 26467 6304 26479 6307
rect 26697 6307 26755 6313
rect 26697 6304 26709 6307
rect 26467 6276 26709 6304
rect 26467 6273 26479 6276
rect 26421 6267 26479 6273
rect 26697 6273 26709 6276
rect 26743 6273 26755 6307
rect 28534 6304 28540 6316
rect 26697 6267 26755 6273
rect 28276 6276 28540 6304
rect 25961 6239 26019 6245
rect 25961 6236 25973 6239
rect 25832 6208 25973 6236
rect 25832 6196 25838 6208
rect 25961 6205 25973 6208
rect 26007 6205 26019 6239
rect 25961 6199 26019 6205
rect 26050 6196 26056 6248
rect 26108 6236 26114 6248
rect 26237 6239 26295 6245
rect 26237 6236 26249 6239
rect 26108 6208 26249 6236
rect 26108 6196 26114 6208
rect 26237 6205 26249 6208
rect 26283 6205 26295 6239
rect 26237 6199 26295 6205
rect 25869 6171 25927 6177
rect 25869 6168 25881 6171
rect 25424 6140 25881 6168
rect 25317 6131 25375 6137
rect 25869 6137 25881 6140
rect 25915 6168 25927 6171
rect 26145 6171 26203 6177
rect 26145 6168 26157 6171
rect 25915 6140 26157 6168
rect 25915 6137 25927 6140
rect 25869 6131 25927 6137
rect 26145 6137 26157 6140
rect 26191 6137 26203 6171
rect 26252 6168 26280 6199
rect 26326 6196 26332 6248
rect 26384 6196 26390 6248
rect 26789 6239 26847 6245
rect 26789 6205 26801 6239
rect 26835 6236 26847 6239
rect 27065 6239 27123 6245
rect 27065 6236 27077 6239
rect 26835 6208 27077 6236
rect 26835 6205 26847 6208
rect 26789 6199 26847 6205
rect 27065 6205 27077 6208
rect 27111 6205 27123 6239
rect 27065 6199 27123 6205
rect 26973 6171 27031 6177
rect 26973 6168 26985 6171
rect 26252 6140 26985 6168
rect 26145 6131 26203 6137
rect 26973 6137 26985 6140
rect 27019 6137 27031 6171
rect 27080 6168 27108 6199
rect 27154 6196 27160 6248
rect 27212 6236 27218 6248
rect 27341 6239 27399 6245
rect 27341 6236 27353 6239
rect 27212 6208 27353 6236
rect 27212 6196 27218 6208
rect 27341 6205 27353 6208
rect 27387 6236 27399 6239
rect 27430 6236 27436 6248
rect 27387 6208 27436 6236
rect 27387 6205 27399 6208
rect 27341 6199 27399 6205
rect 27430 6196 27436 6208
rect 27488 6196 27494 6248
rect 27614 6196 27620 6248
rect 27672 6236 27678 6248
rect 27709 6239 27767 6245
rect 27709 6236 27721 6239
rect 27672 6208 27721 6236
rect 27672 6196 27678 6208
rect 27709 6205 27721 6208
rect 27755 6205 27767 6239
rect 27709 6199 27767 6205
rect 28166 6196 28172 6248
rect 28224 6236 28230 6248
rect 28276 6236 28304 6276
rect 28534 6264 28540 6276
rect 28592 6264 28598 6316
rect 28828 6304 28856 6332
rect 29178 6304 29184 6316
rect 28828 6276 29184 6304
rect 29178 6264 29184 6276
rect 29236 6304 29242 6316
rect 29236 6276 29592 6304
rect 29236 6264 29242 6276
rect 28442 6236 28448 6248
rect 28224 6208 28304 6236
rect 28405 6208 28448 6236
rect 28224 6196 28230 6208
rect 28442 6196 28448 6208
rect 28500 6196 28506 6248
rect 29564 6245 29592 6276
rect 28813 6239 28871 6245
rect 28813 6205 28825 6239
rect 28859 6205 28871 6239
rect 28813 6199 28871 6205
rect 29549 6239 29607 6245
rect 29549 6205 29561 6239
rect 29595 6205 29607 6239
rect 29549 6199 29607 6205
rect 27249 6171 27307 6177
rect 27249 6168 27261 6171
rect 27080 6140 27261 6168
rect 26973 6131 27031 6137
rect 27249 6137 27261 6140
rect 27295 6168 27307 6171
rect 27525 6171 27583 6177
rect 27525 6168 27537 6171
rect 27295 6140 27537 6168
rect 27295 6137 27307 6140
rect 27249 6131 27307 6137
rect 27525 6137 27537 6140
rect 27571 6137 27583 6171
rect 28828 6168 28856 6199
rect 29638 6196 29644 6248
rect 29696 6196 29702 6248
rect 29730 6196 29736 6248
rect 29788 6236 29794 6248
rect 29897 6239 29955 6245
rect 29897 6236 29909 6239
rect 29788 6208 29909 6236
rect 29788 6196 29794 6208
rect 29897 6205 29909 6208
rect 29943 6205 29955 6239
rect 29897 6199 29955 6205
rect 30374 6196 30380 6248
rect 30432 6196 30438 6248
rect 30392 6168 30420 6196
rect 28828 6140 30420 6168
rect 27525 6131 27583 6137
rect 25593 6103 25651 6109
rect 25593 6100 25605 6103
rect 24872 6072 25605 6100
rect 25593 6069 25605 6072
rect 25639 6069 25651 6103
rect 25593 6063 25651 6069
rect 27430 6060 27436 6112
rect 27488 6100 27494 6112
rect 28353 6103 28411 6109
rect 28353 6100 28365 6103
rect 27488 6072 28365 6100
rect 27488 6060 27494 6072
rect 28353 6069 28365 6072
rect 28399 6069 28411 6103
rect 28353 6063 28411 6069
rect 29362 6060 29368 6112
rect 29420 6060 29426 6112
rect 552 6010 31531 6032
rect 552 5958 8102 6010
rect 8154 5958 8166 6010
rect 8218 5958 8230 6010
rect 8282 5958 8294 6010
rect 8346 5958 8358 6010
rect 8410 5958 15807 6010
rect 15859 5958 15871 6010
rect 15923 5958 15935 6010
rect 15987 5958 15999 6010
rect 16051 5958 16063 6010
rect 16115 5958 23512 6010
rect 23564 5958 23576 6010
rect 23628 5958 23640 6010
rect 23692 5958 23704 6010
rect 23756 5958 23768 6010
rect 23820 5958 31217 6010
rect 31269 5958 31281 6010
rect 31333 5958 31345 6010
rect 31397 5958 31409 6010
rect 31461 5958 31473 6010
rect 31525 5958 31531 6010
rect 552 5936 31531 5958
rect 1136 5868 1961 5896
rect 1136 5828 1164 5868
rect 492 5800 1164 5828
rect 1933 5828 1961 5868
rect 2590 5856 2596 5908
rect 2648 5896 2654 5908
rect 2777 5899 2835 5905
rect 2777 5896 2789 5899
rect 2648 5868 2789 5896
rect 2648 5856 2654 5868
rect 2777 5865 2789 5868
rect 2823 5865 2835 5899
rect 4430 5896 4436 5908
rect 2777 5859 2835 5865
rect 3344 5868 4436 5896
rect 2682 5828 2688 5840
rect 1933 5800 2688 5828
rect 1136 5769 1164 5800
rect 2682 5788 2688 5800
rect 2740 5828 2746 5840
rect 3344 5828 3372 5868
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 4614 5856 4620 5908
rect 4672 5856 4678 5908
rect 4890 5856 4896 5908
rect 4948 5856 4954 5908
rect 7193 5899 7251 5905
rect 7193 5865 7205 5899
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 2740 5800 3372 5828
rect 2740 5788 2746 5800
rect 1394 5769 1400 5772
rect 1029 5763 1087 5769
rect 1029 5760 1041 5763
rect 860 5732 1041 5760
rect 860 5556 888 5732
rect 1029 5729 1041 5732
rect 1075 5729 1087 5763
rect 1029 5723 1087 5729
rect 1121 5763 1179 5769
rect 1121 5729 1133 5763
rect 1167 5729 1179 5763
rect 1377 5763 1400 5769
rect 1377 5760 1389 5763
rect 1121 5723 1179 5729
rect 1228 5732 1389 5760
rect 937 5695 995 5701
rect 937 5661 949 5695
rect 983 5692 995 5695
rect 1228 5692 1256 5732
rect 1377 5729 1389 5732
rect 1377 5723 1400 5729
rect 1394 5720 1400 5723
rect 1452 5720 1458 5772
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5760 2927 5763
rect 2958 5760 2964 5772
rect 2915 5732 2964 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 3142 5720 3148 5772
rect 3200 5720 3206 5772
rect 3252 5769 3280 5800
rect 4154 5788 4160 5840
rect 4212 5828 4218 5840
rect 5169 5831 5227 5837
rect 5169 5828 5181 5831
rect 4212 5800 5181 5828
rect 4212 5788 4218 5800
rect 5169 5797 5181 5800
rect 5215 5797 5227 5831
rect 7208 5828 7236 5859
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 9582 5896 9588 5908
rect 8996 5868 9588 5896
rect 8996 5856 9002 5868
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 10318 5856 10324 5908
rect 10376 5856 10382 5908
rect 12342 5896 12348 5908
rect 12084 5868 12348 5896
rect 11606 5828 11612 5840
rect 7208 5800 11612 5828
rect 5169 5791 5227 5797
rect 11606 5788 11612 5800
rect 11664 5788 11670 5840
rect 12084 5837 12112 5868
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 12710 5856 12716 5908
rect 12768 5856 12774 5908
rect 14185 5899 14243 5905
rect 14185 5865 14197 5899
rect 14231 5896 14243 5899
rect 14274 5896 14280 5908
rect 14231 5868 14280 5896
rect 14231 5865 14243 5868
rect 14185 5859 14243 5865
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 15102 5856 15108 5908
rect 15160 5896 15166 5908
rect 19061 5899 19119 5905
rect 19061 5896 19073 5899
rect 15160 5868 19073 5896
rect 15160 5856 15166 5868
rect 19061 5865 19073 5868
rect 19107 5865 19119 5899
rect 19679 5899 19737 5905
rect 19679 5896 19691 5899
rect 19061 5859 19119 5865
rect 19168 5868 19691 5896
rect 12069 5831 12127 5837
rect 12069 5797 12081 5831
rect 12115 5797 12127 5831
rect 12728 5828 12756 5856
rect 12069 5791 12127 5797
rect 12176 5800 12756 5828
rect 3510 5769 3516 5772
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5729 3295 5763
rect 3504 5760 3516 5769
rect 3471 5732 3516 5760
rect 3237 5723 3295 5729
rect 3504 5723 3516 5732
rect 3510 5720 3516 5723
rect 3568 5720 3574 5772
rect 4982 5720 4988 5772
rect 5040 5720 5046 5772
rect 5074 5720 5080 5772
rect 5132 5720 5138 5772
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 5442 5760 5448 5772
rect 5307 5732 5448 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 5718 5720 5724 5772
rect 5776 5760 5782 5772
rect 5813 5763 5871 5769
rect 5813 5760 5825 5763
rect 5776 5732 5825 5760
rect 5776 5720 5782 5732
rect 5813 5729 5825 5732
rect 5859 5729 5871 5763
rect 6069 5763 6127 5769
rect 6069 5760 6081 5763
rect 5813 5723 5871 5729
rect 5920 5732 6081 5760
rect 983 5664 1256 5692
rect 5092 5692 5120 5720
rect 5920 5692 5948 5732
rect 6069 5729 6081 5732
rect 6115 5729 6127 5763
rect 6069 5723 6127 5729
rect 7469 5763 7527 5769
rect 7469 5729 7481 5763
rect 7515 5760 7527 5763
rect 7742 5760 7748 5772
rect 7515 5732 7748 5760
rect 7515 5729 7527 5732
rect 7469 5723 7527 5729
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 8202 5760 8208 5772
rect 7883 5732 8208 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 9674 5720 9680 5772
rect 9732 5720 9738 5772
rect 9950 5720 9956 5772
rect 10008 5720 10014 5772
rect 10410 5720 10416 5772
rect 10468 5720 10474 5772
rect 12176 5760 12204 5800
rect 14090 5788 14096 5840
rect 14148 5828 14154 5840
rect 15013 5831 15071 5837
rect 15013 5828 15025 5831
rect 14148 5800 15025 5828
rect 14148 5788 14154 5800
rect 15013 5797 15025 5800
rect 15059 5797 15071 5831
rect 18049 5831 18107 5837
rect 18049 5828 18061 5831
rect 15013 5791 15071 5797
rect 16868 5800 18061 5828
rect 16868 5772 16896 5800
rect 18049 5797 18061 5800
rect 18095 5797 18107 5831
rect 19168 5828 19196 5868
rect 19679 5865 19691 5868
rect 19725 5896 19737 5899
rect 19978 5896 19984 5908
rect 19725 5868 19984 5896
rect 19725 5865 19737 5868
rect 19679 5859 19737 5865
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 20149 5899 20207 5905
rect 20149 5896 20161 5899
rect 20088 5868 20161 5896
rect 19242 5837 19248 5840
rect 18049 5791 18107 5797
rect 19076 5800 19196 5828
rect 19229 5831 19248 5837
rect 10520 5732 12204 5760
rect 10520 5692 10548 5732
rect 12250 5720 12256 5772
rect 12308 5760 12314 5772
rect 12417 5763 12475 5769
rect 12417 5760 12429 5763
rect 12308 5732 12429 5760
rect 12308 5720 12314 5732
rect 12417 5729 12429 5732
rect 12463 5729 12475 5763
rect 12417 5723 12475 5729
rect 14918 5720 14924 5772
rect 14976 5720 14982 5772
rect 15105 5763 15163 5769
rect 15105 5729 15117 5763
rect 15151 5760 15163 5763
rect 15562 5760 15568 5772
rect 15151 5732 15568 5760
rect 15151 5729 15163 5732
rect 15105 5723 15163 5729
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 16482 5760 16488 5772
rect 16408 5732 16488 5760
rect 5092 5664 5948 5692
rect 7576 5664 10548 5692
rect 983 5661 995 5664
rect 937 5655 995 5661
rect 2406 5584 2412 5636
rect 2464 5584 2470 5636
rect 2501 5627 2559 5633
rect 2501 5593 2513 5627
rect 2547 5624 2559 5627
rect 7576 5624 7604 5664
rect 10686 5652 10692 5704
rect 10744 5652 10750 5704
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5692 11391 5695
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 11379 5664 12173 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 14936 5692 14964 5720
rect 16408 5692 16436 5732
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 16850 5720 16856 5772
rect 16908 5720 16914 5772
rect 16942 5720 16948 5772
rect 17000 5720 17006 5772
rect 17221 5763 17279 5769
rect 17221 5729 17233 5763
rect 17267 5729 17279 5763
rect 17221 5723 17279 5729
rect 14936 5664 16436 5692
rect 12161 5655 12219 5661
rect 2547 5596 3280 5624
rect 2547 5593 2559 5596
rect 2501 5587 2559 5593
rect 2424 5556 2452 5584
rect 860 5528 2452 5556
rect 3050 5516 3056 5568
rect 3108 5516 3114 5568
rect 3252 5556 3280 5596
rect 6748 5596 7604 5624
rect 6748 5556 6776 5596
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 9861 5627 9919 5633
rect 9861 5624 9873 5627
rect 9548 5596 9873 5624
rect 9548 5584 9554 5596
rect 9861 5593 9873 5596
rect 9907 5593 9919 5627
rect 9861 5587 9919 5593
rect 3252 5528 6776 5556
rect 7282 5516 7288 5568
rect 7340 5556 7346 5568
rect 7377 5559 7435 5565
rect 7377 5556 7389 5559
rect 7340 5528 7389 5556
rect 7340 5516 7346 5528
rect 7377 5525 7389 5528
rect 7423 5556 7435 5559
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 7423 5528 7757 5556
rect 7423 5525 7435 5528
rect 7377 5519 7435 5525
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 7745 5519 7803 5525
rect 9030 5516 9036 5568
rect 9088 5556 9094 5568
rect 9306 5556 9312 5568
rect 9088 5528 9312 5556
rect 9088 5516 9094 5528
rect 9306 5516 9312 5528
rect 9364 5556 9370 5568
rect 9585 5559 9643 5565
rect 9585 5556 9597 5559
rect 9364 5528 9597 5556
rect 9364 5516 9370 5528
rect 9585 5525 9597 5528
rect 9631 5556 9643 5559
rect 10704 5556 10732 5652
rect 9631 5528 10732 5556
rect 12176 5556 12204 5655
rect 13541 5627 13599 5633
rect 13541 5593 13553 5627
rect 13587 5624 13599 5627
rect 16960 5624 16988 5720
rect 17236 5692 17264 5723
rect 17310 5720 17316 5772
rect 17368 5760 17374 5772
rect 17773 5763 17831 5769
rect 17773 5760 17785 5763
rect 17368 5732 17785 5760
rect 17368 5720 17374 5732
rect 17773 5729 17785 5732
rect 17819 5760 17831 5763
rect 18874 5760 18880 5772
rect 17819 5732 18880 5760
rect 17819 5729 17831 5732
rect 17773 5723 17831 5729
rect 18874 5720 18880 5732
rect 18932 5760 18938 5772
rect 19076 5760 19104 5800
rect 19229 5797 19241 5831
rect 19229 5791 19248 5797
rect 19242 5788 19248 5791
rect 19300 5788 19306 5840
rect 19429 5831 19487 5837
rect 19429 5797 19441 5831
rect 19475 5828 19487 5831
rect 19794 5828 19800 5840
rect 19475 5800 19800 5828
rect 19475 5797 19487 5800
rect 19429 5791 19487 5797
rect 19794 5788 19800 5800
rect 19852 5788 19858 5840
rect 19886 5788 19892 5840
rect 19944 5788 19950 5840
rect 18932 5732 19104 5760
rect 19244 5760 19272 5788
rect 20088 5760 20116 5868
rect 20149 5865 20161 5868
rect 20195 5896 20207 5899
rect 20599 5899 20657 5905
rect 20599 5896 20611 5899
rect 20195 5868 20611 5896
rect 20195 5865 20207 5868
rect 20149 5859 20207 5865
rect 20599 5865 20611 5868
rect 20645 5865 20657 5899
rect 23566 5896 23572 5908
rect 20599 5859 20657 5865
rect 20824 5868 23572 5896
rect 20824 5837 20852 5868
rect 23566 5856 23572 5868
rect 23624 5856 23630 5908
rect 23937 5899 23995 5905
rect 23937 5865 23949 5899
rect 23983 5896 23995 5899
rect 24486 5896 24492 5908
rect 23983 5868 24492 5896
rect 23983 5865 23995 5868
rect 23937 5859 23995 5865
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 25314 5856 25320 5908
rect 25372 5896 25378 5908
rect 25409 5899 25467 5905
rect 25409 5896 25421 5899
rect 25372 5868 25421 5896
rect 25372 5856 25378 5868
rect 25409 5865 25421 5868
rect 25455 5896 25467 5899
rect 26326 5896 26332 5908
rect 25455 5868 26332 5896
rect 25455 5865 25467 5868
rect 25409 5859 25467 5865
rect 26326 5856 26332 5868
rect 26384 5856 26390 5908
rect 27798 5856 27804 5908
rect 27856 5896 27862 5908
rect 28442 5896 28448 5908
rect 27856 5868 28448 5896
rect 27856 5856 27862 5868
rect 28442 5856 28448 5868
rect 28500 5896 28506 5908
rect 28629 5899 28687 5905
rect 28629 5896 28641 5899
rect 28500 5868 28641 5896
rect 28500 5856 28506 5868
rect 28629 5865 28641 5868
rect 28675 5896 28687 5899
rect 29089 5899 29147 5905
rect 29089 5896 29101 5899
rect 28675 5868 29101 5896
rect 28675 5865 28687 5868
rect 28629 5859 28687 5865
rect 29089 5865 29101 5868
rect 29135 5865 29147 5899
rect 29089 5859 29147 5865
rect 29178 5856 29184 5908
rect 29236 5896 29242 5908
rect 30558 5896 30564 5908
rect 29236 5868 30564 5896
rect 29236 5856 29242 5868
rect 30558 5856 30564 5868
rect 30616 5896 30622 5908
rect 30616 5868 30880 5896
rect 30616 5856 30622 5868
rect 20349 5831 20407 5837
rect 20349 5797 20361 5831
rect 20395 5797 20407 5831
rect 20349 5791 20407 5797
rect 20809 5831 20867 5837
rect 20809 5797 20821 5831
rect 20855 5797 20867 5831
rect 20809 5791 20867 5797
rect 19244 5732 20116 5760
rect 18932 5720 18938 5732
rect 17494 5692 17500 5704
rect 17236 5664 17500 5692
rect 17494 5652 17500 5664
rect 17552 5692 17558 5704
rect 20364 5692 20392 5791
rect 21450 5788 21456 5840
rect 21508 5828 21514 5840
rect 21508 5800 21688 5828
rect 21508 5788 21514 5800
rect 21269 5763 21327 5769
rect 21269 5729 21281 5763
rect 21315 5760 21327 5763
rect 21358 5760 21364 5772
rect 21315 5732 21364 5760
rect 21315 5729 21327 5732
rect 21269 5723 21327 5729
rect 21358 5720 21364 5732
rect 21416 5720 21422 5772
rect 21542 5769 21548 5772
rect 21536 5723 21548 5769
rect 21542 5720 21548 5723
rect 21600 5720 21606 5772
rect 21660 5760 21688 5800
rect 21726 5788 21732 5840
rect 21784 5828 21790 5840
rect 22370 5828 22376 5840
rect 21784 5800 22376 5828
rect 21784 5788 21790 5800
rect 22370 5788 22376 5800
rect 22428 5788 22434 5840
rect 23198 5837 23204 5840
rect 23155 5831 23204 5837
rect 23155 5828 23167 5831
rect 22857 5800 23167 5828
rect 22857 5760 22885 5800
rect 23155 5797 23167 5800
rect 23201 5797 23204 5831
rect 23155 5791 23204 5797
rect 23198 5788 23204 5791
rect 23256 5788 23262 5840
rect 25130 5828 25136 5840
rect 24596 5800 25136 5828
rect 23476 5785 23534 5791
rect 21660 5732 22885 5760
rect 22940 5732 23244 5760
rect 22940 5692 22968 5732
rect 17552 5664 18460 5692
rect 20364 5664 21312 5692
rect 17552 5652 17558 5664
rect 18432 5633 18460 5664
rect 18417 5627 18475 5633
rect 13587 5596 16988 5624
rect 17512 5596 18092 5624
rect 13587 5593 13599 5596
rect 13541 5587 13599 5593
rect 17512 5568 17540 5596
rect 12434 5556 12440 5568
rect 12176 5528 12440 5556
rect 9631 5525 9643 5528
rect 9585 5519 9643 5525
rect 12434 5516 12440 5528
rect 12492 5516 12498 5568
rect 12894 5516 12900 5568
rect 12952 5556 12958 5568
rect 13262 5556 13268 5568
rect 12952 5528 13268 5556
rect 12952 5516 12958 5528
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 17494 5516 17500 5568
rect 17552 5516 17558 5568
rect 17862 5516 17868 5568
rect 17920 5516 17926 5568
rect 18064 5565 18092 5596
rect 18417 5593 18429 5627
rect 18463 5624 18475 5627
rect 18506 5624 18512 5636
rect 18463 5596 18512 5624
rect 18463 5593 18475 5596
rect 18417 5587 18475 5593
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 19521 5627 19579 5633
rect 18800 5596 19472 5624
rect 18800 5568 18828 5596
rect 18049 5559 18107 5565
rect 18049 5525 18061 5559
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 18782 5516 18788 5568
rect 18840 5516 18846 5568
rect 19058 5516 19064 5568
rect 19116 5556 19122 5568
rect 19245 5559 19303 5565
rect 19245 5556 19257 5559
rect 19116 5528 19257 5556
rect 19116 5516 19122 5528
rect 19245 5525 19257 5528
rect 19291 5525 19303 5559
rect 19444 5556 19472 5596
rect 19521 5593 19533 5627
rect 19567 5624 19579 5627
rect 19610 5624 19616 5636
rect 19567 5596 19616 5624
rect 19567 5593 19579 5596
rect 19521 5587 19579 5593
rect 19610 5584 19616 5596
rect 19668 5584 19674 5636
rect 19720 5596 20668 5624
rect 19720 5565 19748 5596
rect 19705 5559 19763 5565
rect 19705 5556 19717 5559
rect 19444 5528 19717 5556
rect 19245 5519 19303 5525
rect 19705 5525 19717 5528
rect 19751 5525 19763 5559
rect 19705 5519 19763 5525
rect 19978 5516 19984 5568
rect 20036 5516 20042 5568
rect 20180 5565 20208 5596
rect 20165 5559 20223 5565
rect 20165 5525 20177 5559
rect 20211 5525 20223 5559
rect 20165 5519 20223 5525
rect 20438 5516 20444 5568
rect 20496 5516 20502 5568
rect 20640 5565 20668 5596
rect 20625 5559 20683 5565
rect 20625 5525 20637 5559
rect 20671 5525 20683 5559
rect 21284 5556 21312 5664
rect 22848 5664 22968 5692
rect 22848 5636 22876 5664
rect 23014 5652 23020 5704
rect 23072 5652 23078 5704
rect 23216 5692 23244 5732
rect 23290 5720 23296 5772
rect 23348 5720 23354 5772
rect 23385 5763 23443 5769
rect 23385 5729 23397 5763
rect 23431 5729 23443 5763
rect 23476 5751 23488 5785
rect 23522 5751 23534 5785
rect 23476 5745 23534 5751
rect 23845 5763 23903 5769
rect 23491 5732 23520 5745
rect 23385 5723 23443 5729
rect 23400 5692 23428 5723
rect 23492 5704 23520 5732
rect 23845 5729 23857 5763
rect 23891 5760 23903 5763
rect 23934 5760 23940 5772
rect 23891 5732 23940 5760
rect 23891 5729 23903 5732
rect 23845 5723 23903 5729
rect 23934 5720 23940 5732
rect 23992 5760 23998 5772
rect 24596 5769 24624 5800
rect 25130 5788 25136 5800
rect 25188 5788 25194 5840
rect 26050 5828 26056 5840
rect 25240 5800 26056 5828
rect 25240 5769 25268 5800
rect 26050 5788 26056 5800
rect 26108 5788 26114 5840
rect 26234 5788 26240 5840
rect 26292 5828 26298 5840
rect 26292 5800 26648 5828
rect 26292 5788 26298 5800
rect 24489 5763 24547 5769
rect 24489 5760 24501 5763
rect 23992 5732 24501 5760
rect 23992 5720 23998 5732
rect 24489 5729 24501 5732
rect 24535 5729 24547 5763
rect 24489 5723 24547 5729
rect 24581 5763 24639 5769
rect 24581 5729 24593 5763
rect 24627 5729 24639 5763
rect 24581 5723 24639 5729
rect 24857 5763 24915 5769
rect 24857 5729 24869 5763
rect 24903 5760 24915 5763
rect 25225 5763 25283 5769
rect 24903 5732 25176 5760
rect 24903 5729 24915 5732
rect 24857 5723 24915 5729
rect 23216 5664 23428 5692
rect 23474 5652 23480 5704
rect 23532 5652 23538 5704
rect 23661 5695 23719 5701
rect 23661 5661 23673 5695
rect 23707 5692 23719 5695
rect 24302 5692 24308 5704
rect 23707 5664 24308 5692
rect 23707 5661 23719 5664
rect 23661 5655 23719 5661
rect 24302 5652 24308 5664
rect 24360 5652 24366 5704
rect 24504 5692 24532 5723
rect 24765 5695 24823 5701
rect 24765 5692 24777 5695
rect 24504 5664 24777 5692
rect 24765 5661 24777 5664
rect 24811 5692 24823 5695
rect 24946 5692 24952 5704
rect 24811 5664 24952 5692
rect 24811 5661 24823 5664
rect 24765 5655 24823 5661
rect 24946 5652 24952 5664
rect 25004 5652 25010 5704
rect 25148 5701 25176 5732
rect 25225 5729 25237 5763
rect 25271 5729 25283 5763
rect 25225 5723 25283 5729
rect 25501 5763 25559 5769
rect 25501 5729 25513 5763
rect 25547 5729 25559 5763
rect 26068 5760 26096 5788
rect 26620 5769 26648 5800
rect 27982 5788 27988 5840
rect 28040 5828 28046 5840
rect 29638 5828 29644 5840
rect 28040 5800 29644 5828
rect 28040 5788 28046 5800
rect 26513 5763 26571 5769
rect 26513 5760 26525 5763
rect 26068 5732 26525 5760
rect 25501 5723 25559 5729
rect 26513 5729 26525 5732
rect 26559 5729 26571 5763
rect 26513 5723 26571 5729
rect 26605 5763 26663 5769
rect 26605 5729 26617 5763
rect 26651 5729 26663 5763
rect 26605 5723 26663 5729
rect 25133 5695 25191 5701
rect 25133 5661 25145 5695
rect 25179 5692 25191 5695
rect 25314 5692 25320 5704
rect 25179 5664 25320 5692
rect 25179 5661 25191 5664
rect 25133 5655 25191 5661
rect 25314 5652 25320 5664
rect 25372 5652 25378 5704
rect 25516 5692 25544 5723
rect 27154 5720 27160 5772
rect 27212 5720 27218 5772
rect 28460 5769 28488 5800
rect 29638 5788 29644 5800
rect 29696 5828 29702 5840
rect 29696 5800 30788 5828
rect 29696 5788 29702 5800
rect 30760 5772 30788 5800
rect 28189 5763 28247 5769
rect 28189 5729 28201 5763
rect 28235 5760 28247 5763
rect 28445 5763 28503 5769
rect 28235 5732 28396 5760
rect 28235 5729 28247 5732
rect 28189 5723 28247 5729
rect 27172 5692 27200 5720
rect 25516 5664 27200 5692
rect 28368 5692 28396 5732
rect 28445 5729 28457 5763
rect 28491 5729 28503 5763
rect 28445 5723 28503 5729
rect 28534 5720 28540 5772
rect 28592 5760 28598 5772
rect 28721 5763 28779 5769
rect 28721 5760 28733 5763
rect 28592 5732 28733 5760
rect 28592 5720 28598 5732
rect 28721 5729 28733 5732
rect 28767 5760 28779 5763
rect 29086 5760 29092 5772
rect 28767 5732 29092 5760
rect 28767 5729 28779 5732
rect 28721 5723 28779 5729
rect 29086 5720 29092 5732
rect 29144 5720 29150 5772
rect 29178 5720 29184 5772
rect 29236 5720 29242 5772
rect 29362 5720 29368 5772
rect 29420 5720 29426 5772
rect 30489 5763 30547 5769
rect 30489 5729 30501 5763
rect 30535 5760 30547 5763
rect 30650 5760 30656 5772
rect 30535 5732 30656 5760
rect 30535 5729 30547 5732
rect 30489 5723 30547 5729
rect 30650 5720 30656 5732
rect 30708 5720 30714 5772
rect 30742 5720 30748 5772
rect 30800 5720 30806 5772
rect 30852 5769 30880 5868
rect 30926 5856 30932 5908
rect 30984 5856 30990 5908
rect 30837 5763 30895 5769
rect 30837 5729 30849 5763
rect 30883 5729 30895 5763
rect 30837 5723 30895 5729
rect 29380 5692 29408 5720
rect 28368 5664 29408 5692
rect 22572 5596 22768 5624
rect 22572 5556 22600 5596
rect 21284 5528 22600 5556
rect 20625 5519 20683 5525
rect 22646 5516 22652 5568
rect 22704 5516 22710 5568
rect 22740 5556 22768 5596
rect 22830 5584 22836 5636
rect 22888 5584 22894 5636
rect 22922 5584 22928 5636
rect 22980 5624 22986 5636
rect 27065 5627 27123 5633
rect 27065 5624 27077 5627
rect 22980 5596 27077 5624
rect 22980 5584 22986 5596
rect 27065 5593 27077 5596
rect 27111 5593 27123 5627
rect 27065 5587 27123 5593
rect 29362 5584 29368 5636
rect 29420 5584 29426 5636
rect 25038 5556 25044 5568
rect 22740 5528 25044 5556
rect 25038 5516 25044 5528
rect 25096 5516 25102 5568
rect 552 5466 31372 5488
rect 552 5414 4250 5466
rect 4302 5414 4314 5466
rect 4366 5414 4378 5466
rect 4430 5414 4442 5466
rect 4494 5414 4506 5466
rect 4558 5414 11955 5466
rect 12007 5414 12019 5466
rect 12071 5414 12083 5466
rect 12135 5414 12147 5466
rect 12199 5414 12211 5466
rect 12263 5414 19660 5466
rect 19712 5414 19724 5466
rect 19776 5414 19788 5466
rect 19840 5414 19852 5466
rect 19904 5414 19916 5466
rect 19968 5414 27365 5466
rect 27417 5414 27429 5466
rect 27481 5414 27493 5466
rect 27545 5414 27557 5466
rect 27609 5414 27621 5466
rect 27673 5414 31372 5466
rect 552 5392 31372 5414
rect 1397 5355 1455 5361
rect 1397 5321 1409 5355
rect 1443 5352 1455 5355
rect 1949 5355 2007 5361
rect 1949 5352 1961 5355
rect 1443 5324 1961 5352
rect 1443 5321 1455 5324
rect 1397 5315 1455 5321
rect 1949 5321 1961 5324
rect 1995 5352 2007 5355
rect 2222 5352 2228 5364
rect 1995 5324 2228 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 2406 5312 2412 5364
rect 2464 5312 2470 5364
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 2590 5352 2596 5364
rect 2547 5324 2596 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 4801 5355 4859 5361
rect 4801 5321 4813 5355
rect 4847 5352 4859 5355
rect 4982 5352 4988 5364
rect 4847 5324 4988 5352
rect 4847 5321 4859 5324
rect 4801 5315 4859 5321
rect 4982 5312 4988 5324
rect 5040 5352 5046 5364
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 5040 5324 5365 5352
rect 5040 5312 5046 5324
rect 2225 5219 2283 5225
rect 2225 5216 2237 5219
rect 2056 5188 2237 5216
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5148 1547 5151
rect 1670 5148 1676 5160
rect 1535 5120 1676 5148
rect 1535 5117 1547 5120
rect 1489 5111 1547 5117
rect 1670 5108 1676 5120
rect 1728 5108 1734 5160
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5148 1823 5151
rect 1946 5148 1952 5160
rect 1811 5120 1952 5148
rect 1811 5117 1823 5120
rect 1765 5111 1823 5117
rect 1946 5108 1952 5120
rect 2004 5108 2010 5160
rect 2056 5157 2084 5188
rect 2225 5185 2237 5188
rect 2271 5216 2283 5219
rect 2424 5216 2452 5312
rect 2271 5188 2452 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2041 5151 2099 5157
rect 2041 5117 2053 5151
rect 2087 5117 2099 5151
rect 2041 5111 2099 5117
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 2409 5151 2467 5157
rect 2409 5148 2421 5151
rect 2363 5120 2421 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 2409 5117 2421 5120
rect 2455 5117 2467 5151
rect 2608 5148 2636 5312
rect 4249 5287 4307 5293
rect 4249 5253 4261 5287
rect 4295 5284 4307 5287
rect 4890 5284 4896 5296
rect 4295 5256 4896 5284
rect 4295 5253 4307 5256
rect 4249 5247 4307 5253
rect 4890 5244 4896 5256
rect 4948 5244 4954 5296
rect 5074 5244 5080 5296
rect 5132 5244 5138 5296
rect 2685 5151 2743 5157
rect 2685 5148 2697 5151
rect 2608 5120 2697 5148
rect 2409 5111 2467 5117
rect 2685 5117 2697 5120
rect 2731 5117 2743 5151
rect 2685 5111 2743 5117
rect 2424 5080 2452 5111
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 3789 5151 3847 5157
rect 3789 5148 3801 5151
rect 3200 5120 3801 5148
rect 3200 5108 3206 5120
rect 3789 5117 3801 5120
rect 3835 5117 3847 5151
rect 3789 5111 3847 5117
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5148 4123 5151
rect 4154 5148 4160 5160
rect 4111 5120 4160 5148
rect 4111 5117 4123 5120
rect 4065 5111 4123 5117
rect 4154 5108 4160 5120
rect 4212 5148 4218 5160
rect 5184 5157 5212 5324
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 5353 5315 5411 5321
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 6181 5355 6239 5361
rect 6181 5352 6193 5355
rect 5500 5324 6193 5352
rect 5500 5312 5506 5324
rect 6181 5321 6193 5324
rect 6227 5352 6239 5355
rect 7009 5355 7067 5361
rect 7009 5352 7021 5355
rect 6227 5324 7021 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 7009 5321 7021 5324
rect 7055 5352 7067 5355
rect 9214 5352 9220 5364
rect 7055 5324 9220 5352
rect 7055 5321 7067 5324
rect 7009 5315 7067 5321
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 9401 5355 9459 5361
rect 9401 5321 9413 5355
rect 9447 5352 9459 5355
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 9447 5324 9689 5352
rect 9447 5321 9459 5324
rect 9401 5315 9459 5321
rect 9677 5321 9689 5324
rect 9723 5352 9735 5355
rect 9950 5352 9956 5364
rect 9723 5324 9956 5352
rect 9723 5321 9735 5324
rect 9677 5315 9735 5321
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 10229 5355 10287 5361
rect 10229 5321 10241 5355
rect 10275 5352 10287 5355
rect 10318 5352 10324 5364
rect 10275 5324 10324 5352
rect 10275 5321 10287 5324
rect 10229 5315 10287 5321
rect 5460 5216 5488 5312
rect 7742 5284 7748 5296
rect 5368 5188 5488 5216
rect 6564 5256 7748 5284
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 4212 5120 4353 5148
rect 4212 5108 4218 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 4893 5151 4951 5157
rect 4893 5117 4905 5151
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 5169 5151 5227 5157
rect 5169 5117 5181 5151
rect 5215 5117 5227 5151
rect 5169 5111 5227 5117
rect 3510 5080 3516 5092
rect 2424 5052 3516 5080
rect 3510 5040 3516 5052
rect 3568 5080 3574 5092
rect 3697 5083 3755 5089
rect 3697 5080 3709 5083
rect 3568 5052 3709 5080
rect 3568 5040 3574 5052
rect 3697 5049 3709 5052
rect 3743 5080 3755 5083
rect 3973 5083 4031 5089
rect 3973 5080 3985 5083
rect 3743 5052 3985 5080
rect 3743 5049 3755 5052
rect 3697 5043 3755 5049
rect 3973 5049 3985 5052
rect 4019 5049 4031 5083
rect 4908 5080 4936 5111
rect 5368 5080 5396 5188
rect 6564 5157 6592 5256
rect 7742 5244 7748 5256
rect 7800 5244 7806 5296
rect 8202 5244 8208 5296
rect 8260 5284 8266 5296
rect 8573 5287 8631 5293
rect 8573 5284 8585 5287
rect 8260 5256 8585 5284
rect 8260 5244 8266 5256
rect 8573 5253 8585 5256
rect 8619 5284 8631 5287
rect 9490 5284 9496 5296
rect 8619 5256 9496 5284
rect 8619 5253 8631 5256
rect 8573 5247 8631 5253
rect 9490 5244 9496 5256
rect 9548 5244 9554 5296
rect 9968 5284 9996 5312
rect 9968 5256 10180 5284
rect 8220 5216 8248 5244
rect 8849 5219 8907 5225
rect 8849 5216 8861 5219
rect 7668 5188 8248 5216
rect 8680 5188 8861 5216
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5148 5503 5151
rect 5537 5151 5595 5157
rect 5537 5148 5549 5151
rect 5491 5120 5549 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 5537 5117 5549 5120
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5997 5151 6055 5157
rect 5997 5148 6009 5151
rect 5675 5120 6009 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5997 5117 6009 5120
rect 6043 5148 6055 5151
rect 6273 5151 6331 5157
rect 6273 5148 6285 5151
rect 6043 5120 6285 5148
rect 6043 5117 6055 5120
rect 5997 5111 6055 5117
rect 6273 5117 6285 5120
rect 6319 5148 6331 5151
rect 6457 5151 6515 5157
rect 6457 5148 6469 5151
rect 6319 5120 6469 5148
rect 6319 5117 6331 5120
rect 6273 5111 6331 5117
rect 6457 5117 6469 5120
rect 6503 5117 6515 5151
rect 6457 5111 6515 5117
rect 6549 5151 6607 5157
rect 6549 5117 6561 5151
rect 6595 5117 6607 5151
rect 6549 5111 6607 5117
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 6871 5120 7113 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 7101 5117 7113 5120
rect 7147 5148 7159 5151
rect 7282 5148 7288 5160
rect 7147 5120 7288 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 4908 5052 5396 5080
rect 5552 5080 5580 5111
rect 7282 5108 7288 5120
rect 7340 5108 7346 5160
rect 7668 5157 7696 5188
rect 8680 5157 8708 5188
rect 8849 5185 8861 5188
rect 8895 5216 8907 5219
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 8895 5188 9965 5216
rect 8895 5185 8907 5188
rect 8849 5179 8907 5185
rect 9232 5157 9260 5188
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 7653 5151 7711 5157
rect 7423 5120 7604 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 7576 5089 7604 5120
rect 7653 5117 7665 5151
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 7975 5120 8125 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 8665 5151 8723 5157
rect 8665 5117 8677 5151
rect 8711 5117 8723 5151
rect 8665 5111 8723 5117
rect 8941 5151 8999 5157
rect 8941 5117 8953 5151
rect 8987 5117 8999 5151
rect 8941 5111 8999 5117
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5117 9275 5151
rect 9217 5111 9275 5117
rect 6733 5083 6791 5089
rect 6733 5080 6745 5083
rect 5552 5052 6745 5080
rect 3973 5043 4031 5049
rect 6733 5049 6745 5052
rect 6779 5080 6791 5083
rect 7561 5083 7619 5089
rect 6779 5052 7328 5080
rect 6779 5049 6791 5052
rect 6733 5043 6791 5049
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 2777 5015 2835 5021
rect 2777 5012 2789 5015
rect 1452 4984 2789 5012
rect 1452 4972 1458 4984
rect 2777 4981 2789 4984
rect 2823 4981 2835 5015
rect 2777 4975 2835 4981
rect 5074 4972 5080 5024
rect 5132 5012 5138 5024
rect 7300 5021 7328 5052
rect 7561 5049 7573 5083
rect 7607 5080 7619 5083
rect 7944 5080 7972 5111
rect 7607 5052 7972 5080
rect 8220 5080 8248 5111
rect 8956 5080 8984 5111
rect 9306 5108 9312 5160
rect 9364 5108 9370 5160
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 10152 5157 10180 5256
rect 10045 5151 10103 5157
rect 10045 5148 10057 5151
rect 9824 5120 10057 5148
rect 9824 5108 9830 5120
rect 10045 5117 10057 5120
rect 10091 5117 10103 5151
rect 10045 5111 10103 5117
rect 10137 5151 10195 5157
rect 10137 5117 10149 5151
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 10244 5080 10272 5315
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 12342 5352 12348 5364
rect 10468 5324 12348 5352
rect 10468 5312 10474 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 13173 5355 13231 5361
rect 13173 5321 13185 5355
rect 13219 5352 13231 5355
rect 14090 5352 14096 5364
rect 13219 5324 14096 5352
rect 13219 5321 13231 5324
rect 13173 5315 13231 5321
rect 14090 5312 14096 5324
rect 14148 5352 14154 5364
rect 14277 5355 14335 5361
rect 14277 5352 14289 5355
rect 14148 5324 14289 5352
rect 14148 5312 14154 5324
rect 14277 5321 14289 5324
rect 14323 5321 14335 5355
rect 14277 5315 14335 5321
rect 14461 5355 14519 5361
rect 14461 5321 14473 5355
rect 14507 5352 14519 5355
rect 15378 5352 15384 5364
rect 14507 5324 15384 5352
rect 14507 5321 14519 5324
rect 14461 5315 14519 5321
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 15930 5312 15936 5364
rect 15988 5352 15994 5364
rect 16298 5352 16304 5364
rect 15988 5324 16304 5352
rect 15988 5312 15994 5324
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 16408 5324 17080 5352
rect 11977 5287 12035 5293
rect 11977 5253 11989 5287
rect 12023 5284 12035 5287
rect 13078 5284 13084 5296
rect 12023 5256 13084 5284
rect 12023 5253 12035 5256
rect 11977 5247 12035 5253
rect 13078 5244 13084 5256
rect 13136 5244 13142 5296
rect 13357 5287 13415 5293
rect 13357 5253 13369 5287
rect 13403 5253 13415 5287
rect 13357 5247 13415 5253
rect 15289 5287 15347 5293
rect 15289 5253 15301 5287
rect 15335 5284 15347 5287
rect 15562 5284 15568 5296
rect 15335 5256 15568 5284
rect 15335 5253 15347 5256
rect 15289 5247 15347 5253
rect 10594 5176 10600 5228
rect 10652 5176 10658 5228
rect 13372 5216 13400 5247
rect 15562 5244 15568 5256
rect 15620 5244 15626 5296
rect 16408 5216 16436 5324
rect 16482 5244 16488 5296
rect 16540 5284 16546 5296
rect 16945 5287 17003 5293
rect 16945 5284 16957 5287
rect 16540 5256 16957 5284
rect 16540 5244 16546 5256
rect 16945 5253 16957 5256
rect 16991 5253 17003 5287
rect 17052 5284 17080 5324
rect 18782 5312 18788 5364
rect 18840 5352 18846 5364
rect 18877 5355 18935 5361
rect 18877 5352 18889 5355
rect 18840 5324 18889 5352
rect 18840 5312 18846 5324
rect 18877 5321 18889 5324
rect 18923 5321 18935 5355
rect 18877 5315 18935 5321
rect 19518 5312 19524 5364
rect 19576 5352 19582 5364
rect 19705 5355 19763 5361
rect 19705 5352 19717 5355
rect 19576 5324 19717 5352
rect 19576 5312 19582 5324
rect 19705 5321 19717 5324
rect 19751 5321 19763 5355
rect 19705 5315 19763 5321
rect 19797 5355 19855 5361
rect 19797 5321 19809 5355
rect 19843 5352 19855 5355
rect 19978 5352 19984 5364
rect 19843 5324 19984 5352
rect 19843 5321 19855 5324
rect 19797 5315 19855 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20254 5312 20260 5364
rect 20312 5312 20318 5364
rect 20438 5312 20444 5364
rect 20496 5352 20502 5364
rect 20625 5355 20683 5361
rect 20625 5352 20637 5355
rect 20496 5324 20637 5352
rect 20496 5312 20502 5324
rect 20625 5321 20637 5324
rect 20671 5321 20683 5355
rect 20625 5315 20683 5321
rect 20714 5312 20720 5364
rect 20772 5312 20778 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 20864 5324 23520 5352
rect 20864 5312 20870 5324
rect 20990 5284 20996 5296
rect 17052 5256 19932 5284
rect 16945 5247 17003 5253
rect 13372 5188 16436 5216
rect 13446 5108 13452 5160
rect 13504 5148 13510 5160
rect 15378 5148 15384 5160
rect 13504 5120 15384 5148
rect 13504 5108 13510 5120
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 15488 5120 15577 5148
rect 10842 5083 10900 5089
rect 10842 5080 10854 5083
rect 8220 5052 10272 5080
rect 10336 5052 10854 5080
rect 7607 5049 7619 5052
rect 7561 5043 7619 5049
rect 5905 5015 5963 5021
rect 5905 5012 5917 5015
rect 5132 4984 5917 5012
rect 5132 4972 5138 4984
rect 5905 4981 5917 4984
rect 5951 4981 5963 5015
rect 5905 4975 5963 4981
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 7374 5012 7380 5024
rect 7331 4984 7380 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 7800 4984 7849 5012
rect 7800 4972 7806 4984
rect 7837 4981 7849 4984
rect 7883 5012 7895 5015
rect 9125 5015 9183 5021
rect 9125 5012 9137 5015
rect 7883 4984 9137 5012
rect 7883 4981 7895 4984
rect 7837 4975 7895 4981
rect 9125 4981 9137 4984
rect 9171 5012 9183 5015
rect 10336 5012 10364 5052
rect 10842 5049 10854 5052
rect 10888 5049 10900 5083
rect 12158 5080 12164 5092
rect 10842 5043 10900 5049
rect 10980 5052 12164 5080
rect 9171 4984 10364 5012
rect 9171 4981 9183 4984
rect 9125 4975 9183 4981
rect 10410 4972 10416 5024
rect 10468 5012 10474 5024
rect 10980 5012 11008 5052
rect 12158 5040 12164 5052
rect 12216 5040 12222 5092
rect 12986 5040 12992 5092
rect 13044 5040 13050 5092
rect 14093 5083 14151 5089
rect 14093 5080 14105 5083
rect 13096 5052 14105 5080
rect 10468 4984 11008 5012
rect 10468 4972 10474 4984
rect 11238 4972 11244 5024
rect 11296 5012 11302 5024
rect 13096 5012 13124 5052
rect 14093 5049 14105 5052
rect 14139 5049 14151 5083
rect 14093 5043 14151 5049
rect 15010 5040 15016 5092
rect 15068 5040 15074 5092
rect 15488 5080 15516 5120
rect 15565 5117 15577 5120
rect 15611 5117 15623 5151
rect 15565 5111 15623 5117
rect 15654 5108 15660 5160
rect 15712 5148 15718 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15712 5120 15761 5148
rect 15712 5108 15718 5120
rect 15749 5117 15761 5120
rect 15795 5117 15807 5151
rect 15749 5111 15807 5117
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5117 16175 5151
rect 16117 5111 16175 5117
rect 16132 5080 16160 5111
rect 16206 5108 16212 5160
rect 16264 5108 16270 5160
rect 16960 5148 16988 5247
rect 18414 5176 18420 5228
rect 18472 5216 18478 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 18472 5188 19441 5216
rect 18472 5176 18478 5188
rect 19429 5185 19441 5188
rect 19475 5185 19487 5219
rect 19429 5179 19487 5185
rect 19518 5176 19524 5228
rect 19576 5176 19582 5228
rect 19904 5225 19932 5256
rect 20180 5256 20996 5284
rect 19889 5219 19947 5225
rect 19889 5185 19901 5219
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 17494 5148 17500 5160
rect 16960 5120 17500 5148
rect 17494 5108 17500 5120
rect 17552 5108 17558 5160
rect 17589 5151 17647 5157
rect 17589 5117 17601 5151
rect 17635 5117 17647 5151
rect 19150 5148 19156 5160
rect 17589 5111 17647 5117
rect 18616 5120 19156 5148
rect 15488 5052 16160 5080
rect 15488 5024 15516 5052
rect 11296 4984 13124 5012
rect 13199 5015 13257 5021
rect 11296 4972 11302 4984
rect 13199 4981 13211 5015
rect 13245 5012 13257 5015
rect 14303 5015 14361 5021
rect 14303 5012 14315 5015
rect 13245 4984 14315 5012
rect 13245 4981 13257 4984
rect 13199 4975 13257 4981
rect 14303 4981 14315 4984
rect 14349 5012 14361 5015
rect 14734 5012 14740 5024
rect 14349 4984 14740 5012
rect 14349 4981 14361 4984
rect 14303 4975 14361 4981
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 15470 4972 15476 5024
rect 15528 4972 15534 5024
rect 16224 5012 16252 5108
rect 16390 5040 16396 5092
rect 16448 5080 16454 5092
rect 16850 5080 16856 5092
rect 16448 5052 16856 5080
rect 16448 5040 16454 5052
rect 16850 5040 16856 5052
rect 16908 5080 16914 5092
rect 17221 5083 17279 5089
rect 17221 5080 17233 5083
rect 16908 5052 17233 5080
rect 16908 5040 16914 5052
rect 17221 5049 17233 5052
rect 17267 5080 17279 5083
rect 17604 5080 17632 5111
rect 17267 5052 17632 5080
rect 17267 5049 17279 5052
rect 17221 5043 17279 5049
rect 16301 5015 16359 5021
rect 16301 5012 16313 5015
rect 16224 4984 16313 5012
rect 16301 4981 16313 4984
rect 16347 4981 16359 5015
rect 16301 4975 16359 4981
rect 16574 4972 16580 5024
rect 16632 5012 16638 5024
rect 16761 5015 16819 5021
rect 16761 5012 16773 5015
rect 16632 4984 16773 5012
rect 16632 4972 16638 4984
rect 16761 4981 16773 4984
rect 16807 4981 16819 5015
rect 16761 4975 16819 4981
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17313 5015 17371 5021
rect 17313 5012 17325 5015
rect 17000 4984 17325 5012
rect 17000 4972 17006 4984
rect 17313 4981 17325 4984
rect 17359 5012 17371 5015
rect 18616 5012 18644 5120
rect 19150 5108 19156 5120
rect 19208 5108 19214 5160
rect 18874 5089 18880 5092
rect 18861 5083 18880 5089
rect 18861 5049 18873 5083
rect 18861 5043 18880 5049
rect 18874 5040 18880 5043
rect 18932 5040 18938 5092
rect 19061 5083 19119 5089
rect 19061 5049 19073 5083
rect 19107 5049 19119 5083
rect 19536 5080 19564 5176
rect 19978 5108 19984 5160
rect 20036 5108 20042 5160
rect 20180 5157 20208 5256
rect 20990 5244 20996 5256
rect 21048 5244 21054 5296
rect 22922 5244 22928 5296
rect 22980 5284 22986 5296
rect 23106 5284 23112 5296
rect 22980 5256 23112 5284
rect 22980 5244 22986 5256
rect 23106 5244 23112 5256
rect 23164 5244 23170 5296
rect 23492 5284 23520 5324
rect 23566 5312 23572 5364
rect 23624 5352 23630 5364
rect 23845 5355 23903 5361
rect 23845 5352 23857 5355
rect 23624 5324 23857 5352
rect 23624 5312 23630 5324
rect 23845 5321 23857 5324
rect 23891 5321 23903 5355
rect 24854 5352 24860 5364
rect 23845 5315 23903 5321
rect 23952 5324 24860 5352
rect 23952 5284 23980 5324
rect 24854 5312 24860 5324
rect 24912 5312 24918 5364
rect 25038 5312 25044 5364
rect 25096 5352 25102 5364
rect 25317 5355 25375 5361
rect 25317 5352 25329 5355
rect 25096 5324 25329 5352
rect 25096 5312 25102 5324
rect 25317 5321 25329 5324
rect 25363 5321 25375 5355
rect 25317 5315 25375 5321
rect 28445 5355 28503 5361
rect 28445 5321 28457 5355
rect 28491 5352 28503 5355
rect 28718 5352 28724 5364
rect 28491 5324 28724 5352
rect 28491 5321 28503 5324
rect 28445 5315 28503 5321
rect 28718 5312 28724 5324
rect 28776 5312 28782 5364
rect 28920 5324 30512 5352
rect 28920 5296 28948 5324
rect 23492 5256 23980 5284
rect 28902 5244 28908 5296
rect 28960 5244 28966 5296
rect 30374 5244 30380 5296
rect 30432 5244 30438 5296
rect 20622 5176 20628 5228
rect 20680 5216 20686 5228
rect 22557 5219 22615 5225
rect 22557 5216 22569 5219
rect 20680 5188 22569 5216
rect 20680 5176 20686 5188
rect 22557 5185 22569 5188
rect 22603 5185 22615 5219
rect 22557 5179 22615 5185
rect 22646 5176 22652 5228
rect 22704 5216 22710 5228
rect 23201 5219 23259 5225
rect 23201 5216 23213 5219
rect 22704 5188 23213 5216
rect 22704 5176 22710 5188
rect 23201 5185 23213 5188
rect 23247 5185 23259 5219
rect 23201 5179 23259 5185
rect 25225 5219 25283 5225
rect 25225 5185 25237 5219
rect 25271 5216 25283 5219
rect 25406 5216 25412 5228
rect 25271 5188 25412 5216
rect 25271 5185 25283 5188
rect 25225 5179 25283 5185
rect 25406 5176 25412 5188
rect 25464 5176 25470 5228
rect 28997 5219 29055 5225
rect 28997 5216 29009 5219
rect 28000 5188 29009 5216
rect 20165 5151 20223 5157
rect 20165 5117 20177 5151
rect 20211 5148 20223 5151
rect 20254 5148 20260 5160
rect 20211 5120 20260 5148
rect 20211 5117 20223 5120
rect 20165 5111 20223 5117
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 20533 5151 20591 5157
rect 20533 5117 20545 5151
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 20548 5080 20576 5111
rect 20990 5108 20996 5160
rect 21048 5108 21054 5160
rect 21634 5108 21640 5160
rect 21692 5148 21698 5160
rect 23106 5157 23112 5160
rect 22741 5151 22799 5157
rect 22741 5148 22753 5151
rect 21692 5120 22753 5148
rect 21692 5108 21698 5120
rect 22741 5117 22753 5120
rect 22787 5117 22799 5151
rect 22741 5111 22799 5117
rect 23063 5151 23112 5157
rect 23063 5117 23075 5151
rect 23109 5117 23112 5151
rect 23063 5111 23112 5117
rect 23106 5108 23112 5111
rect 23164 5108 23170 5160
rect 24946 5108 24952 5160
rect 25004 5157 25010 5160
rect 25004 5111 25016 5157
rect 25424 5148 25452 5176
rect 28000 5160 28028 5188
rect 28997 5185 29009 5188
rect 29043 5185 29055 5219
rect 28997 5179 29055 5185
rect 26697 5151 26755 5157
rect 26697 5148 26709 5151
rect 25424 5120 26709 5148
rect 26697 5117 26709 5120
rect 26743 5117 26755 5151
rect 26697 5111 26755 5117
rect 25004 5108 25010 5111
rect 27154 5108 27160 5160
rect 27212 5108 27218 5160
rect 27982 5108 27988 5160
rect 28040 5108 28046 5160
rect 28537 5151 28595 5157
rect 28537 5117 28549 5151
rect 28583 5148 28595 5151
rect 28626 5148 28632 5160
rect 28583 5120 28632 5148
rect 28583 5117 28595 5120
rect 28537 5111 28595 5117
rect 28626 5108 28632 5120
rect 28684 5108 28690 5160
rect 28813 5151 28871 5157
rect 28813 5117 28825 5151
rect 28859 5148 28871 5151
rect 28902 5148 28908 5160
rect 28859 5120 28908 5148
rect 28859 5117 28871 5120
rect 28813 5111 28871 5117
rect 28902 5108 28908 5120
rect 28960 5108 28966 5160
rect 29270 5157 29276 5160
rect 29264 5148 29276 5157
rect 29231 5120 29276 5148
rect 29264 5111 29276 5120
rect 29270 5108 29276 5111
rect 29328 5108 29334 5160
rect 30392 5148 30420 5244
rect 30484 5216 30512 5324
rect 30558 5312 30564 5364
rect 30616 5312 30622 5364
rect 30484 5188 30788 5216
rect 30760 5157 30788 5188
rect 30653 5151 30711 5157
rect 30653 5148 30665 5151
rect 30392 5120 30665 5148
rect 30653 5117 30665 5120
rect 30699 5117 30711 5151
rect 30653 5111 30711 5117
rect 30745 5151 30803 5157
rect 30745 5117 30757 5151
rect 30791 5117 30803 5151
rect 30745 5111 30803 5117
rect 19536 5052 20576 5080
rect 20916 5052 22784 5080
rect 19061 5043 19119 5049
rect 17359 4984 18644 5012
rect 17359 4981 17371 4984
rect 17313 4975 17371 4981
rect 18690 4972 18696 5024
rect 18748 4972 18754 5024
rect 19076 5012 19104 5043
rect 20806 5012 20812 5024
rect 19076 4984 20812 5012
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 20916 5021 20944 5052
rect 20901 5015 20959 5021
rect 20901 4981 20913 5015
rect 20947 4981 20959 5015
rect 22756 5012 22784 5052
rect 22830 5040 22836 5092
rect 22888 5040 22894 5092
rect 22925 5083 22983 5089
rect 22925 5049 22937 5083
rect 22971 5080 22983 5083
rect 23842 5080 23848 5092
rect 22971 5052 23848 5080
rect 22971 5049 22983 5052
rect 22925 5043 22983 5049
rect 23842 5040 23848 5052
rect 23900 5040 23906 5092
rect 24854 5040 24860 5092
rect 24912 5040 24918 5092
rect 26452 5083 26510 5089
rect 26452 5049 26464 5083
rect 26498 5080 26510 5083
rect 27172 5080 27200 5108
rect 30668 5080 30696 5111
rect 30837 5083 30895 5089
rect 30837 5080 30849 5083
rect 26498 5052 27200 5080
rect 27632 5052 30420 5080
rect 30668 5052 30849 5080
rect 26498 5049 26510 5052
rect 26452 5043 26510 5049
rect 23106 5012 23112 5024
rect 22756 4984 23112 5012
rect 20901 4975 20959 4981
rect 23106 4972 23112 4984
rect 23164 4972 23170 5024
rect 23198 4972 23204 5024
rect 23256 5012 23262 5024
rect 23474 5012 23480 5024
rect 23256 4984 23480 5012
rect 23256 4972 23262 4984
rect 23474 4972 23480 4984
rect 23532 4972 23538 5024
rect 24872 5012 24900 5040
rect 27632 5012 27660 5052
rect 30392 5021 30420 5052
rect 30837 5049 30849 5052
rect 30883 5049 30895 5083
rect 30837 5043 30895 5049
rect 24872 4984 27660 5012
rect 30377 5015 30435 5021
rect 30377 4981 30389 5015
rect 30423 4981 30435 5015
rect 30377 4975 30435 4981
rect 552 4922 31531 4944
rect 552 4870 8102 4922
rect 8154 4870 8166 4922
rect 8218 4870 8230 4922
rect 8282 4870 8294 4922
rect 8346 4870 8358 4922
rect 8410 4870 15807 4922
rect 15859 4870 15871 4922
rect 15923 4870 15935 4922
rect 15987 4870 15999 4922
rect 16051 4870 16063 4922
rect 16115 4870 23512 4922
rect 23564 4870 23576 4922
rect 23628 4870 23640 4922
rect 23692 4870 23704 4922
rect 23756 4870 23768 4922
rect 23820 4870 31217 4922
rect 31269 4870 31281 4922
rect 31333 4870 31345 4922
rect 31397 4870 31409 4922
rect 31461 4870 31473 4922
rect 31525 4870 31531 4922
rect 552 4848 31531 4870
rect 1394 4768 1400 4820
rect 1452 4768 1458 4820
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 1765 4811 1823 4817
rect 1765 4808 1777 4811
rect 1728 4780 1777 4808
rect 1728 4768 1734 4780
rect 1765 4777 1777 4780
rect 1811 4777 1823 4811
rect 1765 4771 1823 4777
rect 1946 4768 1952 4820
rect 2004 4808 2010 4820
rect 3050 4808 3056 4820
rect 2004 4780 3056 4808
rect 2004 4768 2010 4780
rect 3050 4768 3056 4780
rect 3108 4808 3114 4820
rect 3108 4780 3648 4808
rect 3108 4768 3114 4780
rect 1412 4740 1440 4768
rect 1320 4712 1440 4740
rect 1029 4675 1087 4681
rect 1029 4641 1041 4675
rect 1075 4672 1087 4675
rect 1210 4672 1216 4684
rect 1075 4644 1216 4672
rect 1075 4641 1087 4644
rect 1029 4635 1087 4641
rect 1210 4632 1216 4644
rect 1268 4632 1274 4684
rect 1320 4681 1348 4712
rect 1305 4675 1363 4681
rect 1305 4641 1317 4675
rect 1351 4641 1363 4675
rect 1305 4635 1363 4641
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1688 4672 1716 4768
rect 2682 4740 2688 4752
rect 2056 4712 2688 4740
rect 2056 4681 2084 4712
rect 2682 4700 2688 4712
rect 2740 4740 2746 4752
rect 3620 4740 3648 4780
rect 7190 4768 7196 4820
rect 7248 4768 7254 4820
rect 8665 4811 8723 4817
rect 8665 4777 8677 4811
rect 8711 4808 8723 4811
rect 11330 4808 11336 4820
rect 8711 4780 11336 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11451 4811 11509 4817
rect 11451 4777 11463 4811
rect 11497 4808 11509 4811
rect 11497 4780 11836 4808
rect 11497 4777 11509 4780
rect 11451 4771 11509 4777
rect 3758 4743 3816 4749
rect 3758 4740 3770 4743
rect 2740 4712 3556 4740
rect 3620 4712 3770 4740
rect 2740 4700 2746 4712
rect 1443 4644 1716 4672
rect 1857 4675 1915 4681
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1857 4641 1869 4675
rect 1903 4641 1915 4675
rect 1857 4635 1915 4641
rect 2041 4675 2099 4681
rect 2041 4641 2053 4675
rect 2087 4641 2099 4675
rect 2297 4675 2355 4681
rect 2297 4672 2309 4675
rect 2041 4635 2099 4641
rect 2148 4644 2309 4672
rect 1320 4604 1348 4635
rect 1872 4604 1900 4635
rect 2148 4604 2176 4644
rect 2297 4641 2309 4644
rect 2343 4641 2355 4675
rect 2297 4635 2355 4641
rect 3528 4616 3556 4712
rect 3758 4709 3770 4712
rect 3804 4709 3816 4743
rect 6914 4740 6920 4752
rect 3758 4703 3816 4709
rect 5828 4712 6920 4740
rect 5828 4681 5856 4712
rect 6914 4700 6920 4712
rect 6972 4740 6978 4752
rect 6972 4712 7328 4740
rect 6972 4700 6978 4712
rect 5813 4675 5871 4681
rect 5813 4641 5825 4675
rect 5859 4641 5871 4675
rect 6069 4675 6127 4681
rect 6069 4672 6081 4675
rect 5813 4635 5871 4641
rect 5920 4644 6081 4672
rect 1320 4576 1900 4604
rect 2056 4576 2176 4604
rect 2056 4536 2084 4576
rect 3510 4564 3516 4616
rect 3568 4564 3574 4616
rect 5920 4604 5948 4644
rect 6069 4641 6081 4644
rect 6115 4641 6127 4675
rect 6069 4635 6127 4641
rect 7300 4616 7328 4712
rect 7374 4700 7380 4752
rect 7432 4740 7438 4752
rect 9490 4749 9496 4752
rect 7530 4743 7588 4749
rect 7530 4740 7542 4743
rect 7432 4712 7542 4740
rect 7432 4700 7438 4712
rect 7530 4709 7542 4712
rect 7576 4709 7588 4743
rect 9484 4740 9496 4749
rect 9451 4712 9496 4740
rect 7530 4703 7588 4709
rect 9484 4703 9496 4712
rect 9490 4700 9496 4703
rect 9548 4700 9554 4752
rect 10686 4700 10692 4752
rect 10744 4740 10750 4752
rect 11241 4743 11299 4749
rect 11241 4740 11253 4743
rect 10744 4712 11253 4740
rect 10744 4700 10750 4712
rect 11241 4709 11253 4712
rect 11287 4709 11299 4743
rect 11701 4743 11759 4749
rect 11701 4740 11713 4743
rect 11241 4703 11299 4709
rect 11624 4712 11713 4740
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 11624 4672 11652 4712
rect 11701 4709 11713 4712
rect 11747 4709 11759 4743
rect 11701 4703 11759 4709
rect 11808 4684 11836 4780
rect 12066 4768 12072 4820
rect 12124 4768 12130 4820
rect 13262 4808 13268 4820
rect 13162 4780 13268 4808
rect 11931 4709 11989 4715
rect 11931 4706 11943 4709
rect 9180 4644 11652 4672
rect 9180 4632 9186 4644
rect 11790 4632 11796 4684
rect 11848 4672 11854 4684
rect 11926 4675 11943 4706
rect 11977 4675 11989 4709
rect 12158 4700 12164 4752
rect 12216 4700 12222 4752
rect 13162 4749 13190 4780
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 13630 4768 13636 4820
rect 13688 4768 13694 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13872 4780 14105 4808
rect 13872 4768 13878 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14093 4771 14151 4777
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14829 4811 14887 4817
rect 14829 4808 14841 4811
rect 14240 4780 14841 4808
rect 14240 4768 14246 4780
rect 14829 4777 14841 4780
rect 14875 4777 14887 4811
rect 14829 4771 14887 4777
rect 14992 4811 15050 4817
rect 14992 4777 15004 4811
rect 15038 4808 15050 4811
rect 15038 4780 16252 4808
rect 15038 4777 15050 4780
rect 14992 4771 15050 4777
rect 12377 4743 12435 4749
rect 12377 4740 12389 4743
rect 12376 4709 12389 4740
rect 12423 4709 12435 4743
rect 12376 4703 12435 4709
rect 13147 4743 13205 4749
rect 13147 4709 13159 4743
rect 13193 4709 13205 4743
rect 13147 4703 13205 4709
rect 13357 4743 13415 4749
rect 13357 4709 13369 4743
rect 13403 4709 13415 4743
rect 13725 4743 13783 4749
rect 13725 4740 13737 4743
rect 13357 4703 13415 4709
rect 13664 4712 13737 4740
rect 11926 4672 11989 4675
rect 12376 4672 12404 4703
rect 11848 4644 12404 4672
rect 13265 4675 13323 4681
rect 11848 4632 11854 4644
rect 13265 4641 13277 4675
rect 13311 4641 13323 4675
rect 13265 4635 13323 4641
rect 4540 4576 5948 4604
rect 952 4508 2084 4536
rect 3344 4508 3556 4536
rect 952 4480 980 4508
rect 934 4428 940 4480
rect 992 4428 998 4480
rect 1486 4428 1492 4480
rect 1544 4468 1550 4480
rect 3344 4468 3372 4508
rect 1544 4440 3372 4468
rect 1544 4428 1550 4440
rect 3418 4428 3424 4480
rect 3476 4428 3482 4480
rect 3528 4468 3556 4508
rect 4540 4468 4568 4576
rect 7282 4564 7288 4616
rect 7340 4564 7346 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4573 13047 4607
rect 12989 4567 13047 4573
rect 4890 4496 4896 4548
rect 4948 4496 4954 4548
rect 3528 4440 4568 4468
rect 9232 4468 9260 4567
rect 10597 4539 10655 4545
rect 10597 4505 10609 4539
rect 10643 4536 10655 4539
rect 10643 4508 11560 4536
rect 10643 4505 10655 4508
rect 10597 4499 10655 4505
rect 9398 4468 9404 4480
rect 9232 4440 9404 4468
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 11422 4428 11428 4480
rect 11480 4428 11486 4480
rect 11532 4468 11560 4508
rect 11606 4496 11612 4548
rect 11664 4496 11670 4548
rect 13004 4536 13032 4567
rect 13078 4564 13084 4616
rect 13136 4604 13142 4616
rect 13280 4604 13308 4635
rect 13372 4616 13400 4703
rect 13664 4684 13692 4712
rect 13725 4709 13737 4712
rect 13771 4709 13783 4743
rect 13725 4703 13783 4709
rect 13941 4743 13999 4749
rect 13941 4709 13953 4743
rect 13987 4740 13999 4743
rect 13987 4712 14688 4740
rect 13987 4709 13999 4712
rect 13941 4703 13999 4709
rect 13446 4632 13452 4684
rect 13504 4632 13510 4684
rect 13630 4632 13636 4684
rect 13688 4632 13694 4684
rect 14274 4632 14280 4684
rect 14332 4632 14338 4684
rect 13136 4576 13308 4604
rect 13136 4564 13142 4576
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 14292 4604 14320 4632
rect 14660 4616 14688 4712
rect 14734 4700 14740 4752
rect 14792 4740 14798 4752
rect 15012 4740 15040 4771
rect 14792 4712 15040 4740
rect 15197 4743 15255 4749
rect 14792 4700 14798 4712
rect 15197 4709 15209 4743
rect 15243 4740 15255 4743
rect 15378 4740 15384 4752
rect 15243 4712 15384 4740
rect 15243 4709 15255 4712
rect 15197 4703 15255 4709
rect 15378 4700 15384 4712
rect 15436 4700 15442 4752
rect 15654 4700 15660 4752
rect 15712 4700 15718 4752
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 14844 4644 15485 4672
rect 14844 4616 14872 4644
rect 15473 4641 15485 4644
rect 15519 4672 15531 4675
rect 15672 4672 15700 4700
rect 15519 4644 15700 4672
rect 15519 4641 15531 4644
rect 15473 4635 15531 4641
rect 13412 4576 14320 4604
rect 13412 4564 13418 4576
rect 14642 4564 14648 4616
rect 14700 4564 14706 4616
rect 14826 4564 14832 4616
rect 14884 4564 14890 4616
rect 15194 4564 15200 4616
rect 15252 4604 15258 4616
rect 15289 4607 15347 4613
rect 15289 4604 15301 4607
rect 15252 4576 15301 4604
rect 15252 4564 15258 4576
rect 15289 4573 15301 4576
rect 15335 4573 15347 4607
rect 16224 4604 16252 4780
rect 16298 4768 16304 4820
rect 16356 4808 16362 4820
rect 16356 4780 17908 4808
rect 16356 4768 16362 4780
rect 16669 4743 16727 4749
rect 16669 4709 16681 4743
rect 16715 4740 16727 4743
rect 16758 4740 16764 4752
rect 16715 4712 16764 4740
rect 16715 4709 16727 4712
rect 16669 4703 16727 4709
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 17880 4740 17908 4780
rect 18598 4768 18604 4820
rect 18656 4768 18662 4820
rect 18966 4768 18972 4820
rect 19024 4768 19030 4820
rect 19150 4768 19156 4820
rect 19208 4768 19214 4820
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 19613 4811 19671 4817
rect 19613 4808 19625 4811
rect 19484 4780 19625 4808
rect 19484 4768 19490 4780
rect 19613 4777 19625 4780
rect 19659 4777 19671 4811
rect 19613 4771 19671 4777
rect 20162 4768 20168 4820
rect 20220 4808 20226 4820
rect 20349 4811 20407 4817
rect 20349 4808 20361 4811
rect 20220 4780 20361 4808
rect 20220 4768 20226 4780
rect 20349 4777 20361 4780
rect 20395 4777 20407 4811
rect 20349 4771 20407 4777
rect 20993 4811 21051 4817
rect 20993 4777 21005 4811
rect 21039 4808 21051 4811
rect 21039 4780 22885 4808
rect 21039 4777 21051 4780
rect 20993 4771 21051 4777
rect 19168 4740 19196 4768
rect 17880 4712 18920 4740
rect 19168 4712 20116 4740
rect 16776 4672 16804 4700
rect 17880 4681 17908 4712
rect 17129 4675 17187 4681
rect 17129 4672 17141 4675
rect 16776 4644 17141 4672
rect 17129 4641 17141 4644
rect 17175 4672 17187 4675
rect 17313 4675 17371 4681
rect 17313 4672 17325 4675
rect 17175 4644 17325 4672
rect 17175 4641 17187 4644
rect 17129 4635 17187 4641
rect 17313 4641 17325 4644
rect 17359 4641 17371 4675
rect 17313 4635 17371 4641
rect 17865 4675 17923 4681
rect 17865 4641 17877 4675
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 18046 4632 18052 4684
rect 18104 4632 18110 4684
rect 18141 4675 18199 4681
rect 18141 4641 18153 4675
rect 18187 4672 18199 4675
rect 18690 4672 18696 4684
rect 18187 4644 18696 4672
rect 18187 4641 18199 4644
rect 18141 4635 18199 4641
rect 18690 4632 18696 4644
rect 18748 4632 18754 4684
rect 18892 4681 18920 4712
rect 18877 4675 18935 4681
rect 18877 4641 18889 4675
rect 18923 4641 18935 4675
rect 18877 4635 18935 4641
rect 19153 4675 19211 4681
rect 19153 4641 19165 4675
rect 19199 4672 19211 4675
rect 19334 4672 19340 4684
rect 19199 4644 19340 4672
rect 19199 4641 19211 4644
rect 19153 4635 19211 4641
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 20088 4681 20116 4712
rect 20254 4700 20260 4752
rect 20312 4700 20318 4752
rect 21904 4743 21962 4749
rect 20364 4712 21864 4740
rect 20364 4684 20392 4712
rect 20073 4675 20131 4681
rect 20073 4641 20085 4675
rect 20119 4672 20131 4675
rect 20119 4644 20300 4672
rect 20119 4641 20131 4644
rect 20073 4635 20131 4641
rect 20272 4616 20300 4644
rect 20346 4632 20352 4684
rect 20404 4632 20410 4684
rect 21082 4632 21088 4684
rect 21140 4632 21146 4684
rect 21358 4632 21364 4684
rect 21416 4672 21422 4684
rect 21637 4675 21695 4681
rect 21637 4672 21649 4675
rect 21416 4644 21649 4672
rect 21416 4632 21422 4644
rect 21637 4641 21649 4644
rect 21683 4641 21695 4675
rect 21836 4672 21864 4712
rect 21904 4709 21916 4743
rect 21950 4740 21962 4743
rect 22186 4740 22192 4752
rect 21950 4712 22192 4740
rect 21950 4709 21962 4712
rect 21904 4703 21962 4709
rect 22186 4700 22192 4712
rect 22244 4700 22250 4752
rect 22857 4740 22885 4780
rect 23014 4768 23020 4820
rect 23072 4768 23078 4820
rect 23106 4768 23112 4820
rect 23164 4808 23170 4820
rect 29457 4811 29515 4817
rect 29457 4808 29469 4811
rect 23164 4780 29469 4808
rect 23164 4768 23170 4780
rect 29457 4777 29469 4780
rect 29503 4777 29515 4811
rect 29457 4771 29515 4777
rect 28258 4740 28264 4752
rect 22857 4712 28264 4740
rect 28258 4700 28264 4712
rect 28316 4700 28322 4752
rect 28718 4700 28724 4752
rect 28776 4740 28782 4752
rect 28776 4712 29040 4740
rect 28776 4700 28782 4712
rect 24762 4672 24768 4684
rect 21836 4644 24768 4672
rect 21637 4635 21695 4641
rect 24762 4632 24768 4644
rect 24820 4632 24826 4684
rect 27706 4632 27712 4684
rect 27764 4681 27770 4684
rect 27764 4635 27776 4681
rect 27764 4632 27770 4635
rect 28902 4632 28908 4684
rect 28960 4632 28966 4684
rect 29012 4681 29040 4712
rect 29086 4700 29092 4752
rect 29144 4700 29150 4752
rect 28997 4675 29055 4681
rect 28997 4641 29009 4675
rect 29043 4641 29055 4675
rect 28997 4635 29055 4641
rect 30558 4632 30564 4684
rect 30616 4681 30622 4684
rect 30616 4635 30628 4681
rect 30616 4632 30622 4635
rect 30742 4632 30748 4684
rect 30800 4672 30806 4684
rect 30837 4675 30895 4681
rect 30837 4672 30849 4675
rect 30800 4644 30849 4672
rect 30800 4632 30806 4644
rect 30837 4641 30849 4644
rect 30883 4641 30895 4675
rect 30837 4635 30895 4641
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 16224 4576 17509 4604
rect 15289 4567 15347 4573
rect 17497 4573 17509 4576
rect 17543 4604 17555 4607
rect 19889 4607 19947 4613
rect 19889 4604 19901 4607
rect 17543 4576 19901 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 19889 4573 19901 4576
rect 19935 4604 19947 4607
rect 20162 4604 20168 4616
rect 19935 4576 20168 4604
rect 19935 4573 19947 4576
rect 19889 4567 19947 4573
rect 20162 4564 20168 4576
rect 20220 4564 20226 4616
rect 20254 4564 20260 4616
rect 20312 4564 20318 4616
rect 27982 4564 27988 4616
rect 28040 4564 28046 4616
rect 28813 4607 28871 4613
rect 28813 4573 28825 4607
rect 28859 4604 28871 4607
rect 29822 4604 29828 4616
rect 28859 4576 29828 4604
rect 28859 4573 28871 4576
rect 28813 4567 28871 4573
rect 29822 4564 29828 4576
rect 29880 4564 29886 4616
rect 18233 4539 18291 4545
rect 18233 4536 18245 4539
rect 11716 4508 13032 4536
rect 13832 4508 18245 4536
rect 11716 4468 11744 4508
rect 11532 4440 11744 4468
rect 11885 4471 11943 4477
rect 11885 4437 11897 4471
rect 11931 4468 11943 4471
rect 11974 4468 11980 4480
rect 11931 4440 11980 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 11974 4428 11980 4440
rect 12032 4468 12038 4480
rect 12345 4471 12403 4477
rect 12345 4468 12357 4471
rect 12032 4440 12357 4468
rect 12032 4428 12038 4440
rect 12345 4437 12357 4440
rect 12391 4437 12403 4471
rect 12345 4431 12403 4437
rect 12529 4471 12587 4477
rect 12529 4437 12541 4471
rect 12575 4468 12587 4471
rect 13832 4468 13860 4508
rect 18233 4505 18245 4508
rect 18279 4505 18291 4539
rect 18233 4499 18291 4505
rect 19978 4496 19984 4548
rect 20036 4536 20042 4548
rect 20036 4508 20944 4536
rect 20036 4496 20042 4508
rect 12575 4440 13860 4468
rect 13909 4471 13967 4477
rect 12575 4437 12587 4440
rect 12529 4431 12587 4437
rect 13909 4437 13921 4471
rect 13955 4468 13967 4471
rect 13998 4468 14004 4480
rect 13955 4440 14004 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 15013 4471 15071 4477
rect 15013 4437 15025 4471
rect 15059 4468 15071 4471
rect 15470 4468 15476 4480
rect 15059 4440 15476 4468
rect 15059 4437 15071 4440
rect 15013 4431 15071 4437
rect 15470 4428 15476 4440
rect 15528 4428 15534 4480
rect 15657 4471 15715 4477
rect 15657 4437 15669 4471
rect 15703 4468 15715 4471
rect 15838 4468 15844 4480
rect 15703 4440 15844 4468
rect 15703 4437 15715 4440
rect 15657 4431 15715 4437
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 16482 4428 16488 4480
rect 16540 4468 16546 4480
rect 16577 4471 16635 4477
rect 16577 4468 16589 4471
rect 16540 4440 16589 4468
rect 16540 4428 16546 4440
rect 16577 4437 16589 4440
rect 16623 4437 16635 4471
rect 16577 4431 16635 4437
rect 16942 4428 16948 4480
rect 17000 4428 17006 4480
rect 18322 4428 18328 4480
rect 18380 4428 18386 4480
rect 18414 4428 18420 4480
rect 18472 4468 18478 4480
rect 19245 4471 19303 4477
rect 19245 4468 19257 4471
rect 18472 4440 19257 4468
rect 18472 4428 18478 4440
rect 19245 4437 19257 4440
rect 19291 4437 19303 4471
rect 19245 4431 19303 4437
rect 19334 4428 19340 4480
rect 19392 4428 19398 4480
rect 20622 4428 20628 4480
rect 20680 4428 20686 4480
rect 20714 4428 20720 4480
rect 20772 4428 20778 4480
rect 20806 4428 20812 4480
rect 20864 4428 20870 4480
rect 20916 4468 20944 4508
rect 26605 4471 26663 4477
rect 26605 4468 26617 4471
rect 20916 4440 26617 4468
rect 26605 4437 26617 4440
rect 26651 4437 26663 4471
rect 26605 4431 26663 4437
rect 552 4378 31372 4400
rect 552 4326 4250 4378
rect 4302 4326 4314 4378
rect 4366 4326 4378 4378
rect 4430 4326 4442 4378
rect 4494 4326 4506 4378
rect 4558 4326 11955 4378
rect 12007 4326 12019 4378
rect 12071 4326 12083 4378
rect 12135 4326 12147 4378
rect 12199 4326 12211 4378
rect 12263 4326 19660 4378
rect 19712 4326 19724 4378
rect 19776 4326 19788 4378
rect 19840 4326 19852 4378
rect 19904 4326 19916 4378
rect 19968 4326 27365 4378
rect 27417 4326 27429 4378
rect 27481 4326 27493 4378
rect 27545 4326 27557 4378
rect 27609 4326 27621 4378
rect 27673 4326 31372 4378
rect 552 4304 31372 4326
rect 1210 4224 1216 4276
rect 1268 4224 1274 4276
rect 1486 4224 1492 4276
rect 1544 4264 1550 4276
rect 2041 4267 2099 4273
rect 2041 4264 2053 4267
rect 1544 4236 2053 4264
rect 1544 4224 1550 4236
rect 2041 4233 2053 4236
rect 2087 4233 2099 4267
rect 2041 4227 2099 4233
rect 1228 4196 1256 4224
rect 1765 4199 1823 4205
rect 1765 4196 1777 4199
rect 1228 4168 1777 4196
rect 1765 4165 1777 4168
rect 1811 4196 1823 4199
rect 1946 4196 1952 4208
rect 1811 4168 1952 4196
rect 1811 4165 1823 4168
rect 1765 4159 1823 4165
rect 1946 4156 1952 4168
rect 2004 4156 2010 4208
rect 2056 4128 2084 4227
rect 3418 4224 3424 4276
rect 3476 4264 3482 4276
rect 3476 4236 11468 4264
rect 3476 4224 3482 4236
rect 10965 4199 11023 4205
rect 10965 4165 10977 4199
rect 11011 4165 11023 4199
rect 11440 4196 11468 4236
rect 11514 4224 11520 4276
rect 11572 4264 11578 4276
rect 11701 4267 11759 4273
rect 11701 4264 11713 4267
rect 11572 4236 11713 4264
rect 11572 4224 11578 4236
rect 11701 4233 11713 4236
rect 11747 4264 11759 4267
rect 11882 4264 11888 4276
rect 11747 4236 11888 4264
rect 11747 4233 11759 4236
rect 11701 4227 11759 4233
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 13630 4224 13636 4276
rect 13688 4224 13694 4276
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 14461 4267 14519 4273
rect 14461 4264 14473 4267
rect 14056 4236 14473 4264
rect 14056 4224 14062 4236
rect 14461 4233 14473 4236
rect 14507 4264 14519 4267
rect 14826 4264 14832 4276
rect 14507 4236 14832 4264
rect 14507 4233 14519 4236
rect 14461 4227 14519 4233
rect 14826 4224 14832 4236
rect 14884 4224 14890 4276
rect 15096 4267 15154 4273
rect 15096 4233 15108 4267
rect 15142 4264 15154 4267
rect 15194 4264 15200 4276
rect 15142 4236 15200 4264
rect 15142 4233 15154 4236
rect 15096 4227 15154 4233
rect 15194 4224 15200 4236
rect 15252 4224 15258 4276
rect 15286 4224 15292 4276
rect 15344 4224 15350 4276
rect 15565 4267 15623 4273
rect 15565 4233 15577 4267
rect 15611 4264 15623 4267
rect 15654 4264 15660 4276
rect 15611 4236 15660 4264
rect 15611 4233 15623 4236
rect 15565 4227 15623 4233
rect 15654 4224 15660 4236
rect 15712 4224 15718 4276
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 16758 4264 16764 4276
rect 16632 4236 16764 4264
rect 16632 4224 16638 4236
rect 16758 4224 16764 4236
rect 16816 4224 16822 4276
rect 17402 4224 17408 4276
rect 17460 4264 17466 4276
rect 17773 4267 17831 4273
rect 17773 4264 17785 4267
rect 17460 4236 17785 4264
rect 17460 4224 17466 4236
rect 17773 4233 17785 4236
rect 17819 4233 17831 4267
rect 17773 4227 17831 4233
rect 18046 4224 18052 4276
rect 18104 4224 18110 4276
rect 18233 4267 18291 4273
rect 18233 4233 18245 4267
rect 18279 4264 18291 4267
rect 18322 4264 18328 4276
rect 18279 4236 18328 4264
rect 18279 4233 18291 4236
rect 18233 4227 18291 4233
rect 18322 4224 18328 4236
rect 18380 4224 18386 4276
rect 20073 4267 20131 4273
rect 20073 4233 20085 4267
rect 20119 4264 20131 4267
rect 20162 4264 20168 4276
rect 20119 4236 20168 4264
rect 20119 4233 20131 4236
rect 20073 4227 20131 4233
rect 20162 4224 20168 4236
rect 20220 4224 20226 4276
rect 20254 4224 20260 4276
rect 20312 4224 20318 4276
rect 20714 4224 20720 4276
rect 20772 4264 20778 4276
rect 21545 4267 21603 4273
rect 21545 4264 21557 4267
rect 20772 4236 21557 4264
rect 20772 4224 20778 4236
rect 21545 4233 21557 4236
rect 21591 4233 21603 4267
rect 21545 4227 21603 4233
rect 21726 4224 21732 4276
rect 21784 4264 21790 4276
rect 22646 4264 22652 4276
rect 21784 4236 22652 4264
rect 21784 4224 21790 4236
rect 22646 4224 22652 4236
rect 22704 4224 22710 4276
rect 22741 4267 22799 4273
rect 22741 4233 22753 4267
rect 22787 4233 22799 4267
rect 22741 4227 22799 4233
rect 13648 4196 13676 4224
rect 11440 4168 13676 4196
rect 10965 4159 11023 4165
rect 2314 4128 2320 4140
rect 2056 4100 2320 4128
rect 2314 4088 2320 4100
rect 2372 4128 2378 4140
rect 2372 4100 2728 4128
rect 2372 4088 2378 4100
rect 934 4020 940 4072
rect 992 4060 998 4072
rect 1489 4063 1547 4069
rect 1489 4060 1501 4063
rect 992 4032 1501 4060
rect 992 4020 998 4032
rect 1489 4029 1501 4032
rect 1535 4029 1547 4063
rect 1489 4023 1547 4029
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4029 1639 4063
rect 1581 4023 1639 4029
rect 1596 3924 1624 4023
rect 1854 4020 1860 4072
rect 1912 4020 1918 4072
rect 1946 4020 1952 4072
rect 2004 4020 2010 4072
rect 2222 4020 2228 4072
rect 2280 4020 2286 4072
rect 2700 4069 2728 4100
rect 9324 4100 9720 4128
rect 9324 4072 9352 4100
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4029 2743 4063
rect 2685 4023 2743 4029
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 3568 4032 3617 4060
rect 3568 4020 3574 4032
rect 3605 4029 3617 4032
rect 3651 4060 3663 4063
rect 5629 4063 5687 4069
rect 5629 4060 5641 4063
rect 3651 4032 5641 4060
rect 3651 4029 3663 4032
rect 3605 4023 3663 4029
rect 5629 4029 5641 4032
rect 5675 4060 5687 4063
rect 7282 4060 7288 4072
rect 5675 4032 7288 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 9306 4020 9312 4072
rect 9364 4020 9370 4072
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9585 4063 9643 4069
rect 9585 4060 9597 4063
rect 9456 4032 9597 4060
rect 9456 4020 9462 4032
rect 9585 4029 9597 4032
rect 9631 4029 9643 4063
rect 9692 4060 9720 4100
rect 10686 4088 10692 4140
rect 10744 4088 10750 4140
rect 10980 4128 11008 4159
rect 14366 4156 14372 4208
rect 14424 4196 14430 4208
rect 14645 4199 14703 4205
rect 14645 4196 14657 4199
rect 14424 4168 14657 4196
rect 14424 4156 14430 4168
rect 14645 4165 14657 4168
rect 14691 4165 14703 4199
rect 14645 4159 14703 4165
rect 15749 4199 15807 4205
rect 15749 4165 15761 4199
rect 15795 4196 15807 4199
rect 17313 4199 17371 4205
rect 17313 4196 17325 4199
rect 15795 4168 17325 4196
rect 15795 4165 15807 4168
rect 15749 4159 15807 4165
rect 17313 4165 17325 4168
rect 17359 4165 17371 4199
rect 17313 4159 17371 4165
rect 19889 4199 19947 4205
rect 19889 4165 19901 4199
rect 19935 4196 19947 4199
rect 19935 4168 20116 4196
rect 19935 4165 19947 4168
rect 19889 4159 19947 4165
rect 20088 4140 20116 4168
rect 17405 4131 17463 4137
rect 10980 4100 17264 4128
rect 9841 4063 9899 4069
rect 9841 4060 9853 4063
rect 9692 4032 9853 4060
rect 9585 4023 9643 4029
rect 9841 4029 9853 4032
rect 9887 4029 9899 4063
rect 9841 4023 9899 4029
rect 2498 3952 2504 4004
rect 2556 3992 2562 4004
rect 3850 3995 3908 4001
rect 3850 3992 3862 3995
rect 2556 3964 3862 3992
rect 2556 3952 2562 3964
rect 3850 3961 3862 3964
rect 3896 3961 3908 3995
rect 3850 3955 3908 3961
rect 5442 3952 5448 4004
rect 5500 3992 5506 4004
rect 5874 3995 5932 4001
rect 5874 3992 5886 3995
rect 5500 3964 5886 3992
rect 5500 3952 5506 3964
rect 5874 3961 5886 3964
rect 5920 3961 5932 3995
rect 10704 3992 10732 4088
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 11388 4032 14780 4060
rect 11388 4020 11394 4032
rect 5874 3955 5932 3961
rect 6932 3964 10732 3992
rect 2038 3924 2044 3936
rect 1596 3896 2044 3924
rect 2038 3884 2044 3896
rect 2096 3924 2102 3936
rect 2317 3927 2375 3933
rect 2317 3924 2329 3927
rect 2096 3896 2329 3924
rect 2096 3884 2102 3896
rect 2317 3893 2329 3896
rect 2363 3924 2375 3927
rect 2593 3927 2651 3933
rect 2593 3924 2605 3927
rect 2363 3896 2605 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 2593 3893 2605 3896
rect 2639 3893 2651 3927
rect 2593 3887 2651 3893
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 6932 3924 6960 3964
rect 11514 3952 11520 4004
rect 11572 3952 11578 4004
rect 11790 4001 11796 4004
rect 11733 3995 11796 4001
rect 11733 3961 11745 3995
rect 11779 3961 11796 3995
rect 11733 3955 11796 3961
rect 11790 3952 11796 3955
rect 11848 3992 11854 4004
rect 12526 3992 12532 4004
rect 11848 3964 12532 3992
rect 11848 3952 11854 3964
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 12676 3964 13952 3992
rect 12676 3952 12682 3964
rect 5031 3896 6960 3924
rect 7009 3927 7067 3933
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 7009 3893 7021 3927
rect 7055 3924 7067 3927
rect 9122 3924 9128 3936
rect 7055 3896 9128 3924
rect 7055 3893 7067 3896
rect 7009 3887 7067 3893
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 11885 3927 11943 3933
rect 11885 3893 11897 3927
rect 11931 3924 11943 3927
rect 13814 3924 13820 3936
rect 11931 3896 13820 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 13924 3924 13952 3964
rect 14274 3952 14280 4004
rect 14332 3952 14338 4004
rect 14493 3995 14551 4001
rect 14493 3961 14505 3995
rect 14539 3992 14551 3995
rect 14642 3992 14648 4004
rect 14539 3964 14648 3992
rect 14539 3961 14551 3964
rect 14493 3955 14551 3961
rect 14642 3952 14648 3964
rect 14700 3952 14706 4004
rect 14752 3992 14780 4032
rect 14826 4020 14832 4072
rect 14884 4060 14890 4072
rect 14884 4032 15164 4060
rect 14884 4020 14890 4032
rect 15136 4001 15164 4032
rect 15562 4020 15568 4072
rect 15620 4020 15626 4072
rect 15838 4020 15844 4072
rect 15896 4060 15902 4072
rect 17236 4069 17264 4100
rect 17405 4097 17417 4131
rect 17451 4128 17463 4131
rect 19610 4128 19616 4140
rect 17451 4100 19616 4128
rect 17451 4097 17463 4100
rect 17405 4091 17463 4097
rect 19610 4088 19616 4100
rect 19668 4088 19674 4140
rect 20070 4088 20076 4140
rect 20128 4088 20134 4140
rect 17037 4063 17095 4069
rect 17037 4060 17049 4063
rect 15896 4032 17049 4060
rect 15896 4020 15902 4032
rect 17037 4029 17049 4032
rect 17083 4029 17095 4063
rect 17037 4023 17095 4029
rect 17221 4063 17279 4069
rect 17221 4029 17233 4063
rect 17267 4029 17279 4063
rect 17221 4023 17279 4029
rect 17494 4020 17500 4072
rect 17552 4020 17558 4072
rect 20272 4060 20300 4224
rect 22756 4196 22784 4227
rect 22830 4224 22836 4276
rect 22888 4224 22894 4276
rect 22922 4224 22928 4276
rect 22980 4264 22986 4276
rect 23017 4267 23075 4273
rect 23017 4264 23029 4267
rect 22980 4236 23029 4264
rect 22980 4224 22986 4236
rect 23017 4233 23029 4236
rect 23063 4233 23075 4267
rect 23017 4227 23075 4233
rect 23106 4224 23112 4276
rect 23164 4264 23170 4276
rect 23201 4267 23259 4273
rect 23201 4264 23213 4267
rect 23164 4236 23213 4264
rect 23164 4224 23170 4236
rect 23201 4233 23213 4236
rect 23247 4233 23259 4267
rect 24029 4267 24087 4273
rect 24029 4264 24041 4267
rect 23201 4227 23259 4233
rect 23308 4236 24041 4264
rect 22664 4168 22784 4196
rect 22848 4196 22876 4224
rect 23308 4196 23336 4236
rect 24029 4233 24041 4236
rect 24075 4233 24087 4267
rect 24029 4227 24087 4233
rect 24118 4224 24124 4276
rect 24176 4264 24182 4276
rect 24305 4267 24363 4273
rect 24305 4264 24317 4267
rect 24176 4236 24317 4264
rect 24176 4224 24182 4236
rect 24305 4233 24317 4236
rect 24351 4233 24363 4267
rect 24489 4267 24547 4273
rect 24489 4264 24501 4267
rect 24305 4227 24363 4233
rect 24412 4236 24501 4264
rect 22848 4168 23336 4196
rect 23845 4199 23903 4205
rect 22664 4140 22692 4168
rect 23845 4165 23857 4199
rect 23891 4196 23903 4199
rect 23891 4168 24072 4196
rect 23891 4165 23903 4168
rect 23845 4159 23903 4165
rect 24044 4140 24072 4168
rect 22646 4088 22652 4140
rect 22704 4088 22710 4140
rect 23106 4088 23112 4140
rect 23164 4088 23170 4140
rect 24026 4088 24032 4140
rect 24084 4088 24090 4140
rect 20349 4063 20407 4069
rect 20349 4060 20361 4063
rect 17788 4032 20024 4060
rect 20272 4032 20361 4060
rect 14921 3995 14979 4001
rect 14921 3992 14933 3995
rect 14752 3964 14933 3992
rect 14921 3961 14933 3964
rect 14967 3961 14979 3995
rect 14921 3955 14979 3961
rect 15121 3995 15179 4001
rect 15121 3961 15133 3995
rect 15167 3961 15179 3995
rect 15381 3995 15439 4001
rect 15381 3992 15393 3995
rect 15121 3955 15179 3961
rect 15212 3964 15393 3992
rect 15212 3924 15240 3964
rect 15381 3961 15393 3964
rect 15427 3961 15439 3995
rect 15381 3955 15439 3961
rect 15580 3992 15608 4020
rect 16850 3992 16856 4004
rect 15580 3964 16856 3992
rect 13924 3896 15240 3924
rect 15580 3933 15608 3964
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 16942 3952 16948 4004
rect 17000 3952 17006 4004
rect 17310 3952 17316 4004
rect 17368 3992 17374 4004
rect 17788 3992 17816 4032
rect 17368 3964 17816 3992
rect 17865 3995 17923 4001
rect 17368 3952 17374 3964
rect 17865 3961 17877 3995
rect 17911 3992 17923 3995
rect 17954 3992 17960 4004
rect 17911 3964 17960 3992
rect 17911 3961 17923 3964
rect 17865 3955 17923 3961
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 19996 3992 20024 4032
rect 20349 4029 20361 4032
rect 20395 4029 20407 4063
rect 23124 4060 23152 4088
rect 20349 4023 20407 4029
rect 21551 4032 22508 4060
rect 20052 3995 20110 4001
rect 20052 3992 20064 3995
rect 19996 3964 20064 3992
rect 20052 3961 20064 3964
rect 20098 3992 20110 3995
rect 20257 3995 20315 4001
rect 20098 3964 20208 3992
rect 20098 3961 20110 3964
rect 20052 3955 20110 3961
rect 15580 3927 15639 3933
rect 15580 3896 15593 3927
rect 15581 3893 15593 3896
rect 15627 3893 15639 3927
rect 15581 3887 15639 3893
rect 16574 3884 16580 3936
rect 16632 3884 16638 3936
rect 16745 3927 16803 3933
rect 16745 3893 16757 3927
rect 16791 3924 16803 3927
rect 17034 3924 17040 3936
rect 16791 3896 17040 3924
rect 16791 3893 16803 3896
rect 16745 3887 16803 3893
rect 17034 3884 17040 3896
rect 17092 3924 17098 3936
rect 18065 3927 18123 3933
rect 18065 3924 18077 3927
rect 17092 3896 18077 3924
rect 17092 3884 17098 3896
rect 18065 3893 18077 3896
rect 18111 3893 18123 3927
rect 20180 3924 20208 3964
rect 20257 3961 20269 3995
rect 20303 3992 20315 3995
rect 21450 3992 21456 4004
rect 20303 3964 21456 3992
rect 20303 3961 20315 3964
rect 20257 3955 20315 3961
rect 21450 3952 21456 3964
rect 21508 3952 21514 4004
rect 20533 3927 20591 3933
rect 20533 3924 20545 3927
rect 20180 3896 20545 3924
rect 18065 3887 18123 3893
rect 20533 3893 20545 3896
rect 20579 3924 20591 3927
rect 21551 3924 21579 4032
rect 22480 4026 22508 4032
rect 22695 4029 22753 4035
rect 23124 4032 23519 4060
rect 22695 4026 22707 4029
rect 21913 3995 21971 4001
rect 21913 3961 21925 3995
rect 21959 3992 21971 3995
rect 22370 3992 22376 4004
rect 21959 3964 22376 3992
rect 21959 3961 21971 3964
rect 21913 3955 21971 3961
rect 22370 3952 22376 3964
rect 22428 3952 22434 4004
rect 22480 3998 22707 4026
rect 22695 3995 22707 3998
rect 22741 4026 22753 4029
rect 22741 3995 22768 4026
rect 22695 3989 22768 3995
rect 20579 3896 21579 3924
rect 21713 3927 21771 3933
rect 20579 3893 20591 3896
rect 20533 3887 20591 3893
rect 21713 3893 21725 3927
rect 21759 3924 21771 3927
rect 21818 3924 21824 3936
rect 21759 3896 21824 3924
rect 21759 3893 21771 3896
rect 21713 3887 21771 3893
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 22554 3884 22560 3936
rect 22612 3884 22618 3936
rect 22740 3924 22768 3989
rect 22922 3952 22928 4004
rect 22980 3952 22986 4004
rect 23290 3952 23296 4004
rect 23348 3992 23354 4004
rect 23385 3995 23443 4001
rect 23385 3992 23397 3995
rect 23348 3964 23397 3992
rect 23348 3952 23354 3964
rect 23385 3961 23397 3964
rect 23431 3961 23443 3995
rect 23385 3955 23443 3961
rect 23198 3933 23204 3936
rect 23175 3927 23204 3933
rect 23175 3924 23187 3927
rect 22740 3896 23187 3924
rect 23175 3893 23187 3896
rect 23175 3887 23204 3893
rect 23198 3884 23204 3887
rect 23256 3884 23262 3936
rect 23491 3924 23519 4032
rect 23934 4020 23940 4072
rect 23992 4060 23998 4072
rect 23992 4032 24256 4060
rect 23992 4020 23998 4032
rect 24228 4001 24256 4032
rect 24213 3995 24271 4001
rect 24213 3961 24225 3995
rect 24259 3961 24271 3995
rect 24213 3955 24271 3961
rect 24003 3927 24061 3933
rect 24003 3924 24015 3927
rect 23491 3896 24015 3924
rect 24003 3893 24015 3896
rect 24049 3924 24061 3927
rect 24412 3924 24440 4236
rect 24489 4233 24501 4236
rect 24535 4233 24547 4267
rect 24489 4227 24547 4233
rect 24762 4224 24768 4276
rect 24820 4224 24826 4276
rect 29822 4224 29828 4276
rect 29880 4264 29886 4276
rect 30745 4267 30803 4273
rect 30745 4264 30757 4267
rect 29880 4236 30757 4264
rect 29880 4224 29886 4236
rect 30745 4233 30757 4236
rect 30791 4233 30803 4267
rect 30745 4227 30803 4233
rect 29365 4199 29423 4205
rect 29365 4165 29377 4199
rect 29411 4196 29423 4199
rect 30193 4199 30251 4205
rect 30193 4196 30205 4199
rect 29411 4168 30205 4196
rect 29411 4165 29423 4168
rect 29365 4159 29423 4165
rect 30193 4165 30205 4168
rect 30239 4165 30251 4199
rect 30193 4159 30251 4165
rect 30208 4128 30236 4159
rect 30558 4128 30564 4140
rect 28276 4100 29592 4128
rect 26050 4020 26056 4072
rect 26108 4060 26114 4072
rect 26145 4063 26203 4069
rect 26145 4060 26157 4063
rect 26108 4032 26157 4060
rect 26108 4020 26114 4032
rect 26145 4029 26157 4032
rect 26191 4060 26203 4063
rect 27982 4060 27988 4072
rect 26191 4032 27988 4060
rect 26191 4029 26203 4032
rect 26145 4023 26203 4029
rect 27982 4020 27988 4032
rect 28040 4020 28046 4072
rect 28276 4004 28304 4100
rect 29196 4069 29224 4100
rect 29564 4069 29592 4100
rect 29656 4100 30144 4128
rect 30208 4100 30564 4128
rect 29656 4072 29684 4100
rect 28445 4063 28503 4069
rect 28445 4029 28457 4063
rect 28491 4029 28503 4063
rect 28445 4023 28503 4029
rect 29181 4063 29239 4069
rect 29181 4029 29193 4063
rect 29227 4029 29239 4063
rect 29181 4023 29239 4029
rect 29273 4063 29331 4069
rect 29273 4029 29285 4063
rect 29319 4029 29331 4063
rect 29273 4023 29331 4029
rect 29549 4063 29607 4069
rect 29549 4029 29561 4063
rect 29595 4029 29607 4063
rect 29549 4023 29607 4029
rect 24578 3952 24584 4004
rect 24636 3992 24642 4004
rect 24673 3995 24731 4001
rect 24673 3992 24685 3995
rect 24636 3964 24685 3992
rect 24636 3952 24642 3964
rect 24673 3961 24685 3964
rect 24719 3961 24731 3995
rect 24673 3955 24731 3961
rect 25900 3995 25958 4001
rect 25900 3961 25912 3995
rect 25946 3992 25958 3995
rect 26326 3992 26332 4004
rect 25946 3964 26332 3992
rect 25946 3961 25958 3964
rect 25900 3955 25958 3961
rect 26326 3952 26332 3964
rect 26384 3952 26390 4004
rect 27246 3952 27252 4004
rect 27304 3992 27310 4004
rect 27718 3995 27776 4001
rect 27718 3992 27730 3995
rect 27304 3964 27730 3992
rect 27304 3952 27310 3964
rect 27718 3961 27730 3964
rect 27764 3992 27776 3995
rect 28258 3992 28264 4004
rect 27764 3964 28264 3992
rect 27764 3961 27776 3964
rect 27718 3955 27776 3961
rect 28258 3952 28264 3964
rect 28316 3952 28322 4004
rect 24486 3933 24492 3936
rect 24049 3896 24440 3924
rect 24473 3927 24492 3933
rect 24049 3893 24061 3896
rect 24003 3887 24061 3893
rect 24473 3893 24485 3927
rect 24473 3887 24492 3893
rect 24486 3884 24492 3887
rect 24544 3884 24550 3936
rect 26602 3884 26608 3936
rect 26660 3884 26666 3936
rect 27798 3884 27804 3936
rect 27856 3924 27862 3936
rect 28460 3924 28488 4023
rect 28537 3995 28595 4001
rect 28537 3961 28549 3995
rect 28583 3992 28595 3995
rect 29089 3995 29147 4001
rect 29089 3992 29101 3995
rect 28583 3964 29101 3992
rect 28583 3961 28595 3964
rect 28537 3955 28595 3961
rect 29089 3961 29101 3964
rect 29135 3992 29147 3995
rect 29288 3992 29316 4023
rect 29638 4020 29644 4072
rect 29696 4020 29702 4072
rect 30116 4069 30144 4100
rect 30558 4088 30564 4100
rect 30616 4128 30622 4140
rect 30616 4100 30696 4128
rect 30616 4088 30622 4100
rect 30668 4069 30696 4100
rect 29825 4063 29883 4069
rect 29825 4029 29837 4063
rect 29871 4029 29883 4063
rect 29825 4023 29883 4029
rect 30101 4063 30159 4069
rect 30101 4029 30113 4063
rect 30147 4060 30159 4063
rect 30377 4063 30435 4069
rect 30377 4060 30389 4063
rect 30147 4032 30389 4060
rect 30147 4029 30159 4032
rect 30101 4023 30159 4029
rect 30377 4029 30389 4032
rect 30423 4029 30435 4063
rect 30377 4023 30435 4029
rect 30653 4063 30711 4069
rect 30653 4029 30665 4063
rect 30699 4029 30711 4063
rect 30653 4023 30711 4029
rect 29840 3992 29868 4023
rect 29135 3964 29868 3992
rect 29135 3961 29147 3964
rect 29089 3955 29147 3961
rect 27856 3896 28488 3924
rect 27856 3884 27862 3896
rect 29638 3884 29644 3936
rect 29696 3884 29702 3936
rect 29914 3884 29920 3936
rect 29972 3884 29978 3936
rect 30466 3884 30472 3936
rect 30524 3884 30530 3936
rect 552 3834 31531 3856
rect 552 3782 8102 3834
rect 8154 3782 8166 3834
rect 8218 3782 8230 3834
rect 8282 3782 8294 3834
rect 8346 3782 8358 3834
rect 8410 3782 15807 3834
rect 15859 3782 15871 3834
rect 15923 3782 15935 3834
rect 15987 3782 15999 3834
rect 16051 3782 16063 3834
rect 16115 3782 23512 3834
rect 23564 3782 23576 3834
rect 23628 3782 23640 3834
rect 23692 3782 23704 3834
rect 23756 3782 23768 3834
rect 23820 3782 31217 3834
rect 31269 3782 31281 3834
rect 31333 3782 31345 3834
rect 31397 3782 31409 3834
rect 31461 3782 31473 3834
rect 31525 3782 31531 3834
rect 552 3760 31531 3782
rect 934 3680 940 3732
rect 992 3680 998 3732
rect 1854 3680 1860 3732
rect 1912 3720 1918 3732
rect 1949 3723 2007 3729
rect 1949 3720 1961 3723
rect 1912 3692 1961 3720
rect 1912 3680 1918 3692
rect 1949 3689 1961 3692
rect 1995 3720 2007 3723
rect 2498 3720 2504 3732
rect 1995 3692 2504 3720
rect 1995 3689 2007 3692
rect 1949 3683 2007 3689
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 3510 3720 3516 3732
rect 2746 3692 3516 3720
rect 952 3584 980 3680
rect 2225 3655 2283 3661
rect 2225 3652 2237 3655
rect 1596 3624 2237 3652
rect 1596 3593 1624 3624
rect 2225 3621 2237 3624
rect 2271 3652 2283 3655
rect 2271 3624 2452 3652
rect 2271 3621 2283 3624
rect 2225 3615 2283 3621
rect 1305 3587 1363 3593
rect 1305 3584 1317 3587
rect 952 3556 1317 3584
rect 1305 3553 1317 3556
rect 1351 3553 1363 3587
rect 1305 3547 1363 3553
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3584 1455 3587
rect 1581 3587 1639 3593
rect 1581 3584 1593 3587
rect 1443 3556 1593 3584
rect 1443 3553 1455 3556
rect 1397 3547 1455 3553
rect 1581 3553 1593 3556
rect 1627 3553 1639 3587
rect 1581 3547 1639 3553
rect 1320 3516 1348 3547
rect 2038 3544 2044 3596
rect 2096 3544 2102 3596
rect 2314 3544 2320 3596
rect 2372 3544 2378 3596
rect 2424 3593 2452 3624
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3553 2467 3587
rect 2746 3584 2774 3692
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 4157 3723 4215 3729
rect 4157 3689 4169 3723
rect 4203 3720 4215 3723
rect 12739 3723 12797 3729
rect 4203 3692 8524 3720
rect 4203 3689 4215 3692
rect 4157 3683 4215 3689
rect 7282 3652 7288 3664
rect 6564 3624 7288 3652
rect 3050 3593 3056 3596
rect 2746 3556 2820 3584
rect 2409 3547 2467 3553
rect 2130 3516 2136 3528
rect 1320 3488 2136 3516
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 2792 3525 2820 3556
rect 3044 3547 3056 3593
rect 3050 3544 3056 3547
rect 3108 3544 3114 3596
rect 6564 3593 6592 3624
rect 7282 3612 7288 3624
rect 7340 3652 7346 3664
rect 7340 3624 7972 3652
rect 7340 3612 7346 3624
rect 6822 3593 6828 3596
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3553 6607 3587
rect 6549 3547 6607 3553
rect 6816 3547 6828 3593
rect 6822 3544 6828 3547
rect 6880 3544 6886 3596
rect 7944 3528 7972 3624
rect 8110 3544 8116 3596
rect 8168 3584 8174 3596
rect 8277 3587 8335 3593
rect 8277 3584 8289 3587
rect 8168 3556 8289 3584
rect 8168 3544 8174 3556
rect 8277 3553 8289 3556
rect 8323 3553 8335 3587
rect 8496 3584 8524 3692
rect 12739 3689 12751 3723
rect 12785 3720 12797 3723
rect 13817 3723 13875 3729
rect 12785 3692 13242 3720
rect 12785 3689 12797 3692
rect 12739 3683 12797 3689
rect 11606 3612 11612 3664
rect 11664 3652 11670 3664
rect 12529 3655 12587 3661
rect 12529 3652 12541 3655
rect 11664 3624 12541 3652
rect 11664 3612 11670 3624
rect 12529 3621 12541 3624
rect 12575 3621 12587 3655
rect 13015 3655 13073 3661
rect 13015 3652 13027 3655
rect 12529 3615 12587 3621
rect 12728 3624 13027 3652
rect 12728 3596 12756 3624
rect 13015 3621 13027 3624
rect 13061 3621 13073 3655
rect 13214 3652 13242 3692
rect 13817 3689 13829 3723
rect 13863 3720 13875 3723
rect 13906 3720 13912 3732
rect 13863 3692 13912 3720
rect 13863 3689 13875 3692
rect 13817 3683 13875 3689
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 14826 3729 14832 3732
rect 14813 3723 14832 3729
rect 14813 3720 14825 3723
rect 14108 3692 14825 3720
rect 13214 3627 13248 3652
rect 13214 3624 13277 3627
rect 13015 3615 13073 3621
rect 13219 3621 13277 3624
rect 12618 3584 12624 3596
rect 8496 3556 12624 3584
rect 8277 3547 8335 3553
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 12710 3544 12716 3596
rect 12768 3544 12774 3596
rect 13219 3587 13231 3621
rect 13265 3596 13277 3621
rect 13446 3612 13452 3664
rect 13504 3612 13510 3664
rect 13665 3655 13723 3661
rect 13665 3652 13677 3655
rect 13556 3624 13677 3652
rect 13265 3587 13268 3596
rect 13219 3581 13268 3587
rect 13220 3556 13268 3581
rect 13262 3544 13268 3556
rect 13320 3584 13326 3596
rect 13556 3584 13584 3624
rect 13665 3621 13677 3624
rect 13711 3652 13723 3655
rect 14108 3652 14136 3692
rect 14813 3689 14825 3692
rect 14813 3683 14832 3689
rect 14826 3680 14832 3683
rect 14884 3680 14890 3732
rect 15102 3680 15108 3732
rect 15160 3680 15166 3732
rect 15273 3723 15331 3729
rect 15273 3689 15285 3723
rect 15319 3720 15331 3723
rect 16482 3720 16488 3732
rect 16540 3729 16546 3732
rect 16540 3723 16559 3729
rect 15319 3692 16488 3720
rect 15319 3689 15331 3692
rect 15273 3683 15331 3689
rect 13711 3624 14136 3652
rect 13711 3621 13723 3624
rect 13665 3615 13723 3621
rect 14182 3612 14188 3664
rect 14240 3612 14246 3664
rect 14401 3655 14459 3661
rect 14401 3621 14413 3655
rect 14447 3621 14459 3655
rect 14401 3615 14459 3621
rect 13320 3556 13584 3584
rect 14416 3584 14444 3615
rect 14642 3612 14648 3664
rect 14700 3652 14706 3664
rect 15013 3655 15071 3661
rect 15013 3652 15025 3655
rect 14700 3624 15025 3652
rect 14700 3612 14706 3624
rect 15013 3621 15025 3624
rect 15059 3621 15071 3655
rect 15013 3615 15071 3621
rect 15473 3655 15531 3661
rect 15473 3621 15485 3655
rect 15519 3621 15531 3655
rect 15473 3615 15531 3621
rect 14416 3556 14780 3584
rect 13320 3544 13326 3556
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3485 2835 3519
rect 2777 3479 2835 3485
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 7984 3488 8033 3516
rect 7984 3476 7990 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 13446 3516 13452 3528
rect 8021 3479 8079 3485
rect 12820 3488 13452 3516
rect 9401 3451 9459 3457
rect 9401 3417 9413 3451
rect 9447 3448 9459 3451
rect 12820 3448 12848 3488
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 14458 3476 14464 3528
rect 14516 3516 14522 3528
rect 14752 3516 14780 3556
rect 14918 3544 14924 3596
rect 14976 3584 14982 3596
rect 15488 3584 15516 3615
rect 14976 3556 15516 3584
rect 14976 3544 14982 3556
rect 15580 3516 15608 3692
rect 16482 3680 16488 3692
rect 16547 3720 16559 3723
rect 16547 3692 16620 3720
rect 16547 3689 16559 3692
rect 16540 3683 16559 3689
rect 16540 3680 16546 3683
rect 16206 3612 16212 3664
rect 16264 3612 16270 3664
rect 16298 3612 16304 3664
rect 16356 3612 16362 3664
rect 14516 3488 14688 3516
rect 14752 3488 15608 3516
rect 16224 3516 16252 3612
rect 16592 3584 16620 3692
rect 16666 3680 16672 3732
rect 16724 3680 16730 3732
rect 17218 3680 17224 3732
rect 17276 3729 17282 3732
rect 17276 3723 17295 3729
rect 17283 3720 17295 3723
rect 17405 3723 17463 3729
rect 17283 3692 17356 3720
rect 17283 3689 17295 3692
rect 17276 3683 17295 3689
rect 17276 3680 17282 3683
rect 17037 3655 17095 3661
rect 17037 3621 17049 3655
rect 17083 3652 17095 3655
rect 17126 3652 17132 3664
rect 17083 3624 17132 3652
rect 17083 3621 17095 3624
rect 17037 3615 17095 3621
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 17328 3652 17356 3692
rect 17405 3689 17417 3723
rect 17451 3720 17463 3723
rect 17494 3720 17500 3732
rect 17451 3692 17500 3720
rect 17451 3689 17463 3692
rect 17405 3683 17463 3689
rect 17494 3680 17500 3692
rect 17552 3680 17558 3732
rect 18874 3680 18880 3732
rect 18932 3680 18938 3732
rect 19334 3680 19340 3732
rect 19392 3680 19398 3732
rect 19610 3680 19616 3732
rect 19668 3720 19674 3732
rect 20257 3723 20315 3729
rect 19668 3692 20208 3720
rect 19668 3680 19674 3692
rect 19058 3661 19064 3664
rect 19029 3655 19064 3661
rect 19029 3652 19041 3655
rect 17328 3624 19041 3652
rect 19029 3621 19041 3624
rect 19029 3615 19064 3621
rect 19058 3612 19064 3615
rect 19116 3612 19122 3664
rect 19150 3612 19156 3664
rect 19208 3652 19214 3664
rect 19245 3655 19303 3661
rect 19245 3652 19257 3655
rect 19208 3624 19257 3652
rect 19208 3612 19214 3624
rect 19245 3621 19257 3624
rect 19291 3621 19303 3655
rect 19500 3655 19558 3661
rect 19500 3652 19512 3655
rect 19245 3615 19303 3621
rect 19444 3624 19512 3652
rect 19444 3584 19472 3624
rect 19500 3621 19512 3624
rect 19546 3621 19558 3655
rect 19500 3615 19558 3621
rect 19705 3655 19763 3661
rect 19705 3621 19717 3655
rect 19751 3621 19763 3655
rect 19705 3615 19763 3621
rect 19889 3655 19947 3661
rect 19889 3621 19901 3655
rect 19935 3652 19947 3655
rect 19978 3652 19984 3664
rect 19935 3624 19984 3652
rect 19935 3621 19947 3624
rect 19889 3615 19947 3621
rect 19720 3584 19748 3615
rect 19978 3612 19984 3624
rect 20036 3612 20042 3664
rect 20089 3655 20147 3661
rect 20089 3652 20101 3655
rect 20088 3621 20101 3652
rect 20135 3621 20147 3655
rect 20180 3652 20208 3692
rect 20257 3689 20269 3723
rect 20303 3720 20315 3723
rect 20622 3720 20628 3732
rect 20303 3692 20628 3720
rect 20303 3689 20315 3692
rect 20257 3683 20315 3689
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 21266 3680 21272 3732
rect 21324 3680 21330 3732
rect 21910 3729 21916 3732
rect 21729 3723 21787 3729
rect 21729 3720 21741 3723
rect 21376 3692 21741 3720
rect 21376 3652 21404 3692
rect 21729 3689 21741 3692
rect 21775 3689 21787 3723
rect 21729 3683 21787 3689
rect 21897 3723 21916 3729
rect 21897 3689 21909 3723
rect 21968 3720 21974 3732
rect 22646 3720 22652 3732
rect 21968 3692 22652 3720
rect 21897 3683 21916 3689
rect 21910 3680 21916 3683
rect 21968 3680 21974 3692
rect 22646 3680 22652 3692
rect 22704 3680 22710 3732
rect 23198 3680 23204 3732
rect 23256 3720 23262 3732
rect 23493 3723 23551 3729
rect 23493 3720 23505 3723
rect 23256 3692 23505 3720
rect 23256 3680 23262 3692
rect 23493 3689 23505 3692
rect 23539 3720 23551 3723
rect 23661 3723 23719 3729
rect 23539 3692 23612 3720
rect 23539 3689 23551 3692
rect 23493 3683 23551 3689
rect 20180 3624 21404 3652
rect 21437 3655 21495 3661
rect 20088 3615 20147 3621
rect 21437 3621 21449 3655
rect 21483 3652 21495 3655
rect 21483 3621 21496 3652
rect 21437 3615 21496 3621
rect 16592 3556 19472 3584
rect 19058 3516 19064 3528
rect 16224 3488 19064 3516
rect 14516 3476 14522 3488
rect 9447 3420 12848 3448
rect 12897 3451 12955 3457
rect 9447 3417 9459 3420
rect 9401 3411 9459 3417
rect 12897 3417 12909 3451
rect 12943 3448 12955 3451
rect 13357 3451 13415 3457
rect 12943 3420 13308 3448
rect 12943 3417 12955 3420
rect 12897 3411 12955 3417
rect 1673 3383 1731 3389
rect 1673 3349 1685 3383
rect 1719 3380 1731 3383
rect 3050 3380 3056 3392
rect 1719 3352 3056 3380
rect 1719 3349 1731 3352
rect 1673 3343 1731 3349
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 7929 3383 7987 3389
rect 7929 3349 7941 3383
rect 7975 3380 7987 3383
rect 11974 3380 11980 3392
rect 7975 3352 11980 3380
rect 7975 3349 7987 3352
rect 7929 3343 7987 3349
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12713 3383 12771 3389
rect 12713 3349 12725 3383
rect 12759 3380 12771 3383
rect 12802 3380 12808 3392
rect 12759 3352 12808 3380
rect 12759 3349 12771 3352
rect 12713 3343 12771 3349
rect 12802 3340 12808 3352
rect 12860 3380 12866 3392
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 12860 3352 13185 3380
rect 12860 3340 12866 3352
rect 13173 3349 13185 3352
rect 13219 3349 13231 3383
rect 13280 3380 13308 3420
rect 13357 3417 13369 3451
rect 13403 3448 13415 3451
rect 13722 3448 13728 3460
rect 13403 3420 13728 3448
rect 13403 3417 13415 3420
rect 13357 3411 13415 3417
rect 13722 3408 13728 3420
rect 13780 3408 13786 3460
rect 13814 3408 13820 3460
rect 13872 3448 13878 3460
rect 13872 3420 14504 3448
rect 13872 3408 13878 3420
rect 13538 3380 13544 3392
rect 13280 3352 13544 3380
rect 13173 3343 13231 3349
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 14369 3383 14427 3389
rect 14369 3380 14381 3383
rect 13688 3352 14381 3380
rect 13688 3340 13694 3352
rect 14369 3349 14381 3352
rect 14415 3349 14427 3383
rect 14476 3380 14504 3420
rect 14550 3408 14556 3460
rect 14608 3408 14614 3460
rect 14660 3457 14688 3488
rect 19058 3476 19064 3488
rect 19116 3476 19122 3528
rect 14645 3451 14703 3457
rect 14645 3417 14657 3451
rect 14691 3417 14703 3451
rect 18414 3448 18420 3460
rect 14645 3411 14703 3417
rect 14752 3420 18420 3448
rect 14752 3380 14780 3420
rect 18414 3408 18420 3420
rect 18472 3408 18478 3460
rect 19444 3448 19472 3556
rect 19536 3556 19748 3584
rect 20088 3584 20116 3615
rect 21468 3584 21496 3615
rect 21542 3612 21548 3664
rect 21600 3652 21606 3664
rect 21637 3655 21695 3661
rect 21637 3652 21649 3655
rect 21600 3624 21649 3652
rect 21600 3612 21606 3624
rect 21637 3621 21649 3624
rect 21683 3621 21695 3655
rect 21637 3615 21695 3621
rect 21928 3584 21956 3680
rect 22002 3612 22008 3664
rect 22060 3652 22066 3664
rect 22097 3655 22155 3661
rect 22097 3652 22109 3655
rect 22060 3624 22109 3652
rect 22060 3612 22066 3624
rect 22097 3621 22109 3624
rect 22143 3621 22155 3655
rect 22097 3615 22155 3621
rect 20088 3556 21956 3584
rect 19536 3528 19564 3556
rect 19518 3476 19524 3528
rect 19576 3476 19582 3528
rect 20088 3448 20116 3556
rect 19444 3420 20116 3448
rect 14476 3352 14780 3380
rect 14829 3383 14887 3389
rect 14369 3343 14427 3349
rect 14829 3349 14841 3383
rect 14875 3380 14887 3383
rect 15194 3380 15200 3392
rect 14875 3352 15200 3380
rect 14875 3349 14887 3352
rect 14829 3343 14887 3349
rect 15194 3340 15200 3352
rect 15252 3380 15258 3392
rect 15289 3383 15347 3389
rect 15289 3380 15301 3383
rect 15252 3352 15301 3380
rect 15252 3340 15258 3352
rect 15289 3349 15301 3352
rect 15335 3380 15347 3383
rect 16485 3383 16543 3389
rect 16485 3380 16497 3383
rect 15335 3352 16497 3380
rect 15335 3349 15347 3352
rect 15289 3343 15347 3349
rect 16485 3349 16497 3352
rect 16531 3380 16543 3383
rect 16758 3380 16764 3392
rect 16531 3352 16764 3380
rect 16531 3349 16543 3352
rect 16485 3343 16543 3349
rect 16758 3340 16764 3352
rect 16816 3380 16822 3392
rect 17221 3383 17279 3389
rect 17221 3380 17233 3383
rect 16816 3352 17233 3380
rect 16816 3340 16822 3352
rect 17221 3349 17233 3352
rect 17267 3380 17279 3383
rect 18046 3380 18052 3392
rect 17267 3352 18052 3380
rect 17267 3349 17279 3352
rect 17221 3343 17279 3349
rect 18046 3340 18052 3352
rect 18104 3380 18110 3392
rect 18966 3380 18972 3392
rect 18104 3352 18972 3380
rect 18104 3340 18110 3352
rect 18966 3340 18972 3352
rect 19024 3340 19030 3392
rect 19058 3340 19064 3392
rect 19116 3340 19122 3392
rect 19242 3340 19248 3392
rect 19300 3380 19306 3392
rect 19521 3383 19579 3389
rect 19521 3380 19533 3383
rect 19300 3352 19533 3380
rect 19300 3340 19306 3352
rect 19521 3349 19533 3352
rect 19567 3380 19579 3383
rect 20073 3383 20131 3389
rect 20073 3380 20085 3383
rect 19567 3352 20085 3380
rect 19567 3349 19579 3352
rect 19521 3343 19579 3349
rect 20073 3349 20085 3352
rect 20119 3349 20131 3383
rect 20073 3343 20131 3349
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 21453 3383 21511 3389
rect 21453 3380 21465 3383
rect 20772 3352 21465 3380
rect 20772 3340 20778 3352
rect 21453 3349 21465 3352
rect 21499 3380 21511 3383
rect 21726 3380 21732 3392
rect 21499 3352 21732 3380
rect 21499 3349 21511 3352
rect 21453 3343 21511 3349
rect 21726 3340 21732 3352
rect 21784 3380 21790 3392
rect 21913 3383 21971 3389
rect 21913 3380 21925 3383
rect 21784 3352 21925 3380
rect 21784 3340 21790 3352
rect 21913 3349 21925 3352
rect 21959 3349 21971 3383
rect 22664 3380 22692 3680
rect 23293 3655 23351 3661
rect 23293 3621 23305 3655
rect 23339 3621 23351 3655
rect 23584 3652 23612 3692
rect 23661 3689 23673 3723
rect 23707 3720 23719 3723
rect 24394 3720 24400 3732
rect 23707 3692 24400 3720
rect 23707 3689 23719 3692
rect 23661 3683 23719 3689
rect 24394 3680 24400 3692
rect 24452 3680 24458 3732
rect 24578 3680 24584 3732
rect 24636 3680 24642 3732
rect 27246 3680 27252 3732
rect 27304 3680 27310 3732
rect 27525 3723 27583 3729
rect 27525 3689 27537 3723
rect 27571 3720 27583 3723
rect 27706 3720 27712 3732
rect 27571 3692 27712 3720
rect 27571 3689 27583 3692
rect 27525 3683 27583 3689
rect 27706 3680 27712 3692
rect 27764 3720 27770 3732
rect 27801 3723 27859 3729
rect 27801 3720 27813 3723
rect 27764 3692 27813 3720
rect 27764 3680 27770 3692
rect 27801 3689 27813 3692
rect 27847 3689 27859 3723
rect 27801 3683 27859 3689
rect 24486 3652 24492 3664
rect 23584 3624 24492 3652
rect 23293 3615 23351 3621
rect 23308 3584 23336 3615
rect 24486 3612 24492 3624
rect 24544 3612 24550 3664
rect 25590 3612 25596 3664
rect 25648 3652 25654 3664
rect 25694 3655 25752 3661
rect 25694 3652 25706 3655
rect 25648 3624 25706 3652
rect 25648 3612 25654 3624
rect 25694 3621 25706 3624
rect 25740 3652 25752 3655
rect 27816 3652 27844 3683
rect 28258 3680 28264 3732
rect 28316 3720 28322 3732
rect 28721 3723 28779 3729
rect 28721 3720 28733 3723
rect 28316 3692 28733 3720
rect 28316 3680 28322 3692
rect 28721 3689 28733 3692
rect 28767 3689 28779 3723
rect 28721 3683 28779 3689
rect 28902 3680 28908 3732
rect 28960 3720 28966 3732
rect 28997 3723 29055 3729
rect 28997 3720 29009 3723
rect 28960 3692 29009 3720
rect 28960 3680 28966 3692
rect 28997 3689 29009 3692
rect 29043 3689 29055 3723
rect 28997 3683 29055 3689
rect 29365 3723 29423 3729
rect 29365 3689 29377 3723
rect 29411 3720 29423 3723
rect 29638 3720 29644 3732
rect 29411 3692 29644 3720
rect 29411 3689 29423 3692
rect 29365 3683 29423 3689
rect 29012 3652 29040 3683
rect 29638 3680 29644 3692
rect 29696 3680 29702 3732
rect 29794 3655 29852 3661
rect 29794 3652 29806 3655
rect 25740 3624 26832 3652
rect 25740 3621 25752 3624
rect 25694 3615 25752 3621
rect 25406 3584 25412 3596
rect 23308 3556 25412 3584
rect 25406 3544 25412 3556
rect 25464 3544 25470 3596
rect 26804 3593 26832 3624
rect 27172 3624 27752 3652
rect 27816 3624 28120 3652
rect 29012 3624 29806 3652
rect 27172 3596 27200 3624
rect 26789 3587 26847 3593
rect 26789 3553 26801 3587
rect 26835 3553 26847 3587
rect 26789 3547 26847 3553
rect 26881 3587 26939 3593
rect 26881 3553 26893 3587
rect 26927 3584 26939 3587
rect 27154 3584 27160 3596
rect 26927 3556 27160 3584
rect 26927 3553 26939 3556
rect 26881 3547 26939 3553
rect 27154 3544 27160 3556
rect 27212 3544 27218 3596
rect 27246 3544 27252 3596
rect 27304 3584 27310 3596
rect 27724 3593 27752 3624
rect 27433 3587 27491 3593
rect 27433 3584 27445 3587
rect 27304 3556 27445 3584
rect 27304 3544 27310 3556
rect 27433 3553 27445 3556
rect 27479 3553 27491 3587
rect 27433 3547 27491 3553
rect 27709 3587 27767 3593
rect 27709 3553 27721 3587
rect 27755 3553 27767 3587
rect 27709 3547 27767 3553
rect 27982 3544 27988 3596
rect 28040 3544 28046 3596
rect 28092 3584 28120 3624
rect 28353 3587 28411 3593
rect 28353 3584 28365 3587
rect 28092 3556 28365 3584
rect 28353 3553 28365 3556
rect 28399 3553 28411 3587
rect 28353 3547 28411 3553
rect 28445 3587 28503 3593
rect 28445 3553 28457 3587
rect 28491 3584 28503 3587
rect 28813 3587 28871 3593
rect 28813 3584 28825 3587
rect 28491 3556 28825 3584
rect 28491 3553 28503 3556
rect 28445 3547 28503 3553
rect 28813 3553 28825 3556
rect 28859 3584 28871 3587
rect 29086 3584 29092 3596
rect 28859 3556 29092 3584
rect 28859 3553 28871 3556
rect 28813 3547 28871 3553
rect 29086 3544 29092 3556
rect 29144 3544 29150 3596
rect 29288 3593 29316 3624
rect 29794 3621 29806 3624
rect 29840 3652 29852 3655
rect 29914 3652 29920 3664
rect 29840 3624 29920 3652
rect 29840 3621 29852 3624
rect 29794 3615 29852 3621
rect 29914 3612 29920 3624
rect 29972 3612 29978 3664
rect 29273 3587 29331 3593
rect 29273 3553 29285 3587
rect 29319 3553 29331 3587
rect 29273 3547 29331 3553
rect 25961 3519 26019 3525
rect 25961 3485 25973 3519
rect 26007 3516 26019 3519
rect 26050 3516 26056 3528
rect 26007 3488 26056 3516
rect 26007 3485 26019 3488
rect 25961 3479 26019 3485
rect 23477 3383 23535 3389
rect 23477 3380 23489 3383
rect 22664 3352 23489 3380
rect 21913 3343 21971 3349
rect 23477 3349 23489 3352
rect 23523 3349 23535 3383
rect 23477 3343 23535 3349
rect 25222 3340 25228 3392
rect 25280 3380 25286 3392
rect 25976 3380 26004 3479
rect 26050 3476 26056 3488
rect 26108 3476 26114 3528
rect 28000 3516 28028 3544
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 28000 3488 29561 3516
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 25280 3352 26004 3380
rect 25280 3340 25286 3352
rect 30926 3340 30932 3392
rect 30984 3340 30990 3392
rect 552 3290 31372 3312
rect 552 3238 4250 3290
rect 4302 3238 4314 3290
rect 4366 3238 4378 3290
rect 4430 3238 4442 3290
rect 4494 3238 4506 3290
rect 4558 3238 11955 3290
rect 12007 3238 12019 3290
rect 12071 3238 12083 3290
rect 12135 3238 12147 3290
rect 12199 3238 12211 3290
rect 12263 3238 19660 3290
rect 19712 3238 19724 3290
rect 19776 3238 19788 3290
rect 19840 3238 19852 3290
rect 19904 3238 19916 3290
rect 19968 3238 27365 3290
rect 27417 3238 27429 3290
rect 27481 3238 27493 3290
rect 27545 3238 27557 3290
rect 27609 3238 27621 3290
rect 27673 3238 31372 3290
rect 552 3216 31372 3238
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3050 3176 3056 3188
rect 3007 3148 3056 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 8110 3176 8116 3188
rect 7248 3148 8116 3176
rect 7248 3136 7254 3148
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8205 3179 8263 3185
rect 8205 3145 8217 3179
rect 8251 3176 8263 3179
rect 11514 3176 11520 3188
rect 8251 3148 11520 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 12621 3179 12679 3185
rect 12621 3145 12633 3179
rect 12667 3176 12679 3179
rect 12710 3176 12716 3188
rect 12667 3148 12716 3176
rect 12667 3145 12679 3148
rect 12621 3139 12679 3145
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 12989 3179 13047 3185
rect 12989 3176 13001 3179
rect 12860 3148 13001 3176
rect 12860 3136 12866 3148
rect 12989 3145 13001 3148
rect 13035 3145 13047 3179
rect 12989 3139 13047 3145
rect 10965 3111 11023 3117
rect 10965 3077 10977 3111
rect 11011 3108 11023 3111
rect 11238 3108 11244 3120
rect 11011 3080 11244 3108
rect 11011 3077 11023 3080
rect 10965 3071 11023 3077
rect 11238 3068 11244 3080
rect 11296 3068 11302 3120
rect 13004 3108 13032 3139
rect 13170 3136 13176 3188
rect 13228 3136 13234 3188
rect 13354 3136 13360 3188
rect 13412 3136 13418 3188
rect 14458 3136 14464 3188
rect 14516 3136 14522 3188
rect 14918 3136 14924 3188
rect 14976 3136 14982 3188
rect 15028 3148 16896 3176
rect 13372 3108 13400 3136
rect 13004 3080 13400 3108
rect 14476 3108 14504 3136
rect 15028 3108 15056 3148
rect 14476 3080 15056 3108
rect 16868 3108 16896 3148
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17129 3179 17187 3185
rect 17129 3176 17141 3179
rect 17000 3148 17141 3176
rect 17000 3136 17006 3148
rect 17129 3145 17141 3148
rect 17175 3145 17187 3179
rect 17129 3139 17187 3145
rect 18693 3179 18751 3185
rect 18693 3145 18705 3179
rect 18739 3176 18751 3179
rect 19058 3176 19064 3188
rect 18739 3148 19064 3176
rect 18739 3145 18751 3148
rect 18693 3139 18751 3145
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 20806 3176 20812 3188
rect 19168 3148 20812 3176
rect 19168 3108 19196 3148
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 21450 3136 21456 3188
rect 21508 3136 21514 3188
rect 21542 3136 21548 3188
rect 21600 3136 21606 3188
rect 21928 3148 23244 3176
rect 16868 3080 19196 3108
rect 21468 3108 21496 3136
rect 21928 3108 21956 3148
rect 21468 3080 21956 3108
rect 23216 3108 23244 3148
rect 23290 3136 23296 3188
rect 23348 3136 23354 3188
rect 23382 3136 23388 3188
rect 23440 3176 23446 3188
rect 23845 3179 23903 3185
rect 23845 3176 23857 3179
rect 23440 3148 23857 3176
rect 23440 3136 23446 3148
rect 23845 3145 23857 3148
rect 23891 3145 23903 3179
rect 23845 3139 23903 3145
rect 23952 3148 28856 3176
rect 23952 3108 23980 3148
rect 23216 3080 23980 3108
rect 25406 3068 25412 3120
rect 25464 3068 25470 3120
rect 26605 3111 26663 3117
rect 26605 3077 26617 3111
rect 26651 3108 26663 3111
rect 27157 3111 27215 3117
rect 27157 3108 27169 3111
rect 26651 3080 27169 3108
rect 26651 3077 26663 3080
rect 26605 3071 26663 3077
rect 27157 3077 27169 3080
rect 27203 3108 27215 3111
rect 27246 3108 27252 3120
rect 27203 3080 27252 3108
rect 27203 3077 27215 3080
rect 27157 3071 27215 3077
rect 27246 3068 27252 3080
rect 27304 3068 27310 3120
rect 27433 3111 27491 3117
rect 27433 3077 27445 3111
rect 27479 3077 27491 3111
rect 28828 3108 28856 3148
rect 29086 3136 29092 3188
rect 29144 3136 29150 3188
rect 29917 3179 29975 3185
rect 29917 3145 29929 3179
rect 29963 3176 29975 3179
rect 30466 3176 30472 3188
rect 29963 3148 30472 3176
rect 29963 3145 29975 3148
rect 29917 3139 29975 3145
rect 30466 3136 30472 3148
rect 30524 3136 30530 3188
rect 30926 3136 30932 3188
rect 30984 3136 30990 3188
rect 30944 3108 30972 3136
rect 28828 3080 30972 3108
rect 27433 3071 27491 3077
rect 7926 3000 7932 3052
rect 7984 3000 7990 3052
rect 25424 3040 25452 3068
rect 27448 3040 27476 3071
rect 25424 3012 27476 3040
rect 1854 2932 1860 2984
rect 1912 2974 1918 2984
rect 1912 2946 1955 2974
rect 1912 2932 1918 2946
rect 2130 2932 2136 2984
rect 2188 2932 2194 2984
rect 2317 2975 2375 2981
rect 2317 2941 2329 2975
rect 2363 2941 2375 2975
rect 2317 2935 2375 2941
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2904 1823 2907
rect 2041 2907 2099 2913
rect 2041 2904 2053 2907
rect 1811 2876 2053 2904
rect 1811 2873 1823 2876
rect 1765 2867 1823 2873
rect 2041 2873 2053 2876
rect 2087 2904 2099 2907
rect 2332 2904 2360 2935
rect 2498 2932 2504 2984
rect 2556 2972 2562 2984
rect 2777 2975 2835 2981
rect 2777 2972 2789 2975
rect 2556 2944 2789 2972
rect 2556 2932 2562 2944
rect 2777 2941 2789 2944
rect 2823 2941 2835 2975
rect 2777 2935 2835 2941
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2941 2927 2975
rect 2869 2935 2927 2941
rect 3881 2975 3939 2981
rect 3881 2941 3893 2975
rect 3927 2972 3939 2975
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 3927 2944 5365 2972
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 5353 2941 5365 2944
rect 5399 2972 5411 2975
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 5399 2944 6837 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 6825 2941 6837 2944
rect 6871 2972 6883 2975
rect 7944 2972 7972 3000
rect 6871 2944 7972 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 2884 2904 2912 2935
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 9456 2944 9597 2972
rect 9456 2932 9462 2944
rect 9585 2941 9597 2944
rect 9631 2972 9643 2975
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 9631 2944 11253 2972
rect 9631 2941 9643 2944
rect 9585 2935 9643 2941
rect 11241 2941 11253 2944
rect 11287 2972 11299 2975
rect 12434 2972 12440 2984
rect 11287 2944 12440 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 12434 2932 12440 2944
rect 12492 2972 12498 2984
rect 13538 2972 13544 2984
rect 12492 2944 13544 2972
rect 12492 2932 12498 2944
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 15470 2932 15476 2984
rect 15528 2972 15534 2984
rect 15749 2975 15807 2981
rect 15749 2972 15761 2975
rect 15528 2944 15761 2972
rect 15528 2932 15534 2944
rect 15749 2941 15761 2944
rect 15795 2941 15807 2975
rect 15749 2935 15807 2941
rect 20070 2932 20076 2984
rect 20128 2972 20134 2984
rect 20165 2975 20223 2981
rect 20165 2972 20177 2975
rect 20128 2944 20177 2972
rect 20128 2932 20134 2944
rect 20165 2941 20177 2944
rect 20211 2972 20223 2975
rect 21174 2972 21180 2984
rect 20211 2944 21180 2972
rect 20211 2941 20223 2944
rect 20165 2935 20223 2941
rect 21174 2932 21180 2944
rect 21232 2972 21238 2984
rect 21910 2972 21916 2984
rect 21232 2944 21916 2972
rect 21232 2932 21238 2944
rect 21910 2932 21916 2944
rect 21968 2932 21974 2984
rect 25130 2932 25136 2984
rect 25188 2972 25194 2984
rect 25225 2975 25283 2981
rect 25225 2972 25237 2975
rect 25188 2944 25237 2972
rect 25188 2932 25194 2944
rect 25225 2941 25237 2944
rect 25271 2941 25283 2975
rect 25225 2935 25283 2941
rect 25317 2975 25375 2981
rect 25317 2941 25329 2975
rect 25363 2972 25375 2975
rect 25593 2975 25651 2981
rect 25363 2944 25397 2972
rect 25363 2941 25375 2944
rect 25317 2935 25375 2941
rect 25593 2941 25605 2975
rect 25639 2972 25651 2975
rect 25682 2972 25688 2984
rect 25639 2944 25688 2972
rect 25639 2941 25651 2944
rect 25593 2935 25651 2941
rect 2087 2876 2912 2904
rect 2087 2873 2099 2876
rect 2041 2867 2099 2873
rect 3970 2864 3976 2916
rect 4028 2904 4034 2916
rect 4126 2907 4184 2913
rect 4126 2904 4138 2907
rect 4028 2876 4138 2904
rect 4028 2864 4034 2876
rect 4126 2873 4138 2876
rect 4172 2873 4184 2907
rect 4126 2867 4184 2873
rect 5442 2864 5448 2916
rect 5500 2904 5506 2916
rect 7098 2913 7104 2916
rect 5598 2907 5656 2913
rect 5598 2904 5610 2907
rect 5500 2876 5610 2904
rect 5500 2864 5506 2876
rect 5598 2873 5610 2876
rect 5644 2873 5656 2907
rect 5598 2867 5656 2873
rect 7070 2907 7104 2913
rect 7070 2873 7082 2907
rect 7070 2867 7104 2873
rect 7098 2864 7104 2867
rect 7156 2864 7162 2916
rect 9858 2913 9864 2916
rect 9852 2867 9864 2913
rect 9858 2864 9864 2867
rect 9916 2864 9922 2916
rect 10410 2864 10416 2916
rect 10468 2864 10474 2916
rect 11054 2864 11060 2916
rect 11112 2904 11118 2916
rect 11486 2907 11544 2913
rect 11486 2904 11498 2907
rect 11112 2876 11498 2904
rect 11112 2864 11118 2876
rect 11486 2873 11498 2876
rect 11532 2873 11544 2907
rect 11486 2867 11544 2873
rect 12802 2864 12808 2916
rect 12860 2864 12866 2916
rect 12894 2864 12900 2916
rect 12952 2864 12958 2916
rect 13021 2907 13079 2913
rect 13021 2873 13033 2907
rect 13067 2904 13079 2907
rect 13262 2904 13268 2916
rect 13067 2876 13268 2904
rect 13067 2873 13079 2876
rect 13021 2867 13079 2873
rect 13262 2864 13268 2876
rect 13320 2864 13326 2916
rect 13808 2907 13866 2913
rect 13808 2873 13820 2907
rect 13854 2904 13866 2907
rect 14366 2904 14372 2916
rect 13854 2876 14372 2904
rect 13854 2873 13866 2876
rect 13808 2867 13866 2873
rect 14366 2864 14372 2876
rect 14424 2864 14430 2916
rect 16016 2907 16074 2913
rect 16016 2873 16028 2907
rect 16062 2904 16074 2907
rect 16206 2904 16212 2916
rect 16062 2876 16212 2904
rect 16062 2873 16074 2876
rect 16016 2867 16074 2873
rect 16206 2864 16212 2876
rect 16264 2864 16270 2916
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 19806 2907 19864 2913
rect 19806 2904 19818 2907
rect 19484 2876 19818 2904
rect 19484 2864 19490 2876
rect 19806 2873 19818 2876
rect 19852 2873 19864 2907
rect 19806 2867 19864 2873
rect 20254 2864 20260 2916
rect 20312 2904 20318 2916
rect 20410 2907 20468 2913
rect 20410 2904 20422 2907
rect 20312 2876 20422 2904
rect 20312 2864 20318 2876
rect 20410 2873 20422 2876
rect 20456 2873 20468 2907
rect 20410 2867 20468 2873
rect 22180 2907 22238 2913
rect 22180 2873 22192 2907
rect 22226 2904 22238 2907
rect 24026 2904 24032 2916
rect 22226 2876 24032 2904
rect 22226 2873 22238 2876
rect 22180 2867 22238 2873
rect 24026 2864 24032 2876
rect 24084 2864 24090 2916
rect 24946 2864 24952 2916
rect 25004 2913 25010 2916
rect 25004 2904 25016 2913
rect 25332 2904 25360 2935
rect 25682 2932 25688 2944
rect 25740 2932 25746 2984
rect 26053 2975 26111 2981
rect 26053 2941 26065 2975
rect 26099 2972 26111 2975
rect 26145 2975 26203 2981
rect 26145 2972 26157 2975
rect 26099 2944 26157 2972
rect 26099 2941 26111 2944
rect 26053 2935 26111 2941
rect 26145 2941 26157 2944
rect 26191 2941 26203 2975
rect 26145 2935 26203 2941
rect 25004 2876 25049 2904
rect 25332 2876 25728 2904
rect 25004 2867 25016 2876
rect 25004 2864 25010 2867
rect 2406 2796 2412 2848
rect 2464 2796 2470 2848
rect 2682 2796 2688 2848
rect 2740 2796 2746 2848
rect 5258 2796 5264 2848
rect 5316 2796 5322 2848
rect 6733 2839 6791 2845
rect 6733 2805 6745 2839
rect 6779 2836 6791 2839
rect 10428 2836 10456 2864
rect 6779 2808 10456 2836
rect 12912 2836 12940 2864
rect 25332 2848 25360 2876
rect 22554 2836 22560 2848
rect 12912 2808 22560 2836
rect 6779 2805 6791 2808
rect 6733 2799 6791 2805
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 25314 2796 25320 2848
rect 25372 2796 25378 2848
rect 25409 2839 25467 2845
rect 25409 2805 25421 2839
rect 25455 2836 25467 2839
rect 25590 2836 25596 2848
rect 25455 2808 25596 2836
rect 25455 2805 25467 2808
rect 25409 2799 25467 2805
rect 25590 2796 25596 2808
rect 25648 2796 25654 2848
rect 25700 2845 25728 2876
rect 26160 2848 26188 2935
rect 26326 2932 26332 2984
rect 26384 2972 26390 2984
rect 26513 2975 26571 2981
rect 26513 2972 26525 2975
rect 26384 2944 26525 2972
rect 26384 2932 26390 2944
rect 26513 2941 26525 2944
rect 26559 2972 26571 2975
rect 26789 2975 26847 2981
rect 26789 2972 26801 2975
rect 26559 2944 26801 2972
rect 26559 2941 26571 2944
rect 26513 2935 26571 2941
rect 26789 2941 26801 2944
rect 26835 2941 26847 2975
rect 26789 2935 26847 2941
rect 27065 2975 27123 2981
rect 27065 2941 27077 2975
rect 27111 2941 27123 2975
rect 27065 2935 27123 2941
rect 26237 2907 26295 2913
rect 26237 2873 26249 2907
rect 26283 2904 26295 2907
rect 26694 2904 26700 2916
rect 26283 2876 26700 2904
rect 26283 2873 26295 2876
rect 26237 2867 26295 2873
rect 26694 2864 26700 2876
rect 26752 2904 26758 2916
rect 26881 2907 26939 2913
rect 26881 2904 26893 2907
rect 26752 2876 26893 2904
rect 26752 2864 26758 2876
rect 26881 2873 26893 2876
rect 26927 2873 26939 2907
rect 26881 2867 26939 2873
rect 25685 2839 25743 2845
rect 25685 2805 25697 2839
rect 25731 2836 25743 2839
rect 25961 2839 26019 2845
rect 25961 2836 25973 2839
rect 25731 2808 25973 2836
rect 25731 2805 25743 2808
rect 25685 2799 25743 2805
rect 25961 2805 25973 2808
rect 26007 2805 26019 2839
rect 25961 2799 26019 2805
rect 26142 2796 26148 2848
rect 26200 2796 26206 2848
rect 26602 2796 26608 2848
rect 26660 2836 26666 2848
rect 27080 2836 27108 2935
rect 27982 2932 27988 2984
rect 28040 2972 28046 2984
rect 28813 2975 28871 2981
rect 28813 2972 28825 2975
rect 28040 2944 28825 2972
rect 28040 2932 28046 2944
rect 28813 2941 28825 2944
rect 28859 2941 28871 2975
rect 28813 2935 28871 2941
rect 28997 2975 29055 2981
rect 28997 2941 29009 2975
rect 29043 2941 29055 2975
rect 28997 2935 29055 2941
rect 27522 2864 27528 2916
rect 27580 2904 27586 2916
rect 28568 2907 28626 2913
rect 28568 2904 28580 2907
rect 27580 2876 28580 2904
rect 27580 2864 27586 2876
rect 28568 2873 28580 2876
rect 28614 2904 28626 2907
rect 29012 2904 29040 2935
rect 29822 2932 29828 2984
rect 29880 2932 29886 2984
rect 31021 2975 31079 2981
rect 31021 2941 31033 2975
rect 31067 2972 31079 2975
rect 31570 2972 31576 2984
rect 31067 2944 31576 2972
rect 31067 2941 31079 2944
rect 31021 2935 31079 2941
rect 31570 2932 31576 2944
rect 31628 2932 31634 2984
rect 28614 2876 29040 2904
rect 28614 2873 28626 2876
rect 28568 2867 28626 2873
rect 26660 2808 27108 2836
rect 26660 2796 26666 2808
rect 552 2746 31531 2768
rect 552 2694 8102 2746
rect 8154 2694 8166 2746
rect 8218 2694 8230 2746
rect 8282 2694 8294 2746
rect 8346 2694 8358 2746
rect 8410 2694 15807 2746
rect 15859 2694 15871 2746
rect 15923 2694 15935 2746
rect 15987 2694 15999 2746
rect 16051 2694 16063 2746
rect 16115 2694 23512 2746
rect 23564 2694 23576 2746
rect 23628 2694 23640 2746
rect 23692 2694 23704 2746
rect 23756 2694 23768 2746
rect 23820 2694 31217 2746
rect 31269 2694 31281 2746
rect 31333 2694 31345 2746
rect 31397 2694 31409 2746
rect 31461 2694 31473 2746
rect 31525 2694 31531 2746
rect 552 2672 31531 2694
rect 2406 2592 2412 2644
rect 2464 2632 2470 2644
rect 2464 2604 3096 2632
rect 2464 2592 2470 2604
rect 2682 2564 2688 2576
rect 2516 2536 2688 2564
rect 2516 2505 2544 2536
rect 2682 2524 2688 2536
rect 2740 2524 2746 2576
rect 3068 2564 3096 2604
rect 3970 2592 3976 2644
rect 4028 2592 4034 2644
rect 10781 2635 10839 2641
rect 10781 2601 10793 2635
rect 10827 2632 10839 2635
rect 11606 2632 11612 2644
rect 10827 2604 11612 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 11606 2592 11612 2604
rect 11664 2592 11670 2644
rect 12989 2635 13047 2641
rect 12989 2601 13001 2635
rect 13035 2632 13047 2635
rect 13078 2632 13084 2644
rect 13035 2604 13084 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 13078 2592 13084 2604
rect 13136 2592 13142 2644
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 14642 2632 14648 2644
rect 14507 2604 14648 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 14642 2592 14648 2604
rect 14700 2592 14706 2644
rect 15933 2635 15991 2641
rect 15933 2601 15945 2635
rect 15979 2632 15991 2635
rect 16298 2632 16304 2644
rect 15979 2604 16304 2632
rect 15979 2601 15991 2604
rect 15933 2595 15991 2601
rect 16298 2592 16304 2604
rect 16356 2592 16362 2644
rect 17954 2592 17960 2644
rect 18012 2592 18018 2644
rect 19518 2592 19524 2644
rect 19576 2592 19582 2644
rect 20254 2592 20260 2644
rect 20312 2592 20318 2644
rect 24026 2592 24032 2644
rect 24084 2632 24090 2644
rect 24084 2604 24854 2632
rect 24084 2592 24090 2604
rect 3988 2564 4016 2592
rect 3068 2536 4016 2564
rect 2501 2499 2559 2505
rect 2501 2465 2513 2499
rect 2547 2465 2559 2499
rect 2501 2459 2559 2465
rect 2593 2499 2651 2505
rect 2593 2465 2605 2499
rect 2639 2496 2651 2499
rect 2774 2496 2780 2508
rect 2639 2468 2780 2496
rect 2639 2465 2651 2468
rect 2593 2459 2651 2465
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 3068 2505 3096 2536
rect 3988 2505 4016 2536
rect 5350 2524 5356 2576
rect 5408 2524 5414 2576
rect 7006 2524 7012 2576
rect 7064 2524 7070 2576
rect 13630 2564 13636 2576
rect 11624 2536 13636 2564
rect 3053 2499 3111 2505
rect 3053 2465 3065 2499
rect 3099 2465 3111 2499
rect 3053 2459 3111 2465
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3421 2499 3479 2505
rect 3421 2496 3433 2499
rect 3191 2468 3433 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 3421 2465 3433 2468
rect 3467 2465 3479 2499
rect 3421 2459 3479 2465
rect 3697 2499 3755 2505
rect 3697 2465 3709 2499
rect 3743 2465 3755 2499
rect 3697 2459 3755 2465
rect 3973 2499 4031 2505
rect 3973 2465 3985 2499
rect 4019 2465 4031 2499
rect 4433 2499 4491 2505
rect 4433 2496 4445 2499
rect 3973 2459 4031 2465
rect 4080 2468 4445 2496
rect 3160 2428 3188 2459
rect 2976 2400 3188 2428
rect 2976 2369 3004 2400
rect 2685 2363 2743 2369
rect 2685 2329 2697 2363
rect 2731 2360 2743 2363
rect 2961 2363 3019 2369
rect 2961 2360 2973 2363
rect 2731 2332 2973 2360
rect 2731 2329 2743 2332
rect 2685 2323 2743 2329
rect 2961 2329 2973 2332
rect 3007 2329 3019 2363
rect 2961 2323 3019 2329
rect 3237 2363 3295 2369
rect 3237 2329 3249 2363
rect 3283 2360 3295 2363
rect 3326 2360 3332 2372
rect 3283 2332 3332 2360
rect 3283 2329 3295 2332
rect 3237 2323 3295 2329
rect 3326 2320 3332 2332
rect 3384 2360 3390 2372
rect 3712 2360 3740 2459
rect 4080 2437 4108 2468
rect 4433 2465 4445 2468
rect 4479 2496 4491 2499
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4479 2468 4629 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2496 5319 2499
rect 5368 2496 5396 2524
rect 5307 2468 5396 2496
rect 7024 2496 7052 2524
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 7024 2468 7205 2496
rect 5307 2465 5319 2468
rect 5261 2459 5319 2465
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7193 2459 7251 2465
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2428 3847 2431
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 3835 2400 4077 2428
rect 3835 2397 3847 2400
rect 3789 2391 3847 2397
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 5276 2360 5304 2459
rect 7926 2456 7932 2508
rect 7984 2456 7990 2508
rect 8202 2505 8208 2508
rect 8196 2459 8208 2505
rect 8202 2456 8208 2459
rect 8260 2456 8266 2508
rect 9398 2456 9404 2508
rect 9456 2456 9462 2508
rect 9674 2505 9680 2508
rect 9668 2459 9680 2505
rect 9674 2456 9680 2459
rect 9732 2456 9738 2508
rect 11514 2456 11520 2508
rect 11572 2496 11578 2508
rect 11624 2505 11652 2536
rect 11609 2499 11667 2505
rect 11609 2496 11621 2499
rect 11572 2468 11621 2496
rect 11572 2456 11578 2468
rect 11609 2465 11621 2468
rect 11655 2465 11667 2499
rect 11609 2459 11667 2465
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 13096 2505 13124 2536
rect 13630 2524 13636 2536
rect 13688 2564 13694 2576
rect 15470 2564 15476 2576
rect 13688 2536 15476 2564
rect 13688 2524 13694 2536
rect 11865 2499 11923 2505
rect 11865 2496 11877 2499
rect 11756 2468 11877 2496
rect 11756 2456 11762 2468
rect 11865 2465 11877 2468
rect 11911 2465 11923 2499
rect 11865 2459 11923 2465
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2465 13139 2499
rect 13081 2459 13139 2465
rect 13170 2456 13176 2508
rect 13228 2496 13234 2508
rect 13337 2499 13395 2505
rect 13337 2496 13349 2499
rect 13228 2468 13349 2496
rect 13228 2456 13234 2468
rect 13337 2465 13349 2468
rect 13383 2465 13395 2499
rect 13337 2459 13395 2465
rect 13722 2456 13728 2508
rect 13780 2496 13786 2508
rect 14568 2505 14596 2536
rect 15470 2524 15476 2536
rect 15528 2524 15534 2576
rect 16592 2536 18184 2564
rect 14553 2499 14611 2505
rect 13780 2468 14136 2496
rect 13780 2456 13786 2468
rect 14108 2428 14136 2468
rect 14553 2465 14565 2499
rect 14599 2465 14611 2499
rect 14809 2499 14867 2505
rect 14809 2496 14821 2499
rect 14553 2459 14611 2465
rect 14660 2468 14821 2496
rect 14660 2428 14688 2468
rect 14809 2465 14821 2468
rect 14855 2465 14867 2499
rect 14809 2459 14867 2465
rect 14108 2400 14688 2428
rect 16206 2388 16212 2440
rect 16264 2428 16270 2440
rect 16592 2437 16620 2536
rect 16850 2505 16856 2508
rect 16844 2496 16856 2505
rect 16811 2468 16856 2496
rect 16844 2459 16856 2468
rect 16850 2456 16856 2459
rect 16908 2456 16914 2508
rect 18156 2505 18184 2536
rect 21910 2524 21916 2576
rect 21968 2564 21974 2576
rect 24826 2564 24854 2604
rect 25590 2592 25596 2644
rect 25648 2632 25654 2644
rect 26602 2632 26608 2644
rect 25648 2604 26608 2632
rect 25648 2592 25654 2604
rect 26602 2592 26608 2604
rect 26660 2592 26666 2644
rect 26694 2592 26700 2644
rect 26752 2592 26758 2644
rect 27154 2592 27160 2644
rect 27212 2632 27218 2644
rect 27249 2635 27307 2641
rect 27249 2632 27261 2635
rect 27212 2604 27261 2632
rect 27212 2592 27218 2604
rect 27249 2601 27261 2604
rect 27295 2601 27307 2635
rect 27249 2595 27307 2601
rect 27522 2592 27528 2644
rect 27580 2592 27586 2644
rect 26142 2564 26148 2576
rect 21968 2536 23152 2564
rect 24826 2536 26148 2564
rect 21968 2524 21974 2536
rect 18141 2499 18199 2505
rect 18141 2465 18153 2499
rect 18187 2465 18199 2499
rect 18141 2459 18199 2465
rect 18230 2456 18236 2508
rect 18288 2496 18294 2508
rect 18397 2499 18455 2505
rect 18397 2496 18409 2499
rect 18288 2468 18409 2496
rect 18288 2456 18294 2468
rect 18397 2465 18409 2468
rect 18443 2465 18455 2499
rect 18397 2459 18455 2465
rect 20162 2456 20168 2508
rect 20220 2456 20226 2508
rect 22830 2456 22836 2508
rect 22888 2505 22894 2508
rect 23124 2505 23152 2536
rect 26142 2524 26148 2536
rect 26200 2524 26206 2576
rect 22888 2459 22900 2505
rect 23109 2499 23167 2505
rect 23109 2465 23121 2499
rect 23155 2465 23167 2499
rect 23109 2459 23167 2465
rect 22888 2456 22894 2459
rect 24118 2456 24124 2508
rect 24176 2496 24182 2508
rect 24213 2499 24271 2505
rect 24213 2496 24225 2499
rect 24176 2468 24225 2496
rect 24176 2456 24182 2468
rect 24213 2465 24225 2468
rect 24259 2465 24271 2499
rect 24213 2459 24271 2465
rect 25314 2456 25320 2508
rect 25372 2496 25378 2508
rect 25409 2499 25467 2505
rect 25409 2496 25421 2499
rect 25372 2468 25421 2496
rect 25372 2456 25378 2468
rect 25409 2465 25421 2468
rect 25455 2465 25467 2499
rect 25409 2459 25467 2465
rect 25501 2499 25559 2505
rect 25501 2465 25513 2499
rect 25547 2465 25559 2499
rect 25501 2459 25559 2465
rect 16577 2431 16635 2437
rect 16577 2428 16589 2431
rect 16264 2400 16589 2428
rect 16264 2388 16270 2400
rect 16577 2397 16589 2400
rect 16623 2397 16635 2431
rect 25516 2428 25544 2459
rect 25590 2456 25596 2508
rect 25648 2496 25654 2508
rect 26712 2505 26740 2592
rect 26881 2567 26939 2573
rect 26881 2533 26893 2567
rect 26927 2564 26939 2567
rect 27540 2564 27568 2592
rect 26927 2536 27568 2564
rect 26927 2533 26939 2536
rect 26881 2527 26939 2533
rect 25961 2499 26019 2505
rect 25961 2496 25973 2499
rect 25648 2468 25973 2496
rect 25648 2456 25654 2468
rect 25961 2465 25973 2468
rect 26007 2496 26019 2499
rect 26053 2499 26111 2505
rect 26053 2496 26065 2499
rect 26007 2468 26065 2496
rect 26007 2465 26019 2468
rect 25961 2459 26019 2465
rect 26053 2465 26065 2468
rect 26099 2465 26111 2499
rect 26053 2459 26111 2465
rect 26697 2499 26755 2505
rect 26697 2465 26709 2499
rect 26743 2496 26755 2499
rect 26789 2499 26847 2505
rect 26789 2496 26801 2499
rect 26743 2468 26801 2496
rect 26743 2465 26755 2468
rect 26697 2459 26755 2465
rect 26789 2465 26801 2468
rect 26835 2465 26847 2499
rect 26789 2459 26847 2465
rect 27246 2456 27252 2508
rect 27304 2456 27310 2508
rect 27356 2505 27384 2536
rect 27341 2499 27399 2505
rect 27341 2465 27353 2499
rect 27387 2465 27399 2499
rect 27341 2459 27399 2465
rect 27433 2499 27491 2505
rect 27433 2465 27445 2499
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 25682 2428 25688 2440
rect 16577 2391 16635 2397
rect 24964 2400 25688 2428
rect 3384 2332 5304 2360
rect 10704 2332 10916 2360
rect 3384 2320 3390 2332
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 4341 2295 4399 2301
rect 4341 2292 4353 2295
rect 3559 2264 4353 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 4341 2261 4353 2264
rect 4387 2292 4399 2295
rect 4614 2292 4620 2304
rect 4387 2264 4620 2292
rect 4387 2261 4399 2264
rect 4341 2255 4399 2261
rect 4614 2252 4620 2264
rect 4672 2252 4678 2304
rect 4706 2252 4712 2304
rect 4764 2252 4770 2304
rect 5166 2252 5172 2304
rect 5224 2252 5230 2304
rect 7282 2252 7288 2304
rect 7340 2252 7346 2304
rect 9309 2295 9367 2301
rect 9309 2261 9321 2295
rect 9355 2292 9367 2295
rect 10704 2292 10732 2332
rect 9355 2264 10732 2292
rect 10888 2292 10916 2332
rect 24964 2304 24992 2400
rect 25682 2388 25688 2400
rect 25740 2388 25746 2440
rect 27264 2428 27292 2456
rect 27448 2428 27476 2459
rect 27264 2400 27476 2428
rect 25317 2363 25375 2369
rect 25317 2329 25329 2363
rect 25363 2360 25375 2363
rect 25869 2363 25927 2369
rect 25869 2360 25881 2363
rect 25363 2332 25881 2360
rect 25363 2329 25375 2332
rect 25317 2323 25375 2329
rect 25869 2329 25881 2332
rect 25915 2360 25927 2363
rect 26326 2360 26332 2372
rect 25915 2332 26332 2360
rect 25915 2329 25927 2332
rect 25869 2323 25927 2329
rect 26326 2320 26332 2332
rect 26384 2320 26390 2372
rect 14182 2292 14188 2304
rect 10888 2264 14188 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 15562 2252 15568 2304
rect 15620 2292 15626 2304
rect 21729 2295 21787 2301
rect 21729 2292 21741 2295
rect 15620 2264 21741 2292
rect 15620 2252 15626 2264
rect 21729 2261 21741 2264
rect 21775 2261 21787 2295
rect 21729 2255 21787 2261
rect 24305 2295 24363 2301
rect 24305 2261 24317 2295
rect 24351 2292 24363 2295
rect 24486 2292 24492 2304
rect 24351 2264 24492 2292
rect 24351 2261 24363 2264
rect 24305 2255 24363 2261
rect 24486 2252 24492 2264
rect 24544 2292 24550 2304
rect 24946 2292 24952 2304
rect 24544 2264 24952 2292
rect 24544 2252 24550 2264
rect 24946 2252 24952 2264
rect 25004 2252 25010 2304
rect 25406 2252 25412 2304
rect 25464 2292 25470 2304
rect 25590 2292 25596 2304
rect 25464 2264 25596 2292
rect 25464 2252 25470 2264
rect 25590 2252 25596 2264
rect 25648 2252 25654 2304
rect 31018 2252 31024 2304
rect 31076 2252 31082 2304
rect 552 2202 31372 2224
rect 552 2150 4250 2202
rect 4302 2150 4314 2202
rect 4366 2150 4378 2202
rect 4430 2150 4442 2202
rect 4494 2150 4506 2202
rect 4558 2150 11955 2202
rect 12007 2150 12019 2202
rect 12071 2150 12083 2202
rect 12135 2150 12147 2202
rect 12199 2150 12211 2202
rect 12263 2150 19660 2202
rect 19712 2150 19724 2202
rect 19776 2150 19788 2202
rect 19840 2150 19852 2202
rect 19904 2150 19916 2202
rect 19968 2150 27365 2202
rect 27417 2150 27429 2202
rect 27481 2150 27493 2202
rect 27545 2150 27557 2202
rect 27609 2150 27621 2202
rect 27673 2150 31372 2202
rect 552 2128 31372 2150
rect 2682 2048 2688 2100
rect 2740 2048 2746 2100
rect 3326 2048 3332 2100
rect 3384 2048 3390 2100
rect 6365 2091 6423 2097
rect 6365 2057 6377 2091
rect 6411 2088 6423 2091
rect 7190 2088 7196 2100
rect 6411 2060 7196 2088
rect 6411 2057 6423 2060
rect 6365 2051 6423 2057
rect 7190 2048 7196 2060
rect 7248 2048 7254 2100
rect 7469 2091 7527 2097
rect 7469 2057 7481 2091
rect 7515 2088 7527 2091
rect 7834 2088 7840 2100
rect 7515 2060 7840 2088
rect 7515 2057 7527 2060
rect 7469 2051 7527 2057
rect 7834 2048 7840 2060
rect 7892 2088 7898 2100
rect 8113 2091 8171 2097
rect 8113 2088 8125 2091
rect 7892 2060 8125 2088
rect 7892 2048 7898 2060
rect 8113 2057 8125 2060
rect 8159 2088 8171 2091
rect 8202 2088 8208 2100
rect 8159 2060 8208 2088
rect 8159 2057 8171 2060
rect 8113 2051 8171 2057
rect 8202 2048 8208 2060
rect 8260 2048 8266 2100
rect 9674 2048 9680 2100
rect 9732 2048 9738 2100
rect 11146 2088 11152 2100
rect 10796 2060 11152 2088
rect 2700 1952 2728 2048
rect 4706 1980 4712 2032
rect 4764 2020 4770 2032
rect 4985 2023 5043 2029
rect 4985 2020 4997 2023
rect 4764 1992 4997 2020
rect 4764 1980 4770 1992
rect 4985 1989 4997 1992
rect 5031 2020 5043 2023
rect 6822 2020 6828 2032
rect 5031 1992 6828 2020
rect 5031 1989 5043 1992
rect 4985 1983 5043 1989
rect 2700 1924 3280 1952
rect 2774 1844 2780 1896
rect 2832 1844 2838 1896
rect 3252 1893 3280 1924
rect 3237 1887 3295 1893
rect 3237 1853 3249 1887
rect 3283 1853 3295 1887
rect 3237 1847 3295 1853
rect 4614 1844 4620 1896
rect 4672 1844 4678 1896
rect 5166 1893 5172 1896
rect 4709 1887 4767 1893
rect 4709 1853 4721 1887
rect 4755 1884 4767 1887
rect 5053 1887 5111 1893
rect 5053 1884 5065 1887
rect 4755 1856 5065 1884
rect 4755 1853 4767 1856
rect 4709 1847 4767 1853
rect 5053 1853 5065 1856
rect 5099 1886 5111 1887
rect 5161 1886 5172 1893
rect 5099 1858 5172 1886
rect 5099 1856 5120 1858
rect 5099 1853 5111 1856
rect 5053 1847 5111 1853
rect 5161 1847 5172 1858
rect 5224 1884 5230 1896
rect 5224 1856 5261 1884
rect 5166 1844 5172 1847
rect 5224 1844 5230 1856
rect 5442 1844 5448 1896
rect 5500 1844 5506 1896
rect 5920 1893 5948 1992
rect 6822 1980 6828 1992
rect 6880 1980 6886 2032
rect 7006 1980 7012 2032
rect 7064 1980 7070 2032
rect 7282 1980 7288 2032
rect 7340 1980 7346 2032
rect 6089 1955 6147 1961
rect 6089 1921 6101 1955
rect 6135 1952 6147 1955
rect 7024 1952 7052 1980
rect 6135 1924 7052 1952
rect 7300 1952 7328 1980
rect 7300 1924 7788 1952
rect 6135 1921 6147 1924
rect 6089 1915 6147 1921
rect 6564 1893 6592 1924
rect 5905 1887 5963 1893
rect 5905 1853 5917 1887
rect 5951 1853 5963 1887
rect 5905 1847 5963 1853
rect 6181 1887 6239 1893
rect 6181 1853 6193 1887
rect 6227 1884 6239 1887
rect 6273 1887 6331 1893
rect 6273 1884 6285 1887
rect 6227 1856 6285 1884
rect 6227 1853 6239 1856
rect 6181 1847 6239 1853
rect 6273 1853 6285 1856
rect 6319 1853 6331 1887
rect 6273 1847 6331 1853
rect 6549 1887 6607 1893
rect 6549 1853 6561 1887
rect 6595 1853 6607 1887
rect 6549 1847 6607 1853
rect 4632 1816 4660 1844
rect 5460 1816 5488 1844
rect 4632 1788 5488 1816
rect 5537 1819 5595 1825
rect 5537 1785 5549 1819
rect 5583 1816 5595 1819
rect 5813 1819 5871 1825
rect 5813 1816 5825 1819
rect 5583 1788 5825 1816
rect 5583 1785 5595 1788
rect 5537 1779 5595 1785
rect 5813 1785 5825 1788
rect 5859 1816 5871 1819
rect 6196 1816 6224 1847
rect 5859 1788 6224 1816
rect 5859 1785 5871 1788
rect 5813 1779 5871 1785
rect 5261 1751 5319 1757
rect 5261 1717 5273 1751
rect 5307 1748 5319 1751
rect 6564 1748 6592 1847
rect 6822 1844 6828 1896
rect 6880 1844 6886 1896
rect 7760 1893 7788 1924
rect 7285 1887 7343 1893
rect 7285 1853 7297 1887
rect 7331 1884 7343 1887
rect 7377 1887 7435 1893
rect 7377 1884 7389 1887
rect 7331 1856 7389 1884
rect 7331 1853 7343 1856
rect 7285 1847 7343 1853
rect 7377 1853 7389 1856
rect 7423 1853 7435 1887
rect 7377 1847 7435 1853
rect 7745 1887 7803 1893
rect 7745 1853 7757 1887
rect 7791 1884 7803 1887
rect 8021 1887 8079 1893
rect 8021 1884 8033 1887
rect 7791 1856 8033 1884
rect 7791 1853 7803 1856
rect 7745 1847 7803 1853
rect 8021 1853 8033 1856
rect 8067 1853 8079 1887
rect 8021 1847 8079 1853
rect 6641 1819 6699 1825
rect 6641 1785 6653 1819
rect 6687 1816 6699 1819
rect 6917 1819 6975 1825
rect 6917 1816 6929 1819
rect 6687 1788 6929 1816
rect 6687 1785 6699 1788
rect 6641 1779 6699 1785
rect 6917 1785 6929 1788
rect 6963 1816 6975 1819
rect 7300 1816 7328 1847
rect 8110 1844 8116 1896
rect 8168 1884 8174 1896
rect 8389 1887 8447 1893
rect 8389 1884 8401 1887
rect 8168 1856 8401 1884
rect 8168 1844 8174 1856
rect 8389 1853 8401 1856
rect 8435 1853 8447 1887
rect 8389 1847 8447 1853
rect 9490 1844 9496 1896
rect 9548 1884 9554 1896
rect 9585 1887 9643 1893
rect 9585 1884 9597 1887
rect 9548 1856 9597 1884
rect 9548 1844 9554 1856
rect 9585 1853 9597 1856
rect 9631 1884 9643 1887
rect 9692 1884 9720 2048
rect 10796 1961 10824 2060
rect 11146 2048 11152 2060
rect 11204 2088 11210 2100
rect 11514 2088 11520 2100
rect 11204 2060 11520 2088
rect 11204 2048 11210 2060
rect 11514 2048 11520 2060
rect 11572 2048 11578 2100
rect 12161 2091 12219 2097
rect 12161 2057 12173 2091
rect 12207 2088 12219 2091
rect 12986 2088 12992 2100
rect 12207 2060 12992 2088
rect 12207 2057 12219 2060
rect 12161 2051 12219 2057
rect 12986 2048 12992 2060
rect 13044 2048 13050 2100
rect 16114 2048 16120 2100
rect 16172 2088 16178 2100
rect 17129 2091 17187 2097
rect 17129 2088 17141 2091
rect 16172 2060 17141 2088
rect 16172 2048 16178 2060
rect 17129 2057 17141 2060
rect 17175 2088 17187 2091
rect 17954 2088 17960 2100
rect 17175 2060 17960 2088
rect 17175 2057 17187 2060
rect 17129 2051 17187 2057
rect 17954 2048 17960 2060
rect 18012 2048 18018 2100
rect 18049 2091 18107 2097
rect 18049 2057 18061 2091
rect 18095 2088 18107 2091
rect 18230 2088 18236 2100
rect 18095 2060 18236 2088
rect 18095 2057 18107 2060
rect 18049 2051 18107 2057
rect 18230 2048 18236 2060
rect 18288 2048 18294 2100
rect 19797 2091 19855 2097
rect 19797 2057 19809 2091
rect 19843 2088 19855 2091
rect 20073 2091 20131 2097
rect 20073 2088 20085 2091
rect 19843 2060 20085 2088
rect 19843 2057 19855 2060
rect 19797 2051 19855 2057
rect 20073 2057 20085 2060
rect 20119 2088 20131 2091
rect 20162 2088 20168 2100
rect 20119 2060 20168 2088
rect 20119 2057 20131 2060
rect 20073 2051 20131 2057
rect 20162 2048 20168 2060
rect 20220 2048 20226 2100
rect 21729 2091 21787 2097
rect 21729 2057 21741 2091
rect 21775 2088 21787 2091
rect 22002 2088 22008 2100
rect 21775 2060 22008 2088
rect 21775 2057 21787 2060
rect 21729 2051 21787 2057
rect 22002 2048 22008 2060
rect 22060 2048 22066 2100
rect 22370 2048 22376 2100
rect 22428 2048 22434 2100
rect 23937 2091 23995 2097
rect 23937 2057 23949 2091
rect 23983 2088 23995 2091
rect 24118 2088 24124 2100
rect 23983 2060 24124 2088
rect 23983 2057 23995 2060
rect 23937 2051 23995 2057
rect 24118 2048 24124 2060
rect 24176 2088 24182 2100
rect 24213 2091 24271 2097
rect 24213 2088 24225 2091
rect 24176 2060 24225 2088
rect 24176 2048 24182 2060
rect 24213 2057 24225 2060
rect 24259 2057 24271 2091
rect 24213 2051 24271 2057
rect 24486 2048 24492 2100
rect 24544 2048 24550 2100
rect 25133 2091 25191 2097
rect 25133 2088 25145 2091
rect 24826 2060 25145 2088
rect 18248 2020 18276 2048
rect 22388 2020 22416 2048
rect 24826 2020 24854 2060
rect 25133 2057 25145 2060
rect 25179 2057 25191 2091
rect 25133 2051 25191 2057
rect 18248 1992 18644 2020
rect 22388 1992 24854 2020
rect 10781 1955 10839 1961
rect 10781 1921 10793 1955
rect 10827 1921 10839 1955
rect 10781 1915 10839 1921
rect 15289 1955 15347 1961
rect 15289 1921 15301 1955
rect 15335 1952 15347 1955
rect 15841 1955 15899 1961
rect 15841 1952 15853 1955
rect 15335 1924 15853 1952
rect 15335 1921 15347 1924
rect 15289 1915 15347 1921
rect 15841 1921 15853 1924
rect 15887 1952 15899 1955
rect 16850 1952 16856 1964
rect 15887 1924 16856 1952
rect 15887 1921 15899 1924
rect 15841 1915 15899 1921
rect 16850 1912 16856 1924
rect 16908 1952 16914 1964
rect 16908 1924 17356 1952
rect 16908 1912 16914 1924
rect 9631 1856 9720 1884
rect 9631 1853 9643 1856
rect 9585 1847 9643 1853
rect 9858 1844 9864 1896
rect 9916 1844 9922 1896
rect 11606 1844 11612 1896
rect 11664 1884 11670 1896
rect 12437 1887 12495 1893
rect 12437 1884 12449 1887
rect 11664 1856 12449 1884
rect 11664 1844 11670 1856
rect 12437 1853 12449 1856
rect 12483 1884 12495 1887
rect 12529 1887 12587 1893
rect 12529 1884 12541 1887
rect 12483 1856 12541 1884
rect 12483 1853 12495 1856
rect 12437 1847 12495 1853
rect 12529 1853 12541 1856
rect 12575 1853 12587 1887
rect 12529 1847 12587 1853
rect 14553 1887 14611 1893
rect 14553 1853 14565 1887
rect 14599 1853 14611 1887
rect 14553 1847 14611 1853
rect 6963 1788 7328 1816
rect 7837 1819 7895 1825
rect 6963 1785 6975 1788
rect 6917 1779 6975 1785
rect 7837 1785 7849 1819
rect 7883 1816 7895 1819
rect 8481 1819 8539 1825
rect 8481 1816 8493 1819
rect 7883 1788 8493 1816
rect 7883 1785 7895 1788
rect 7837 1779 7895 1785
rect 8481 1785 8493 1788
rect 8527 1816 8539 1819
rect 9876 1816 9904 1844
rect 8527 1788 9904 1816
rect 8527 1785 8539 1788
rect 8481 1779 8539 1785
rect 10594 1776 10600 1828
rect 10652 1816 10658 1828
rect 11026 1819 11084 1825
rect 11026 1816 11038 1819
rect 10652 1788 11038 1816
rect 10652 1776 10658 1788
rect 11026 1785 11038 1788
rect 11072 1785 11084 1819
rect 11026 1779 11084 1785
rect 14568 1760 14596 1847
rect 15194 1844 15200 1896
rect 15252 1844 15258 1896
rect 15470 1884 15476 1896
rect 15433 1856 15476 1884
rect 15470 1844 15476 1856
rect 15528 1844 15534 1896
rect 15565 1887 15623 1893
rect 15565 1853 15577 1887
rect 15611 1884 15623 1887
rect 15654 1884 15660 1896
rect 15611 1856 15660 1884
rect 15611 1853 15623 1856
rect 15565 1847 15623 1853
rect 15654 1844 15660 1856
rect 15712 1884 15718 1896
rect 15749 1887 15807 1893
rect 15749 1884 15761 1887
rect 15712 1856 15761 1884
rect 15712 1844 15718 1856
rect 15749 1853 15761 1856
rect 15795 1884 15807 1887
rect 16025 1887 16083 1893
rect 16025 1884 16037 1887
rect 15795 1856 16037 1884
rect 15795 1853 15807 1856
rect 15749 1847 15807 1853
rect 16025 1853 16037 1856
rect 16071 1853 16083 1887
rect 16025 1847 16083 1853
rect 16298 1844 16304 1896
rect 16356 1844 16362 1896
rect 16960 1893 16988 1924
rect 17328 1893 17356 1924
rect 16945 1887 17003 1893
rect 16945 1853 16957 1887
rect 16991 1853 17003 1887
rect 16945 1847 17003 1853
rect 17045 1887 17103 1893
rect 17045 1853 17057 1887
rect 17091 1884 17103 1887
rect 17313 1887 17371 1893
rect 17091 1856 17172 1884
rect 17091 1853 17103 1856
rect 17045 1847 17103 1853
rect 5307 1720 6592 1748
rect 5307 1717 5319 1720
rect 5261 1711 5319 1717
rect 9398 1708 9404 1760
rect 9456 1708 9462 1760
rect 9674 1708 9680 1760
rect 9732 1708 9738 1760
rect 12342 1708 12348 1760
rect 12400 1708 12406 1760
rect 12618 1708 12624 1760
rect 12676 1708 12682 1760
rect 14458 1708 14464 1760
rect 14516 1708 14522 1760
rect 14550 1708 14556 1760
rect 14608 1708 14614 1760
rect 16393 1751 16451 1757
rect 16393 1717 16405 1751
rect 16439 1748 16451 1751
rect 16850 1748 16856 1760
rect 16439 1720 16856 1748
rect 16439 1717 16451 1720
rect 16393 1711 16451 1717
rect 16850 1708 16856 1720
rect 16908 1748 16914 1760
rect 17144 1748 17172 1856
rect 17313 1853 17325 1887
rect 17359 1853 17371 1887
rect 17313 1847 17371 1853
rect 17405 1887 17463 1893
rect 17405 1853 17417 1887
rect 17451 1884 17463 1887
rect 17954 1884 17960 1896
rect 17451 1856 17960 1884
rect 17451 1853 17463 1856
rect 17405 1847 17463 1853
rect 17954 1844 17960 1856
rect 18012 1844 18018 1896
rect 18233 1887 18291 1893
rect 18233 1853 18245 1887
rect 18279 1853 18291 1887
rect 18616 1884 18644 1992
rect 18690 1912 18696 1964
rect 18748 1952 18754 1964
rect 20070 1952 20076 1964
rect 18748 1924 20076 1952
rect 18748 1912 18754 1924
rect 20070 1912 20076 1924
rect 20128 1952 20134 1964
rect 20349 1955 20407 1961
rect 20349 1952 20361 1955
rect 20128 1924 20361 1952
rect 20128 1912 20134 1924
rect 20349 1921 20361 1924
rect 20395 1921 20407 1955
rect 20349 1915 20407 1921
rect 23569 1955 23627 1961
rect 23569 1921 23581 1955
rect 23615 1952 23627 1955
rect 24486 1952 24492 1964
rect 23615 1924 24492 1952
rect 23615 1921 23627 1924
rect 23569 1915 23627 1921
rect 24486 1912 24492 1924
rect 24544 1952 24550 1964
rect 24544 1924 24624 1952
rect 24544 1912 24550 1924
rect 19058 1884 19064 1896
rect 18616 1856 19064 1884
rect 18233 1847 18291 1853
rect 17586 1776 17592 1828
rect 17644 1816 17650 1828
rect 18248 1816 18276 1847
rect 19058 1844 19064 1856
rect 19116 1884 19122 1896
rect 19705 1887 19763 1893
rect 19705 1884 19717 1887
rect 19116 1856 19717 1884
rect 19116 1844 19122 1856
rect 19705 1853 19717 1856
rect 19751 1853 19763 1887
rect 19705 1847 19763 1853
rect 19981 1887 20039 1893
rect 19981 1853 19993 1887
rect 20027 1853 20039 1887
rect 19981 1847 20039 1853
rect 22005 1887 22063 1893
rect 22005 1853 22017 1887
rect 22051 1884 22063 1887
rect 22051 1856 22140 1884
rect 22051 1853 22063 1856
rect 22005 1847 22063 1853
rect 17644 1788 19334 1816
rect 17644 1776 17650 1788
rect 16908 1720 17172 1748
rect 18325 1751 18383 1757
rect 16908 1708 16914 1720
rect 18325 1717 18337 1751
rect 18371 1748 18383 1751
rect 18782 1748 18788 1760
rect 18371 1720 18788 1748
rect 18371 1717 18383 1720
rect 18325 1711 18383 1717
rect 18782 1708 18788 1720
rect 18840 1708 18846 1760
rect 19306 1748 19334 1788
rect 19426 1776 19432 1828
rect 19484 1816 19490 1828
rect 19996 1816 20024 1847
rect 19484 1788 20024 1816
rect 19484 1776 19490 1788
rect 20438 1776 20444 1828
rect 20496 1816 20502 1828
rect 20594 1819 20652 1825
rect 20594 1816 20606 1819
rect 20496 1788 20606 1816
rect 20496 1776 20502 1788
rect 20594 1785 20606 1788
rect 20640 1785 20652 1819
rect 20594 1779 20652 1785
rect 22112 1760 22140 1856
rect 22830 1844 22836 1896
rect 22888 1884 22894 1896
rect 24596 1893 24624 1924
rect 25130 1912 25136 1964
rect 25188 1912 25194 1964
rect 23477 1887 23535 1893
rect 23477 1884 23489 1887
rect 22888 1856 23489 1884
rect 22888 1844 22894 1856
rect 23477 1853 23489 1856
rect 23523 1884 23535 1887
rect 23845 1887 23903 1893
rect 23845 1884 23857 1887
rect 23523 1856 23857 1884
rect 23523 1853 23535 1856
rect 23477 1847 23535 1853
rect 23845 1853 23857 1856
rect 23891 1853 23903 1887
rect 24305 1887 24363 1893
rect 24305 1884 24317 1887
rect 23845 1847 23903 1853
rect 24228 1856 24317 1884
rect 24228 1816 24256 1856
rect 24305 1853 24317 1856
rect 24351 1853 24363 1887
rect 24305 1847 24363 1853
rect 24581 1887 24639 1893
rect 24581 1853 24593 1887
rect 24627 1884 24639 1887
rect 24673 1887 24731 1893
rect 24673 1884 24685 1887
rect 24627 1856 24685 1884
rect 24627 1853 24639 1856
rect 24581 1847 24639 1853
rect 24673 1853 24685 1856
rect 24719 1853 24731 1887
rect 25148 1884 25176 1912
rect 26513 1887 26571 1893
rect 26513 1884 26525 1887
rect 25148 1856 26525 1884
rect 24673 1847 24731 1853
rect 26513 1853 26525 1856
rect 26559 1853 26571 1887
rect 26513 1847 26571 1853
rect 31018 1844 31024 1896
rect 31076 1844 31082 1896
rect 24765 1819 24823 1825
rect 24765 1816 24777 1819
rect 24228 1788 24777 1816
rect 24228 1760 24256 1788
rect 24765 1785 24777 1788
rect 24811 1816 24823 1819
rect 26246 1819 26304 1825
rect 26246 1816 26258 1819
rect 24811 1788 26258 1816
rect 24811 1785 24823 1788
rect 24765 1779 24823 1785
rect 26246 1785 26258 1788
rect 26292 1785 26304 1819
rect 26246 1779 26304 1785
rect 19518 1748 19524 1760
rect 19306 1720 19524 1748
rect 19518 1708 19524 1720
rect 19576 1708 19582 1760
rect 21913 1751 21971 1757
rect 21913 1717 21925 1751
rect 21959 1748 21971 1751
rect 22002 1748 22008 1760
rect 21959 1720 22008 1748
rect 21959 1717 21971 1720
rect 21913 1711 21971 1717
rect 22002 1708 22008 1720
rect 22060 1708 22066 1760
rect 22094 1708 22100 1760
rect 22152 1708 22158 1760
rect 24210 1708 24216 1760
rect 24268 1708 24274 1760
rect 552 1658 31531 1680
rect 552 1606 8102 1658
rect 8154 1606 8166 1658
rect 8218 1606 8230 1658
rect 8282 1606 8294 1658
rect 8346 1606 8358 1658
rect 8410 1606 15807 1658
rect 15859 1606 15871 1658
rect 15923 1606 15935 1658
rect 15987 1606 15999 1658
rect 16051 1606 16063 1658
rect 16115 1606 23512 1658
rect 23564 1606 23576 1658
rect 23628 1606 23640 1658
rect 23692 1606 23704 1658
rect 23756 1606 23768 1658
rect 23820 1606 31217 1658
rect 31269 1606 31281 1658
rect 31333 1606 31345 1658
rect 31397 1606 31409 1658
rect 31461 1606 31473 1658
rect 31525 1606 31531 1658
rect 552 1584 31531 1606
rect 7190 1504 7196 1556
rect 7248 1504 7254 1556
rect 7282 1504 7288 1556
rect 7340 1544 7346 1556
rect 7377 1547 7435 1553
rect 7377 1544 7389 1547
rect 7340 1516 7389 1544
rect 7340 1504 7346 1516
rect 7377 1513 7389 1516
rect 7423 1513 7435 1547
rect 7377 1507 7435 1513
rect 7834 1504 7840 1556
rect 7892 1504 7898 1556
rect 8205 1547 8263 1553
rect 8205 1513 8217 1547
rect 8251 1544 8263 1547
rect 9490 1544 9496 1556
rect 8251 1516 9496 1544
rect 8251 1513 8263 1516
rect 8205 1507 8263 1513
rect 7208 1408 7236 1504
rect 7852 1417 7880 1504
rect 8478 1476 8484 1488
rect 8128 1448 8484 1476
rect 8128 1417 8156 1448
rect 8478 1436 8484 1448
rect 8536 1476 8542 1488
rect 8536 1448 8708 1476
rect 8536 1436 8542 1448
rect 8680 1417 8708 1448
rect 7469 1411 7527 1417
rect 7469 1408 7481 1411
rect 7208 1380 7481 1408
rect 7469 1377 7481 1380
rect 7515 1408 7527 1411
rect 7561 1411 7619 1417
rect 7561 1408 7573 1411
rect 7515 1380 7573 1408
rect 7515 1377 7527 1380
rect 7469 1371 7527 1377
rect 7561 1377 7573 1380
rect 7607 1377 7619 1411
rect 7561 1371 7619 1377
rect 7837 1411 7895 1417
rect 7837 1377 7849 1411
rect 7883 1377 7895 1411
rect 7837 1371 7895 1377
rect 7929 1411 7987 1417
rect 7929 1377 7941 1411
rect 7975 1408 7987 1411
rect 8113 1411 8171 1417
rect 8113 1408 8125 1411
rect 7975 1380 8125 1408
rect 7975 1377 7987 1380
rect 7929 1371 7987 1377
rect 8113 1377 8125 1380
rect 8159 1377 8171 1411
rect 8389 1411 8447 1417
rect 8389 1408 8401 1411
rect 8113 1371 8171 1377
rect 8220 1380 8401 1408
rect 7653 1343 7711 1349
rect 7653 1309 7665 1343
rect 7699 1340 7711 1343
rect 8018 1340 8024 1352
rect 7699 1312 8024 1340
rect 7699 1309 7711 1312
rect 7653 1303 7711 1309
rect 8018 1300 8024 1312
rect 8076 1340 8082 1352
rect 8220 1340 8248 1380
rect 8389 1377 8401 1380
rect 8435 1377 8447 1411
rect 8389 1371 8447 1377
rect 8665 1411 8723 1417
rect 8665 1377 8677 1411
rect 8711 1377 8723 1411
rect 8665 1371 8723 1377
rect 8076 1312 8248 1340
rect 8481 1343 8539 1349
rect 8076 1300 8082 1312
rect 8481 1309 8493 1343
rect 8527 1340 8539 1343
rect 8772 1340 8800 1516
rect 9490 1504 9496 1516
rect 9548 1504 9554 1556
rect 9861 1547 9919 1553
rect 9861 1513 9873 1547
rect 9907 1544 9919 1547
rect 10137 1547 10195 1553
rect 10137 1544 10149 1547
rect 9907 1516 10149 1544
rect 9907 1513 9919 1516
rect 9861 1507 9919 1513
rect 10137 1513 10149 1516
rect 10183 1544 10195 1547
rect 10183 1516 11376 1544
rect 10183 1513 10195 1516
rect 10137 1507 10195 1513
rect 9398 1476 9404 1488
rect 9232 1448 9404 1476
rect 9232 1417 9260 1448
rect 9398 1436 9404 1448
rect 9456 1436 9462 1488
rect 10413 1479 10471 1485
rect 10413 1445 10425 1479
rect 10459 1476 10471 1479
rect 10689 1479 10747 1485
rect 10689 1476 10701 1479
rect 10459 1448 10701 1476
rect 10459 1445 10471 1448
rect 10413 1439 10471 1445
rect 10689 1445 10701 1448
rect 10735 1476 10747 1479
rect 10735 1448 11008 1476
rect 10735 1445 10747 1448
rect 10689 1439 10747 1445
rect 9033 1411 9091 1417
rect 9033 1377 9045 1411
rect 9079 1377 9091 1411
rect 9033 1371 9091 1377
rect 9125 1411 9183 1417
rect 9125 1377 9137 1411
rect 9171 1408 9183 1411
rect 9217 1411 9275 1417
rect 9217 1408 9229 1411
rect 9171 1380 9229 1408
rect 9171 1377 9183 1380
rect 9125 1371 9183 1377
rect 9217 1377 9229 1380
rect 9263 1377 9275 1411
rect 9217 1371 9275 1377
rect 8527 1312 8800 1340
rect 9048 1340 9076 1371
rect 9674 1368 9680 1420
rect 9732 1408 9738 1420
rect 9769 1411 9827 1417
rect 9769 1408 9781 1411
rect 9732 1380 9781 1408
rect 9732 1368 9738 1380
rect 9769 1377 9781 1380
rect 9815 1377 9827 1411
rect 9769 1371 9827 1377
rect 10229 1411 10287 1417
rect 10229 1377 10241 1411
rect 10275 1408 10287 1411
rect 10428 1408 10456 1439
rect 10275 1380 10456 1408
rect 10505 1411 10563 1417
rect 10275 1377 10287 1380
rect 10229 1371 10287 1377
rect 10505 1377 10517 1411
rect 10551 1408 10563 1411
rect 10594 1408 10600 1420
rect 10551 1380 10600 1408
rect 10551 1377 10563 1380
rect 10505 1371 10563 1377
rect 10520 1340 10548 1371
rect 10594 1368 10600 1380
rect 10652 1368 10658 1420
rect 10980 1417 11008 1448
rect 11054 1436 11060 1488
rect 11112 1436 11118 1488
rect 11146 1436 11152 1488
rect 11204 1436 11210 1488
rect 10781 1411 10839 1417
rect 10781 1408 10793 1411
rect 10704 1380 10793 1408
rect 9048 1312 10548 1340
rect 8527 1309 8539 1312
rect 8481 1303 8539 1309
rect 8757 1275 8815 1281
rect 8757 1241 8769 1275
rect 8803 1272 8815 1275
rect 9048 1272 9076 1312
rect 8803 1244 9076 1272
rect 9309 1275 9367 1281
rect 8803 1241 8815 1244
rect 8757 1235 8815 1241
rect 9309 1241 9321 1275
rect 9355 1272 9367 1275
rect 9585 1275 9643 1281
rect 9585 1272 9597 1275
rect 9355 1244 9597 1272
rect 9355 1241 9367 1244
rect 9309 1235 9367 1241
rect 9585 1241 9597 1244
rect 9631 1272 9643 1275
rect 10704 1272 10732 1380
rect 10781 1377 10793 1380
rect 10827 1408 10839 1411
rect 10965 1411 11023 1417
rect 10827 1380 10916 1408
rect 10827 1377 10839 1380
rect 10781 1371 10839 1377
rect 10888 1340 10916 1380
rect 10965 1377 10977 1411
rect 11011 1377 11023 1411
rect 11164 1408 11192 1436
rect 11241 1411 11299 1417
rect 11241 1408 11253 1411
rect 11164 1380 11253 1408
rect 10965 1371 11023 1377
rect 11241 1377 11253 1380
rect 11287 1377 11299 1411
rect 11348 1408 11376 1516
rect 11606 1504 11612 1556
rect 11664 1504 11670 1556
rect 12621 1547 12679 1553
rect 12621 1513 12633 1547
rect 12667 1544 12679 1547
rect 12802 1544 12808 1556
rect 12667 1516 12808 1544
rect 12667 1513 12679 1516
rect 12621 1507 12679 1513
rect 12802 1504 12808 1516
rect 12860 1504 12866 1556
rect 13081 1547 13139 1553
rect 13081 1513 13093 1547
rect 13127 1544 13139 1547
rect 13170 1544 13176 1556
rect 13127 1516 13176 1544
rect 13127 1513 13139 1516
rect 13081 1507 13139 1513
rect 13170 1504 13176 1516
rect 13228 1544 13234 1556
rect 13909 1547 13967 1553
rect 13909 1544 13921 1547
rect 13228 1516 13921 1544
rect 13228 1504 13234 1516
rect 13909 1513 13921 1516
rect 13955 1544 13967 1547
rect 14550 1544 14556 1556
rect 13955 1516 14556 1544
rect 13955 1513 13967 1516
rect 13909 1507 13967 1513
rect 14550 1504 14556 1516
rect 14608 1544 14614 1556
rect 14608 1516 14688 1544
rect 14608 1504 14614 1516
rect 11508 1411 11566 1417
rect 11508 1408 11520 1411
rect 11348 1380 11520 1408
rect 11241 1371 11299 1377
rect 11508 1377 11520 1380
rect 11554 1408 11566 1411
rect 11624 1408 11652 1504
rect 13357 1479 13415 1485
rect 13357 1445 13369 1479
rect 13403 1476 13415 1479
rect 13403 1448 13676 1476
rect 13403 1445 13415 1448
rect 13357 1439 13415 1445
rect 11554 1380 11652 1408
rect 11554 1377 11566 1380
rect 11508 1371 11566 1377
rect 12618 1368 12624 1420
rect 12676 1408 12682 1420
rect 12713 1411 12771 1417
rect 12713 1408 12725 1411
rect 12676 1380 12725 1408
rect 12676 1368 12682 1380
rect 12713 1377 12725 1380
rect 12759 1408 12771 1411
rect 12989 1411 13047 1417
rect 12989 1408 13001 1411
rect 12759 1380 13001 1408
rect 12759 1377 12771 1380
rect 12713 1371 12771 1377
rect 12989 1377 13001 1380
rect 13035 1377 13047 1411
rect 12989 1371 13047 1377
rect 13170 1368 13176 1420
rect 13228 1408 13234 1420
rect 13648 1417 13676 1448
rect 14458 1436 14464 1488
rect 14516 1436 14522 1488
rect 13265 1411 13323 1417
rect 13265 1408 13277 1411
rect 13228 1380 13277 1408
rect 13228 1368 13234 1380
rect 13265 1377 13277 1380
rect 13311 1377 13323 1411
rect 13265 1371 13323 1377
rect 13541 1411 13599 1417
rect 13541 1377 13553 1411
rect 13587 1377 13599 1411
rect 13541 1371 13599 1377
rect 13633 1411 13691 1417
rect 13633 1377 13645 1411
rect 13679 1408 13691 1411
rect 14001 1411 14059 1417
rect 14001 1408 14013 1411
rect 13679 1380 14013 1408
rect 13679 1377 13691 1380
rect 13633 1371 13691 1377
rect 14001 1377 14013 1380
rect 14047 1377 14059 1411
rect 14001 1371 14059 1377
rect 14277 1411 14335 1417
rect 14277 1377 14289 1411
rect 14323 1408 14335 1411
rect 14369 1411 14427 1417
rect 14369 1408 14381 1411
rect 14323 1380 14381 1408
rect 14323 1377 14335 1380
rect 14277 1371 14335 1377
rect 14369 1377 14381 1380
rect 14415 1408 14427 1411
rect 14476 1408 14504 1436
rect 14660 1417 14688 1516
rect 14734 1504 14740 1556
rect 14792 1544 14798 1556
rect 15470 1544 15476 1556
rect 14792 1516 15476 1544
rect 14792 1504 14798 1516
rect 15194 1436 15200 1488
rect 15252 1436 15258 1488
rect 15304 1476 15332 1516
rect 15470 1504 15476 1516
rect 15528 1504 15534 1556
rect 15654 1504 15660 1556
rect 15712 1544 15718 1556
rect 15841 1547 15899 1553
rect 15841 1544 15853 1547
rect 15712 1516 15853 1544
rect 15712 1504 15718 1516
rect 15841 1513 15853 1516
rect 15887 1513 15899 1547
rect 15841 1507 15899 1513
rect 16298 1504 16304 1556
rect 16356 1504 16362 1556
rect 16390 1504 16396 1556
rect 16448 1504 16454 1556
rect 16850 1504 16856 1556
rect 16908 1504 16914 1556
rect 17313 1547 17371 1553
rect 17313 1513 17325 1547
rect 17359 1544 17371 1547
rect 17586 1544 17592 1556
rect 17359 1516 17592 1544
rect 17359 1513 17371 1516
rect 17313 1507 17371 1513
rect 17586 1504 17592 1516
rect 17644 1504 17650 1556
rect 17681 1547 17739 1553
rect 17681 1513 17693 1547
rect 17727 1544 17739 1547
rect 17770 1544 17776 1556
rect 17727 1516 17776 1544
rect 17727 1513 17739 1516
rect 17681 1507 17739 1513
rect 17770 1504 17776 1516
rect 17828 1504 17834 1556
rect 17954 1504 17960 1556
rect 18012 1504 18018 1556
rect 18046 1504 18052 1556
rect 18104 1504 18110 1556
rect 18506 1504 18512 1556
rect 18564 1504 18570 1556
rect 18782 1504 18788 1556
rect 18840 1504 18846 1556
rect 19058 1504 19064 1556
rect 19116 1504 19122 1556
rect 19337 1547 19395 1553
rect 19337 1513 19349 1547
rect 19383 1544 19395 1547
rect 19426 1544 19432 1556
rect 19383 1516 19432 1544
rect 19383 1513 19395 1516
rect 19337 1507 19395 1513
rect 19426 1504 19432 1516
rect 19484 1544 19490 1556
rect 20070 1544 20076 1556
rect 19484 1516 20076 1544
rect 19484 1504 19490 1516
rect 20070 1504 20076 1516
rect 20128 1544 20134 1556
rect 20165 1547 20223 1553
rect 20165 1544 20177 1547
rect 20128 1516 20177 1544
rect 20128 1504 20134 1516
rect 20165 1513 20177 1516
rect 20211 1513 20223 1547
rect 20165 1507 20223 1513
rect 20254 1504 20260 1556
rect 20312 1544 20318 1556
rect 20717 1547 20775 1553
rect 20717 1544 20729 1547
rect 20312 1516 20729 1544
rect 20312 1504 20318 1516
rect 20717 1513 20729 1516
rect 20763 1513 20775 1547
rect 20717 1507 20775 1513
rect 16316 1476 16344 1504
rect 15304 1448 16344 1476
rect 16868 1476 16896 1504
rect 16868 1448 17264 1476
rect 14415 1380 14504 1408
rect 14645 1411 14703 1417
rect 14415 1377 14427 1380
rect 14369 1371 14427 1377
rect 14645 1377 14657 1411
rect 14691 1377 14703 1411
rect 14645 1371 14703 1377
rect 14737 1411 14795 1417
rect 14737 1377 14749 1411
rect 14783 1408 14795 1411
rect 15212 1408 15240 1436
rect 15289 1411 15347 1417
rect 15289 1408 15301 1411
rect 14783 1380 15301 1408
rect 14783 1377 14795 1380
rect 14737 1371 14795 1377
rect 15289 1377 15301 1380
rect 15335 1408 15347 1411
rect 15473 1411 15531 1417
rect 15473 1408 15485 1411
rect 15335 1380 15485 1408
rect 15335 1377 15347 1380
rect 15289 1371 15347 1377
rect 15473 1377 15485 1380
rect 15519 1377 15531 1411
rect 15473 1371 15531 1377
rect 15565 1411 15623 1417
rect 15565 1377 15577 1411
rect 15611 1408 15623 1411
rect 15933 1411 15991 1417
rect 15933 1408 15945 1411
rect 15611 1380 15945 1408
rect 15611 1377 15623 1380
rect 15565 1371 15623 1377
rect 15933 1377 15945 1380
rect 15979 1377 15991 1411
rect 15933 1371 15991 1377
rect 12805 1343 12863 1349
rect 10888 1312 11100 1340
rect 9631 1244 10732 1272
rect 9631 1241 9643 1244
rect 9585 1235 9643 1241
rect 11072 1204 11100 1312
rect 12805 1309 12817 1343
rect 12851 1340 12863 1343
rect 13556 1340 13584 1371
rect 13722 1340 13728 1352
rect 12851 1312 13728 1340
rect 12851 1309 12863 1312
rect 12805 1303 12863 1309
rect 13722 1300 13728 1312
rect 13780 1300 13786 1352
rect 14016 1340 14044 1371
rect 15580 1340 15608 1371
rect 14016 1312 14688 1340
rect 14366 1232 14372 1284
rect 14424 1272 14430 1284
rect 14461 1275 14519 1281
rect 14461 1272 14473 1275
rect 14424 1244 14473 1272
rect 14424 1232 14430 1244
rect 14461 1241 14473 1244
rect 14507 1241 14519 1275
rect 14461 1235 14519 1241
rect 14660 1216 14688 1312
rect 14752 1312 15608 1340
rect 14752 1216 14780 1312
rect 15197 1275 15255 1281
rect 15197 1241 15209 1275
rect 15243 1272 15255 1275
rect 16031 1272 16059 1448
rect 16209 1411 16267 1417
rect 16209 1377 16221 1411
rect 16255 1408 16267 1411
rect 16298 1408 16304 1420
rect 16255 1380 16304 1408
rect 16255 1377 16267 1380
rect 16209 1371 16267 1377
rect 16298 1368 16304 1380
rect 16356 1368 16362 1420
rect 17236 1417 17264 1448
rect 17129 1411 17187 1417
rect 17129 1377 17141 1411
rect 17175 1377 17187 1411
rect 17129 1371 17187 1377
rect 17221 1411 17279 1417
rect 17221 1377 17233 1411
rect 17267 1377 17279 1411
rect 17221 1371 17279 1377
rect 17144 1340 17172 1371
rect 17494 1368 17500 1420
rect 17552 1368 17558 1420
rect 17972 1340 18000 1504
rect 18064 1476 18092 1504
rect 18064 1448 18736 1476
rect 18064 1417 18092 1448
rect 18049 1411 18107 1417
rect 18049 1377 18061 1411
rect 18095 1377 18107 1411
rect 18049 1371 18107 1377
rect 18230 1368 18236 1420
rect 18288 1368 18294 1420
rect 18708 1417 18736 1448
rect 18693 1411 18751 1417
rect 18693 1377 18705 1411
rect 18739 1377 18751 1411
rect 18800 1408 18828 1504
rect 19076 1476 19104 1504
rect 20732 1476 20760 1507
rect 22002 1504 22008 1556
rect 22060 1544 22066 1556
rect 22462 1544 22468 1556
rect 22060 1516 22468 1544
rect 22060 1504 22066 1516
rect 22462 1504 22468 1516
rect 22520 1504 22526 1556
rect 22741 1547 22799 1553
rect 22741 1513 22753 1547
rect 22787 1544 22799 1547
rect 22830 1544 22836 1556
rect 22787 1516 22836 1544
rect 22787 1513 22799 1516
rect 22741 1507 22799 1513
rect 22830 1504 22836 1516
rect 22888 1544 22894 1556
rect 23477 1547 23535 1553
rect 23477 1544 23489 1547
rect 22888 1516 23489 1544
rect 22888 1504 22894 1516
rect 23477 1513 23489 1516
rect 23523 1513 23535 1547
rect 23477 1507 23535 1513
rect 23753 1547 23811 1553
rect 23753 1513 23765 1547
rect 23799 1544 23811 1547
rect 23842 1544 23848 1556
rect 23799 1516 23848 1544
rect 23799 1513 23811 1516
rect 23753 1507 23811 1513
rect 23842 1504 23848 1516
rect 23900 1504 23906 1556
rect 25406 1504 25412 1556
rect 25464 1504 25470 1556
rect 19076 1448 19840 1476
rect 19153 1411 19211 1417
rect 19153 1408 19165 1411
rect 18800 1380 19165 1408
rect 18693 1371 18751 1377
rect 19153 1377 19165 1380
rect 19199 1408 19211 1411
rect 19245 1411 19303 1417
rect 19245 1408 19257 1411
rect 19199 1380 19257 1408
rect 19199 1377 19211 1380
rect 19153 1371 19211 1377
rect 19245 1377 19257 1380
rect 19291 1377 19303 1411
rect 19245 1371 19303 1377
rect 19518 1368 19524 1420
rect 19576 1368 19582 1420
rect 19812 1417 19840 1448
rect 20272 1448 20668 1476
rect 20732 1448 21496 1476
rect 20272 1417 20300 1448
rect 19797 1411 19855 1417
rect 19797 1377 19809 1411
rect 19843 1377 19855 1411
rect 20257 1411 20315 1417
rect 20257 1408 20269 1411
rect 19797 1371 19855 1377
rect 19904 1380 20269 1408
rect 17144 1312 18000 1340
rect 15243 1244 16059 1272
rect 17037 1275 17095 1281
rect 15243 1241 15255 1244
rect 15197 1235 15255 1241
rect 17037 1241 17049 1275
rect 17083 1272 17095 1275
rect 17586 1272 17592 1284
rect 17083 1244 17592 1272
rect 17083 1241 17095 1244
rect 17037 1235 17095 1241
rect 17586 1232 17592 1244
rect 17644 1232 17650 1284
rect 19904 1281 19932 1380
rect 20257 1377 20269 1380
rect 20303 1377 20315 1411
rect 20257 1371 20315 1377
rect 20349 1411 20407 1417
rect 20349 1377 20361 1411
rect 20395 1377 20407 1411
rect 20349 1371 20407 1377
rect 20162 1300 20168 1352
rect 20220 1340 20226 1352
rect 20364 1340 20392 1371
rect 20438 1368 20444 1420
rect 20496 1368 20502 1420
rect 20640 1417 20668 1448
rect 21468 1417 21496 1448
rect 24210 1436 24216 1488
rect 24268 1476 24274 1488
rect 24268 1448 25360 1476
rect 24268 1436 24274 1448
rect 20625 1411 20683 1417
rect 20625 1377 20637 1411
rect 20671 1377 20683 1411
rect 20625 1371 20683 1377
rect 20901 1411 20959 1417
rect 20901 1377 20913 1411
rect 20947 1377 20959 1411
rect 20901 1371 20959 1377
rect 21453 1411 21511 1417
rect 21453 1377 21465 1411
rect 21499 1408 21511 1411
rect 21545 1411 21603 1417
rect 21545 1408 21557 1411
rect 21499 1380 21557 1408
rect 21499 1377 21511 1380
rect 21453 1371 21511 1377
rect 21545 1377 21557 1380
rect 21591 1377 21603 1411
rect 21545 1371 21603 1377
rect 20220 1312 20392 1340
rect 20220 1300 20226 1312
rect 19613 1275 19671 1281
rect 19613 1241 19625 1275
rect 19659 1272 19671 1275
rect 19889 1275 19947 1281
rect 19889 1272 19901 1275
rect 19659 1244 19901 1272
rect 19659 1241 19671 1244
rect 19613 1235 19671 1241
rect 19889 1241 19901 1244
rect 19935 1241 19947 1275
rect 19889 1235 19947 1241
rect 20070 1232 20076 1284
rect 20128 1272 20134 1284
rect 20916 1272 20944 1371
rect 21818 1368 21824 1420
rect 21876 1408 21882 1420
rect 22097 1411 22155 1417
rect 22097 1408 22109 1411
rect 21876 1380 22109 1408
rect 21876 1368 21882 1380
rect 22097 1377 22109 1380
rect 22143 1377 22155 1411
rect 22097 1371 22155 1377
rect 22373 1411 22431 1417
rect 22373 1377 22385 1411
rect 22419 1377 22431 1411
rect 22373 1371 22431 1377
rect 22649 1411 22707 1417
rect 22649 1377 22661 1411
rect 22695 1377 22707 1411
rect 22649 1371 22707 1377
rect 21637 1343 21695 1349
rect 21637 1309 21649 1343
rect 21683 1340 21695 1343
rect 21726 1340 21732 1352
rect 21683 1312 21732 1340
rect 21683 1309 21695 1312
rect 21637 1303 21695 1309
rect 21726 1300 21732 1312
rect 21784 1340 21790 1352
rect 21913 1343 21971 1349
rect 21913 1340 21925 1343
rect 21784 1312 21925 1340
rect 21784 1300 21790 1312
rect 21913 1309 21925 1312
rect 21959 1340 21971 1343
rect 22388 1340 22416 1371
rect 21959 1312 22416 1340
rect 21959 1309 21971 1312
rect 21913 1303 21971 1309
rect 22664 1272 22692 1371
rect 22922 1368 22928 1420
rect 22980 1368 22986 1420
rect 23017 1411 23075 1417
rect 23017 1377 23029 1411
rect 23063 1408 23075 1411
rect 23566 1408 23572 1420
rect 23063 1380 23572 1408
rect 23063 1377 23075 1380
rect 23017 1371 23075 1377
rect 23566 1368 23572 1380
rect 23624 1368 23630 1420
rect 24578 1368 24584 1420
rect 24636 1408 24642 1420
rect 24866 1411 24924 1417
rect 24866 1408 24878 1411
rect 24636 1380 24878 1408
rect 24636 1368 24642 1380
rect 24866 1377 24878 1380
rect 24912 1377 24924 1411
rect 24866 1371 24924 1377
rect 25130 1368 25136 1420
rect 25188 1368 25194 1420
rect 25332 1417 25360 1448
rect 25317 1411 25375 1417
rect 25317 1377 25329 1411
rect 25363 1377 25375 1411
rect 25317 1371 25375 1377
rect 20128 1244 20944 1272
rect 22204 1244 22692 1272
rect 20128 1232 20134 1244
rect 11606 1204 11612 1216
rect 11072 1176 11612 1204
rect 11606 1164 11612 1176
rect 11664 1164 11670 1216
rect 14182 1164 14188 1216
rect 14240 1164 14246 1216
rect 14642 1164 14648 1216
rect 14700 1164 14706 1216
rect 14734 1164 14740 1216
rect 14792 1164 14798 1216
rect 20993 1207 21051 1213
rect 20993 1173 21005 1207
rect 21039 1204 21051 1207
rect 21266 1204 21272 1216
rect 21039 1176 21272 1204
rect 21039 1173 21051 1176
rect 20993 1167 21051 1173
rect 21266 1164 21272 1176
rect 21324 1204 21330 1216
rect 21361 1207 21419 1213
rect 21361 1204 21373 1207
rect 21324 1176 21373 1204
rect 21324 1164 21330 1176
rect 21361 1173 21373 1176
rect 21407 1173 21419 1207
rect 21361 1167 21419 1173
rect 22094 1164 22100 1216
rect 22152 1204 22158 1216
rect 22204 1213 22232 1244
rect 22189 1207 22247 1213
rect 22189 1204 22201 1207
rect 22152 1176 22201 1204
rect 22152 1164 22158 1176
rect 22189 1173 22201 1176
rect 22235 1173 22247 1207
rect 22189 1167 22247 1173
rect 552 1114 31372 1136
rect 552 1062 4250 1114
rect 4302 1062 4314 1114
rect 4366 1062 4378 1114
rect 4430 1062 4442 1114
rect 4494 1062 4506 1114
rect 4558 1062 11955 1114
rect 12007 1062 12019 1114
rect 12071 1062 12083 1114
rect 12135 1062 12147 1114
rect 12199 1062 12211 1114
rect 12263 1062 19660 1114
rect 19712 1062 19724 1114
rect 19776 1062 19788 1114
rect 19840 1062 19852 1114
rect 19904 1062 19916 1114
rect 19968 1062 27365 1114
rect 27417 1062 27429 1114
rect 27481 1062 27493 1114
rect 27545 1062 27557 1114
rect 27609 1062 27621 1114
rect 27673 1062 31372 1114
rect 552 1040 31372 1062
rect 8018 960 8024 1012
rect 8076 1000 8082 1012
rect 8113 1003 8171 1009
rect 8113 1000 8125 1003
rect 8076 972 8125 1000
rect 8076 960 8082 972
rect 8113 969 8125 972
rect 8159 969 8171 1003
rect 8113 963 8171 969
rect 8478 960 8484 1012
rect 8536 960 8542 1012
rect 9398 960 9404 1012
rect 9456 960 9462 1012
rect 9674 960 9680 1012
rect 9732 1000 9738 1012
rect 9861 1003 9919 1009
rect 9861 1000 9873 1003
rect 9732 972 9873 1000
rect 9732 960 9738 972
rect 9861 969 9873 972
rect 9907 969 9919 1003
rect 9861 963 9919 969
rect 11054 960 11060 1012
rect 11112 1000 11118 1012
rect 12253 1003 12311 1009
rect 12253 1000 12265 1003
rect 11112 972 12265 1000
rect 11112 960 11118 972
rect 12253 969 12265 972
rect 12299 1000 12311 1003
rect 12299 972 12434 1000
rect 12299 969 12311 972
rect 12253 963 12311 969
rect 11698 892 11704 944
rect 11756 892 11762 944
rect 9858 824 9864 876
rect 9916 824 9922 876
rect 7834 756 7840 808
rect 7892 796 7898 808
rect 8021 799 8079 805
rect 8021 796 8033 799
rect 7892 768 8033 796
rect 7892 756 7898 768
rect 8021 765 8033 768
rect 8067 765 8079 799
rect 8021 759 8079 765
rect 8573 799 8631 805
rect 8573 765 8585 799
rect 8619 796 8631 799
rect 9493 799 9551 805
rect 9493 796 9505 799
rect 8619 768 9505 796
rect 8619 765 8631 768
rect 8573 759 8631 765
rect 9493 765 9505 768
rect 9539 796 9551 799
rect 9876 796 9904 824
rect 9539 768 9904 796
rect 9953 799 10011 805
rect 9539 765 9551 768
rect 9493 759 9551 765
rect 9953 765 9965 799
rect 9999 796 10011 799
rect 10594 796 10600 808
rect 9999 768 10600 796
rect 9999 765 10011 768
rect 9953 759 10011 765
rect 10594 756 10600 768
rect 10652 756 10658 808
rect 11716 796 11744 892
rect 12406 864 12434 972
rect 12618 960 12624 1012
rect 12676 1000 12682 1012
rect 13081 1003 13139 1009
rect 13081 1000 13093 1003
rect 12676 972 13093 1000
rect 12676 960 12682 972
rect 13081 969 13093 972
rect 13127 969 13139 1003
rect 13081 963 13139 969
rect 14182 960 14188 1012
rect 14240 960 14246 1012
rect 14458 960 14464 1012
rect 14516 960 14522 1012
rect 15010 960 15016 1012
rect 15068 1000 15074 1012
rect 15749 1003 15807 1009
rect 15749 1000 15761 1003
rect 15068 972 15761 1000
rect 15068 960 15074 972
rect 15749 969 15761 972
rect 15795 969 15807 1003
rect 15749 963 15807 969
rect 17126 960 17132 1012
rect 17184 1000 17190 1012
rect 17497 1003 17555 1009
rect 17497 1000 17509 1003
rect 17184 972 17509 1000
rect 17184 960 17190 972
rect 17497 969 17509 972
rect 17543 969 17555 1003
rect 17497 963 17555 969
rect 19978 960 19984 1012
rect 20036 1000 20042 1012
rect 20073 1003 20131 1009
rect 20073 1000 20085 1003
rect 20036 972 20085 1000
rect 20036 960 20042 972
rect 20073 969 20085 972
rect 20119 969 20131 1003
rect 20073 963 20131 969
rect 20438 960 20444 1012
rect 20496 1000 20502 1012
rect 20717 1003 20775 1009
rect 20717 1000 20729 1003
rect 20496 972 20729 1000
rect 20496 960 20502 972
rect 20717 969 20729 972
rect 20763 1000 20775 1003
rect 21818 1000 21824 1012
rect 20763 972 21824 1000
rect 20763 969 20775 972
rect 20717 963 20775 969
rect 21818 960 21824 972
rect 21876 960 21882 1012
rect 21913 1003 21971 1009
rect 21913 969 21925 1003
rect 21959 1000 21971 1003
rect 22094 1000 22100 1012
rect 21959 972 22100 1000
rect 21959 969 21971 972
rect 21913 963 21971 969
rect 22094 960 22100 972
rect 22152 960 22158 1012
rect 22462 960 22468 1012
rect 22520 1000 22526 1012
rect 22520 972 23428 1000
rect 22520 960 22526 972
rect 14200 932 14228 960
rect 14734 932 14740 944
rect 14200 904 14740 932
rect 14734 892 14740 904
rect 14792 892 14798 944
rect 12406 836 13032 864
rect 11885 799 11943 805
rect 11885 796 11897 799
rect 11716 768 11897 796
rect 11885 765 11897 768
rect 11931 765 11943 799
rect 11885 759 11943 765
rect 11977 799 12035 805
rect 11977 765 11989 799
rect 12023 796 12035 799
rect 12342 796 12348 808
rect 12023 768 12348 796
rect 12023 765 12035 768
rect 11977 759 12035 765
rect 12342 756 12348 768
rect 12400 796 12406 808
rect 12621 799 12679 805
rect 12621 796 12633 799
rect 12400 768 12633 796
rect 12400 756 12406 768
rect 12621 765 12633 768
rect 12667 765 12679 799
rect 13004 796 13032 836
rect 13170 796 13176 808
rect 13004 768 13176 796
rect 12621 759 12679 765
rect 13170 756 13176 768
rect 13228 756 13234 808
rect 13722 756 13728 808
rect 13780 796 13786 808
rect 14553 799 14611 805
rect 14553 796 14565 799
rect 13780 768 14565 796
rect 13780 756 13786 768
rect 14553 765 14565 768
rect 14599 765 14611 799
rect 14553 759 14611 765
rect 14642 756 14648 808
rect 14700 756 14706 808
rect 14752 796 14780 892
rect 18690 864 18696 876
rect 17512 836 18696 864
rect 16117 799 16175 805
rect 14752 768 15792 796
rect 12713 731 12771 737
rect 12713 697 12725 731
rect 12759 728 12771 731
rect 13740 728 13768 756
rect 12759 700 13768 728
rect 12759 697 12771 700
rect 12713 691 12771 697
rect 15654 688 15660 740
rect 15712 688 15718 740
rect 15764 728 15792 768
rect 16117 765 16129 799
rect 16163 796 16175 799
rect 16206 796 16212 808
rect 16163 768 16212 796
rect 16163 765 16175 768
rect 16117 759 16175 765
rect 16206 756 16212 768
rect 16264 796 16270 808
rect 17512 796 17540 836
rect 18690 824 18696 836
rect 18748 824 18754 876
rect 21361 867 21419 873
rect 21361 833 21373 867
rect 21407 864 21419 867
rect 21637 867 21695 873
rect 21637 864 21649 867
rect 21407 836 21649 864
rect 21407 833 21419 836
rect 21361 827 21419 833
rect 21637 833 21649 836
rect 21683 864 21695 867
rect 21683 836 21864 864
rect 21683 833 21695 836
rect 21637 827 21695 833
rect 16264 768 17540 796
rect 17589 799 17647 805
rect 16264 756 16270 768
rect 17589 765 17601 799
rect 17635 765 17647 799
rect 17589 759 17647 765
rect 16362 731 16420 737
rect 16362 728 16374 731
rect 15764 700 16374 728
rect 16362 697 16374 700
rect 16408 697 16420 731
rect 16362 691 16420 697
rect 16758 688 16764 740
rect 16816 728 16822 740
rect 17604 728 17632 759
rect 17862 756 17868 808
rect 17920 756 17926 808
rect 18960 799 19018 805
rect 18960 765 18972 799
rect 19006 796 19018 799
rect 19518 796 19524 808
rect 19006 768 19524 796
rect 19006 765 19018 768
rect 18960 759 19018 765
rect 19518 756 19524 768
rect 19576 756 19582 808
rect 20809 799 20867 805
rect 20809 765 20821 799
rect 20855 796 20867 799
rect 21266 796 21272 808
rect 20855 768 21272 796
rect 20855 765 20867 768
rect 20809 759 20867 765
rect 21266 756 21272 768
rect 21324 756 21330 808
rect 21726 756 21732 808
rect 21784 756 21790 808
rect 21836 805 21864 836
rect 21910 824 21916 876
rect 21968 864 21974 876
rect 22097 867 22155 873
rect 22097 864 22109 867
rect 21968 836 22109 864
rect 21968 824 21974 836
rect 22097 833 22109 836
rect 22143 833 22155 867
rect 22097 827 22155 833
rect 21821 799 21879 805
rect 21821 765 21833 799
rect 21867 796 21879 799
rect 22364 799 22422 805
rect 22364 796 22376 799
rect 21867 768 22376 796
rect 21867 765 21879 768
rect 21821 759 21879 765
rect 22364 765 22376 768
rect 22410 796 22422 799
rect 22922 796 22928 808
rect 22410 768 22928 796
rect 22410 765 22422 768
rect 22364 759 22422 765
rect 22922 756 22928 768
rect 22980 756 22986 808
rect 23400 796 23428 972
rect 23566 960 23572 1012
rect 23624 1000 23630 1012
rect 23937 1003 23995 1009
rect 23937 1000 23949 1003
rect 23624 972 23949 1000
rect 23624 960 23630 972
rect 23937 969 23949 972
rect 23983 969 23995 1003
rect 23937 963 23995 969
rect 23477 935 23535 941
rect 23477 901 23489 935
rect 23523 932 23535 935
rect 23842 932 23848 944
rect 23523 904 23848 932
rect 23523 901 23535 904
rect 23477 895 23535 901
rect 23842 892 23848 904
rect 23900 892 23906 944
rect 23952 864 23980 963
rect 24210 960 24216 1012
rect 24268 960 24274 1012
rect 24486 960 24492 1012
rect 24544 960 24550 1012
rect 23952 836 24164 864
rect 24136 805 24164 836
rect 24029 799 24087 805
rect 24029 796 24041 799
rect 23400 768 24041 796
rect 24029 765 24041 768
rect 24075 765 24087 799
rect 24029 759 24087 765
rect 24121 799 24179 805
rect 24121 765 24133 799
rect 24167 765 24179 799
rect 24121 759 24179 765
rect 16816 700 17632 728
rect 24044 728 24072 759
rect 24578 756 24584 808
rect 24636 756 24642 808
rect 31018 756 31024 808
rect 31076 756 31082 808
rect 24596 728 24624 756
rect 24044 700 24624 728
rect 16816 688 16822 700
rect 552 570 31531 592
rect 552 518 8102 570
rect 8154 518 8166 570
rect 8218 518 8230 570
rect 8282 518 8294 570
rect 8346 518 8358 570
rect 8410 518 15807 570
rect 15859 518 15871 570
rect 15923 518 15935 570
rect 15987 518 15999 570
rect 16051 518 16063 570
rect 16115 518 23512 570
rect 23564 518 23576 570
rect 23628 518 23640 570
rect 23692 518 23704 570
rect 23756 518 23768 570
rect 23820 518 31217 570
rect 31269 518 31281 570
rect 31333 518 31345 570
rect 31397 518 31409 570
rect 31461 518 31473 570
rect 31525 518 31531 570
rect 552 496 31531 518
rect 16114 348 16120 400
rect 16172 388 16178 400
rect 16298 388 16304 400
rect 16172 360 16304 388
rect 16172 348 16178 360
rect 16298 348 16304 360
rect 16356 348 16362 400
<< via1 >>
rect 8102 19014 8154 19066
rect 8166 19014 8218 19066
rect 8230 19014 8282 19066
rect 8294 19014 8346 19066
rect 8358 19014 8410 19066
rect 15807 19014 15859 19066
rect 15871 19014 15923 19066
rect 15935 19014 15987 19066
rect 15999 19014 16051 19066
rect 16063 19014 16115 19066
rect 23512 19014 23564 19066
rect 23576 19014 23628 19066
rect 23640 19014 23692 19066
rect 23704 19014 23756 19066
rect 23768 19014 23820 19066
rect 31217 19014 31269 19066
rect 31281 19014 31333 19066
rect 31345 19014 31397 19066
rect 31409 19014 31461 19066
rect 31473 19014 31525 19066
rect 756 18776 808 18828
rect 6460 18776 6512 18828
rect 7104 18776 7156 18828
rect 7748 18776 7800 18828
rect 1124 18751 1176 18760
rect 1124 18717 1133 18751
rect 1133 18717 1167 18751
rect 1167 18717 1176 18751
rect 1124 18708 1176 18717
rect 9496 18776 9548 18828
rect 10140 18776 10192 18828
rect 10508 18819 10560 18828
rect 10508 18785 10517 18819
rect 10517 18785 10551 18819
rect 10551 18785 10560 18819
rect 10508 18776 10560 18785
rect 10784 18776 10836 18828
rect 11428 18819 11480 18828
rect 11428 18785 11451 18819
rect 11451 18785 11480 18819
rect 11428 18776 11480 18785
rect 14188 18776 14240 18828
rect 16212 18776 16264 18828
rect 16948 18776 17000 18828
rect 20812 18819 20864 18828
rect 20812 18785 20821 18819
rect 20821 18785 20855 18819
rect 20855 18785 20864 18819
rect 20812 18776 20864 18785
rect 20996 18776 21048 18828
rect 848 18615 900 18624
rect 848 18581 857 18615
rect 857 18581 891 18615
rect 891 18581 900 18615
rect 848 18572 900 18581
rect 7932 18572 7984 18624
rect 8484 18615 8536 18624
rect 8484 18581 8493 18615
rect 8493 18581 8527 18615
rect 8527 18581 8536 18615
rect 8484 18572 8536 18581
rect 8944 18572 8996 18624
rect 9864 18572 9916 18624
rect 13636 18751 13688 18760
rect 13636 18717 13645 18751
rect 13645 18717 13679 18751
rect 13679 18717 13688 18751
rect 13636 18708 13688 18717
rect 17868 18708 17920 18760
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 15016 18615 15068 18624
rect 15016 18581 15025 18615
rect 15025 18581 15059 18615
rect 15059 18581 15068 18615
rect 15016 18572 15068 18581
rect 17040 18572 17092 18624
rect 19984 18572 20036 18624
rect 20720 18572 20772 18624
rect 23204 18776 23256 18828
rect 27712 18776 27764 18828
rect 28356 18776 28408 18828
rect 31668 18776 31720 18828
rect 25228 18751 25280 18760
rect 25228 18717 25237 18751
rect 25237 18717 25271 18751
rect 25271 18717 25280 18751
rect 25228 18708 25280 18717
rect 22284 18572 22336 18624
rect 22744 18615 22796 18624
rect 22744 18581 22753 18615
rect 22753 18581 22787 18615
rect 22787 18581 22796 18615
rect 22744 18572 22796 18581
rect 23020 18572 23072 18624
rect 24032 18572 24084 18624
rect 31024 18615 31076 18624
rect 31024 18581 31033 18615
rect 31033 18581 31067 18615
rect 31067 18581 31076 18615
rect 31024 18572 31076 18581
rect 4250 18470 4302 18522
rect 4314 18470 4366 18522
rect 4378 18470 4430 18522
rect 4442 18470 4494 18522
rect 4506 18470 4558 18522
rect 11955 18470 12007 18522
rect 12019 18470 12071 18522
rect 12083 18470 12135 18522
rect 12147 18470 12199 18522
rect 12211 18470 12263 18522
rect 19660 18470 19712 18522
rect 19724 18470 19776 18522
rect 19788 18470 19840 18522
rect 19852 18470 19904 18522
rect 19916 18470 19968 18522
rect 27365 18470 27417 18522
rect 27429 18470 27481 18522
rect 27493 18470 27545 18522
rect 27557 18470 27609 18522
rect 27621 18470 27673 18522
rect 9496 18411 9548 18420
rect 9496 18377 9505 18411
rect 9505 18377 9539 18411
rect 9539 18377 9548 18411
rect 9496 18368 9548 18377
rect 8576 18300 8628 18352
rect 7380 18232 7432 18284
rect 7748 18232 7800 18284
rect 848 18207 900 18216
rect 848 18173 857 18207
rect 857 18173 891 18207
rect 891 18173 900 18207
rect 848 18164 900 18173
rect 7104 18028 7156 18080
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 8484 18164 8536 18216
rect 8944 18207 8996 18216
rect 8944 18173 8953 18207
rect 8953 18173 8987 18207
rect 8987 18173 8996 18207
rect 8944 18164 8996 18173
rect 10140 18368 10192 18420
rect 10600 18368 10652 18420
rect 11428 18300 11480 18352
rect 9772 18232 9824 18284
rect 9864 18207 9916 18216
rect 9864 18173 9873 18207
rect 9873 18173 9907 18207
rect 9907 18173 9916 18207
rect 9864 18164 9916 18173
rect 14188 18411 14240 18420
rect 14188 18377 14197 18411
rect 14197 18377 14231 18411
rect 14231 18377 14240 18411
rect 14188 18368 14240 18377
rect 20812 18368 20864 18420
rect 20996 18411 21048 18420
rect 20996 18377 21005 18411
rect 21005 18377 21039 18411
rect 21039 18377 21048 18411
rect 20996 18368 21048 18377
rect 22744 18411 22796 18420
rect 22744 18377 22753 18411
rect 22753 18377 22787 18411
rect 22787 18377 22796 18411
rect 22744 18368 22796 18377
rect 23020 18411 23072 18420
rect 23020 18377 23029 18411
rect 23029 18377 23063 18411
rect 23063 18377 23072 18411
rect 23020 18368 23072 18377
rect 10324 18096 10376 18148
rect 12256 18207 12308 18216
rect 12256 18173 12265 18207
rect 12265 18173 12299 18207
rect 12299 18173 12308 18207
rect 12256 18164 12308 18173
rect 7932 18028 7984 18080
rect 9220 18071 9272 18080
rect 9220 18037 9229 18071
rect 9229 18037 9263 18071
rect 9263 18037 9272 18071
rect 9220 18028 9272 18037
rect 11612 18028 11664 18080
rect 14004 18300 14056 18352
rect 12992 18207 13044 18216
rect 12992 18173 13001 18207
rect 13001 18173 13035 18207
rect 13035 18173 13044 18207
rect 12992 18164 13044 18173
rect 13728 18207 13780 18216
rect 13728 18173 13737 18207
rect 13737 18173 13771 18207
rect 13771 18173 13780 18207
rect 13728 18164 13780 18173
rect 16212 18164 16264 18216
rect 16948 18164 17000 18216
rect 19984 18232 20036 18284
rect 13360 18028 13412 18080
rect 18696 18096 18748 18148
rect 16304 18028 16356 18080
rect 16580 18028 16632 18080
rect 16948 18071 17000 18080
rect 16948 18037 16957 18071
rect 16957 18037 16991 18071
rect 16991 18037 17000 18071
rect 16948 18028 17000 18037
rect 18788 18028 18840 18080
rect 19248 18071 19300 18080
rect 19248 18037 19257 18071
rect 19257 18037 19291 18071
rect 19291 18037 19300 18071
rect 19248 18028 19300 18037
rect 22836 18207 22888 18216
rect 22836 18173 22845 18207
rect 22845 18173 22879 18207
rect 22879 18173 22888 18207
rect 22836 18164 22888 18173
rect 23204 18164 23256 18216
rect 22284 18139 22336 18148
rect 22284 18105 22293 18139
rect 22293 18105 22327 18139
rect 22327 18105 22336 18139
rect 22284 18096 22336 18105
rect 24308 18164 24360 18216
rect 24952 18207 25004 18216
rect 24952 18173 24961 18207
rect 24961 18173 24995 18207
rect 24995 18173 25004 18207
rect 24952 18164 25004 18173
rect 22376 18028 22428 18080
rect 8102 17926 8154 17978
rect 8166 17926 8218 17978
rect 8230 17926 8282 17978
rect 8294 17926 8346 17978
rect 8358 17926 8410 17978
rect 15807 17926 15859 17978
rect 15871 17926 15923 17978
rect 15935 17926 15987 17978
rect 15999 17926 16051 17978
rect 16063 17926 16115 17978
rect 23512 17926 23564 17978
rect 23576 17926 23628 17978
rect 23640 17926 23692 17978
rect 23704 17926 23756 17978
rect 23768 17926 23820 17978
rect 31217 17926 31269 17978
rect 31281 17926 31333 17978
rect 31345 17926 31397 17978
rect 31409 17926 31461 17978
rect 31473 17926 31525 17978
rect 7104 17824 7156 17876
rect 12256 17867 12308 17876
rect 12256 17833 12265 17867
rect 12265 17833 12299 17867
rect 12299 17833 12308 17867
rect 12256 17824 12308 17833
rect 8576 17799 8628 17808
rect 8576 17765 8588 17799
rect 8588 17765 8628 17799
rect 8576 17756 8628 17765
rect 7748 17731 7800 17740
rect 7748 17697 7757 17731
rect 7757 17697 7791 17731
rect 7791 17697 7800 17731
rect 7748 17688 7800 17697
rect 7932 17688 7984 17740
rect 8024 17620 8076 17672
rect 12348 17731 12400 17740
rect 12348 17697 12357 17731
rect 12357 17697 12391 17731
rect 12391 17697 12400 17731
rect 12348 17688 12400 17697
rect 12992 17824 13044 17876
rect 13360 17867 13412 17876
rect 13360 17833 13369 17867
rect 13369 17833 13403 17867
rect 13403 17833 13412 17867
rect 13360 17824 13412 17833
rect 13728 17824 13780 17876
rect 12900 17731 12952 17740
rect 12900 17697 12909 17731
rect 12909 17697 12943 17731
rect 12943 17697 12952 17731
rect 12900 17688 12952 17697
rect 12992 17688 13044 17740
rect 13636 17731 13688 17740
rect 13636 17697 13645 17731
rect 13645 17697 13679 17731
rect 13679 17697 13688 17731
rect 13636 17688 13688 17697
rect 16488 17756 16540 17808
rect 16212 17688 16264 17740
rect 18696 17756 18748 17808
rect 24308 17867 24360 17876
rect 24308 17833 24317 17867
rect 24317 17833 24351 17867
rect 24351 17833 24360 17867
rect 24308 17824 24360 17833
rect 24952 17824 25004 17876
rect 16948 17688 17000 17740
rect 19248 17756 19300 17808
rect 22376 17799 22428 17808
rect 22376 17765 22394 17799
rect 22394 17765 22428 17799
rect 22376 17756 22428 17765
rect 22836 17756 22888 17808
rect 21916 17688 21968 17740
rect 24308 17688 24360 17740
rect 25320 17731 25372 17740
rect 25320 17697 25329 17731
rect 25329 17697 25363 17731
rect 25363 17697 25372 17731
rect 25320 17688 25372 17697
rect 25596 17731 25648 17740
rect 25596 17697 25605 17731
rect 25605 17697 25639 17731
rect 25639 17697 25648 17731
rect 25596 17688 25648 17697
rect 26148 17731 26200 17740
rect 26148 17697 26157 17731
rect 26157 17697 26191 17731
rect 26191 17697 26200 17731
rect 26148 17688 26200 17697
rect 6460 17527 6512 17536
rect 6460 17493 6469 17527
rect 6469 17493 6503 17527
rect 6503 17493 6512 17527
rect 6460 17484 6512 17493
rect 7012 17527 7064 17536
rect 7012 17493 7021 17527
rect 7021 17493 7055 17527
rect 7055 17493 7064 17527
rect 7012 17484 7064 17493
rect 7932 17527 7984 17536
rect 7932 17493 7941 17527
rect 7941 17493 7975 17527
rect 7975 17493 7984 17527
rect 7932 17484 7984 17493
rect 14648 17484 14700 17536
rect 15660 17484 15712 17536
rect 17776 17527 17828 17536
rect 17776 17493 17785 17527
rect 17785 17493 17819 17527
rect 17819 17493 17828 17527
rect 17776 17484 17828 17493
rect 19248 17527 19300 17536
rect 19248 17493 19257 17527
rect 19257 17493 19291 17527
rect 19291 17493 19300 17527
rect 19248 17484 19300 17493
rect 19524 17527 19576 17536
rect 19524 17493 19533 17527
rect 19533 17493 19567 17527
rect 19567 17493 19576 17527
rect 19524 17484 19576 17493
rect 19984 17484 20036 17536
rect 21272 17527 21324 17536
rect 21272 17493 21281 17527
rect 21281 17493 21315 17527
rect 21315 17493 21324 17527
rect 21272 17484 21324 17493
rect 23204 17484 23256 17536
rect 23848 17484 23900 17536
rect 25228 17620 25280 17672
rect 4250 17382 4302 17434
rect 4314 17382 4366 17434
rect 4378 17382 4430 17434
rect 4442 17382 4494 17434
rect 4506 17382 4558 17434
rect 11955 17382 12007 17434
rect 12019 17382 12071 17434
rect 12083 17382 12135 17434
rect 12147 17382 12199 17434
rect 12211 17382 12263 17434
rect 19660 17382 19712 17434
rect 19724 17382 19776 17434
rect 19788 17382 19840 17434
rect 19852 17382 19904 17434
rect 19916 17382 19968 17434
rect 27365 17382 27417 17434
rect 27429 17382 27481 17434
rect 27493 17382 27545 17434
rect 27557 17382 27609 17434
rect 27621 17382 27673 17434
rect 6460 17280 6512 17332
rect 7012 17280 7064 17332
rect 6000 17212 6052 17264
rect 848 17119 900 17128
rect 848 17085 857 17119
rect 857 17085 891 17119
rect 891 17085 900 17119
rect 848 17076 900 17085
rect 5632 17144 5684 17196
rect 7380 17119 7432 17128
rect 7380 17085 7389 17119
rect 7389 17085 7423 17119
rect 7423 17085 7432 17119
rect 7380 17076 7432 17085
rect 7932 17076 7984 17128
rect 9772 17076 9824 17128
rect 10784 17076 10836 17128
rect 9220 17008 9272 17060
rect 12348 17280 12400 17332
rect 19524 17280 19576 17332
rect 12808 17212 12860 17264
rect 16856 17212 16908 17264
rect 11888 17119 11940 17128
rect 11888 17085 11897 17119
rect 11897 17085 11931 17119
rect 11931 17085 11940 17119
rect 11888 17076 11940 17085
rect 12164 17119 12216 17128
rect 12164 17085 12173 17119
rect 12173 17085 12207 17119
rect 12207 17085 12216 17119
rect 12164 17076 12216 17085
rect 12440 17076 12492 17128
rect 13636 17144 13688 17196
rect 17868 17187 17920 17196
rect 17868 17153 17877 17187
rect 17877 17153 17911 17187
rect 17911 17153 17920 17187
rect 20444 17212 20496 17264
rect 17868 17144 17920 17153
rect 19524 17144 19576 17196
rect 19984 17076 20036 17128
rect 21916 17280 21968 17332
rect 25320 17323 25372 17332
rect 25320 17289 25329 17323
rect 25329 17289 25363 17323
rect 25363 17289 25372 17323
rect 25320 17280 25372 17289
rect 25320 17144 25372 17196
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 5724 16983 5776 16992
rect 5724 16949 5733 16983
rect 5733 16949 5767 16983
rect 5767 16949 5776 16983
rect 5724 16940 5776 16949
rect 8484 16940 8536 16992
rect 11704 16940 11756 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 17408 16940 17460 16992
rect 19248 16940 19300 16992
rect 24308 17008 24360 17060
rect 25412 17119 25464 17128
rect 25412 17085 25421 17119
rect 25421 17085 25455 17119
rect 25455 17085 25464 17119
rect 25412 17076 25464 17085
rect 25688 17119 25740 17128
rect 25688 17085 25697 17119
rect 25697 17085 25731 17119
rect 25731 17085 25740 17119
rect 25688 17076 25740 17085
rect 27068 17076 27120 17128
rect 26148 17051 26200 17060
rect 26148 17017 26157 17051
rect 26157 17017 26191 17051
rect 26191 17017 26200 17051
rect 27436 17051 27488 17060
rect 26148 17008 26200 17017
rect 27436 17017 27454 17051
rect 27454 17017 27488 17051
rect 27436 17008 27488 17017
rect 21088 16983 21140 16992
rect 21088 16949 21097 16983
rect 21097 16949 21131 16983
rect 21131 16949 21140 16983
rect 21088 16940 21140 16949
rect 21548 16983 21600 16992
rect 21548 16949 21557 16983
rect 21557 16949 21591 16983
rect 21591 16949 21600 16983
rect 21548 16940 21600 16949
rect 23112 16983 23164 16992
rect 23112 16949 23121 16983
rect 23121 16949 23155 16983
rect 23155 16949 23164 16983
rect 23112 16940 23164 16949
rect 25596 16983 25648 16992
rect 25596 16949 25605 16983
rect 25605 16949 25639 16983
rect 25639 16949 25648 16983
rect 25596 16940 25648 16949
rect 26332 16983 26384 16992
rect 26332 16949 26341 16983
rect 26341 16949 26375 16983
rect 26375 16949 26384 16983
rect 26332 16940 26384 16949
rect 30012 16940 30064 16992
rect 8102 16838 8154 16890
rect 8166 16838 8218 16890
rect 8230 16838 8282 16890
rect 8294 16838 8346 16890
rect 8358 16838 8410 16890
rect 15807 16838 15859 16890
rect 15871 16838 15923 16890
rect 15935 16838 15987 16890
rect 15999 16838 16051 16890
rect 16063 16838 16115 16890
rect 23512 16838 23564 16890
rect 23576 16838 23628 16890
rect 23640 16838 23692 16890
rect 23704 16838 23756 16890
rect 23768 16838 23820 16890
rect 31217 16838 31269 16890
rect 31281 16838 31333 16890
rect 31345 16838 31397 16890
rect 31409 16838 31461 16890
rect 31473 16838 31525 16890
rect 5448 16736 5500 16788
rect 2412 16600 2464 16652
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 5724 16600 5776 16652
rect 6552 16736 6604 16788
rect 8024 16736 8076 16788
rect 11888 16736 11940 16788
rect 12440 16779 12492 16788
rect 12440 16745 12449 16779
rect 12449 16745 12483 16779
rect 12483 16745 12492 16779
rect 12440 16736 12492 16745
rect 12900 16736 12952 16788
rect 6460 16668 6512 16720
rect 8392 16668 8444 16720
rect 8116 16600 8168 16652
rect 10140 16643 10192 16652
rect 10140 16609 10149 16643
rect 10149 16609 10183 16643
rect 10183 16609 10192 16643
rect 10140 16600 10192 16609
rect 11428 16600 11480 16652
rect 13636 16668 13688 16720
rect 19248 16668 19300 16720
rect 1952 16439 2004 16448
rect 1952 16405 1961 16439
rect 1961 16405 1995 16439
rect 1995 16405 2004 16439
rect 1952 16396 2004 16405
rect 3516 16396 3568 16448
rect 4160 16439 4212 16448
rect 4160 16405 4169 16439
rect 4169 16405 4203 16439
rect 4203 16405 4212 16439
rect 4160 16396 4212 16405
rect 11796 16600 11848 16652
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 12624 16532 12676 16584
rect 17868 16600 17920 16652
rect 21088 16736 21140 16788
rect 25688 16779 25740 16788
rect 25688 16745 25697 16779
rect 25697 16745 25731 16779
rect 25731 16745 25740 16779
rect 25688 16736 25740 16745
rect 27160 16779 27212 16788
rect 20444 16668 20496 16720
rect 20720 16643 20772 16652
rect 20720 16609 20729 16643
rect 20729 16609 20763 16643
rect 20763 16609 20772 16643
rect 20720 16600 20772 16609
rect 21548 16600 21600 16652
rect 22376 16600 22428 16652
rect 23664 16600 23716 16652
rect 24308 16600 24360 16652
rect 25412 16600 25464 16652
rect 27160 16745 27169 16779
rect 27169 16745 27203 16779
rect 27203 16745 27212 16779
rect 27160 16736 27212 16745
rect 11796 16464 11848 16516
rect 6552 16396 6604 16448
rect 7748 16439 7800 16448
rect 7748 16405 7757 16439
rect 7757 16405 7791 16439
rect 7791 16405 7800 16439
rect 7748 16396 7800 16405
rect 9404 16439 9456 16448
rect 9404 16405 9413 16439
rect 9413 16405 9447 16439
rect 9447 16405 9456 16439
rect 9404 16396 9456 16405
rect 10232 16439 10284 16448
rect 10232 16405 10241 16439
rect 10241 16405 10275 16439
rect 10275 16405 10284 16439
rect 10232 16396 10284 16405
rect 11060 16396 11112 16448
rect 11428 16439 11480 16448
rect 11428 16405 11437 16439
rect 11437 16405 11471 16439
rect 11471 16405 11480 16439
rect 11428 16396 11480 16405
rect 14556 16439 14608 16448
rect 14556 16405 14565 16439
rect 14565 16405 14599 16439
rect 14599 16405 14608 16439
rect 14556 16396 14608 16405
rect 18144 16396 18196 16448
rect 19432 16464 19484 16516
rect 19156 16439 19208 16448
rect 19156 16405 19165 16439
rect 19165 16405 19199 16439
rect 19199 16405 19208 16439
rect 19156 16396 19208 16405
rect 19984 16464 20036 16516
rect 26424 16532 26476 16584
rect 21456 16396 21508 16448
rect 27436 16643 27488 16652
rect 27436 16609 27445 16643
rect 27445 16609 27479 16643
rect 27479 16609 27488 16643
rect 27436 16600 27488 16609
rect 28724 16600 28776 16652
rect 29184 16600 29236 16652
rect 27160 16532 27212 16584
rect 30012 16575 30064 16584
rect 30012 16541 30021 16575
rect 30021 16541 30055 16575
rect 30055 16541 30064 16575
rect 30012 16532 30064 16541
rect 22008 16396 22060 16448
rect 24952 16439 25004 16448
rect 24952 16405 24961 16439
rect 24961 16405 24995 16439
rect 24995 16405 25004 16439
rect 24952 16396 25004 16405
rect 26884 16439 26936 16448
rect 26884 16405 26893 16439
rect 26893 16405 26927 16439
rect 26927 16405 26936 16439
rect 26884 16396 26936 16405
rect 28264 16396 28316 16448
rect 4250 16294 4302 16346
rect 4314 16294 4366 16346
rect 4378 16294 4430 16346
rect 4442 16294 4494 16346
rect 4506 16294 4558 16346
rect 11955 16294 12007 16346
rect 12019 16294 12071 16346
rect 12083 16294 12135 16346
rect 12147 16294 12199 16346
rect 12211 16294 12263 16346
rect 19660 16294 19712 16346
rect 19724 16294 19776 16346
rect 19788 16294 19840 16346
rect 19852 16294 19904 16346
rect 19916 16294 19968 16346
rect 27365 16294 27417 16346
rect 27429 16294 27481 16346
rect 27493 16294 27545 16346
rect 27557 16294 27609 16346
rect 27621 16294 27673 16346
rect 1952 16192 2004 16244
rect 11060 16235 11112 16244
rect 11060 16201 11069 16235
rect 11069 16201 11103 16235
rect 11103 16201 11112 16235
rect 11060 16192 11112 16201
rect 11428 16235 11480 16244
rect 11428 16201 11437 16235
rect 11437 16201 11471 16235
rect 11471 16201 11480 16235
rect 11428 16192 11480 16201
rect 11612 16192 11664 16244
rect 14832 16192 14884 16244
rect 2412 16167 2464 16176
rect 2412 16133 2421 16167
rect 2421 16133 2455 16167
rect 2455 16133 2464 16167
rect 2412 16124 2464 16133
rect 3240 15988 3292 16040
rect 1492 15852 1544 15904
rect 2412 15852 2464 15904
rect 2688 15895 2740 15904
rect 2688 15861 2697 15895
rect 2697 15861 2731 15895
rect 2731 15861 2740 15895
rect 2688 15852 2740 15861
rect 10876 16124 10928 16176
rect 8392 16099 8444 16108
rect 8392 16065 8401 16099
rect 8401 16065 8435 16099
rect 8435 16065 8444 16099
rect 8392 16056 8444 16065
rect 3516 16031 3568 16040
rect 3516 15997 3525 16031
rect 3525 15997 3559 16031
rect 3559 15997 3568 16031
rect 3516 15988 3568 15997
rect 5632 15988 5684 16040
rect 6460 15988 6512 16040
rect 8484 15988 8536 16040
rect 10140 16056 10192 16108
rect 10232 16056 10284 16108
rect 10692 15988 10744 16040
rect 17868 16056 17920 16108
rect 20536 16192 20588 16244
rect 19984 16124 20036 16176
rect 20720 16124 20772 16176
rect 11888 15988 11940 16040
rect 12624 15988 12676 16040
rect 18144 15988 18196 16040
rect 12348 15920 12400 15972
rect 15476 15920 15528 15972
rect 4160 15852 4212 15904
rect 6368 15895 6420 15904
rect 6368 15861 6377 15895
rect 6377 15861 6411 15895
rect 6411 15861 6420 15895
rect 6368 15852 6420 15861
rect 11796 15852 11848 15904
rect 13452 15852 13504 15904
rect 16028 15895 16080 15904
rect 16028 15861 16037 15895
rect 16037 15861 16071 15895
rect 16071 15861 16080 15895
rect 16028 15852 16080 15861
rect 16488 15852 16540 15904
rect 18328 15852 18380 15904
rect 18512 15852 18564 15904
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 19432 16031 19484 16040
rect 19432 15997 19449 16031
rect 19449 15997 19483 16031
rect 19483 15997 19484 16031
rect 19432 15988 19484 15997
rect 20536 15988 20588 16040
rect 26884 16235 26936 16244
rect 26884 16201 26893 16235
rect 26893 16201 26927 16235
rect 26927 16201 26936 16235
rect 26884 16192 26936 16201
rect 28724 16235 28776 16244
rect 28724 16201 28733 16235
rect 28733 16201 28767 16235
rect 28767 16201 28776 16235
rect 28724 16192 28776 16201
rect 23940 16124 23992 16176
rect 29184 16192 29236 16244
rect 22008 16056 22060 16108
rect 21456 15988 21508 16040
rect 21916 15988 21968 16040
rect 22376 16031 22428 16040
rect 22376 15997 22410 16031
rect 22410 15997 22428 16031
rect 22376 15988 22428 15997
rect 23664 15988 23716 16040
rect 27068 16056 27120 16108
rect 27528 16031 27580 16040
rect 27528 15997 27537 16031
rect 27537 15997 27571 16031
rect 27571 15997 27580 16031
rect 27528 15988 27580 15997
rect 20996 15920 21048 15972
rect 19248 15852 19300 15904
rect 19984 15852 20036 15904
rect 25412 15920 25464 15972
rect 26424 15963 26476 15972
rect 26424 15929 26442 15963
rect 26442 15929 26476 15963
rect 26424 15920 26476 15929
rect 23848 15895 23900 15904
rect 23848 15861 23857 15895
rect 23857 15861 23891 15895
rect 23891 15861 23900 15895
rect 23848 15852 23900 15861
rect 24768 15852 24820 15904
rect 29000 15920 29052 15972
rect 28448 15895 28500 15904
rect 28448 15861 28457 15895
rect 28457 15861 28491 15895
rect 28491 15861 28500 15895
rect 28448 15852 28500 15861
rect 28632 15852 28684 15904
rect 29276 15852 29328 15904
rect 8102 15750 8154 15802
rect 8166 15750 8218 15802
rect 8230 15750 8282 15802
rect 8294 15750 8346 15802
rect 8358 15750 8410 15802
rect 15807 15750 15859 15802
rect 15871 15750 15923 15802
rect 15935 15750 15987 15802
rect 15999 15750 16051 15802
rect 16063 15750 16115 15802
rect 23512 15750 23564 15802
rect 23576 15750 23628 15802
rect 23640 15750 23692 15802
rect 23704 15750 23756 15802
rect 23768 15750 23820 15802
rect 31217 15750 31269 15802
rect 31281 15750 31333 15802
rect 31345 15750 31397 15802
rect 31409 15750 31461 15802
rect 31473 15750 31525 15802
rect 1952 15648 2004 15700
rect 2688 15648 2740 15700
rect 10140 15648 10192 15700
rect 10232 15648 10284 15700
rect 1492 15512 1544 15564
rect 6552 15580 6604 15632
rect 2136 15376 2188 15428
rect 4252 15512 4304 15564
rect 6460 15555 6512 15564
rect 6460 15521 6469 15555
rect 6469 15521 6503 15555
rect 6503 15521 6512 15555
rect 6460 15512 6512 15521
rect 2688 15487 2740 15496
rect 2688 15453 2697 15487
rect 2697 15453 2731 15487
rect 2731 15453 2740 15487
rect 2688 15444 2740 15453
rect 9496 15512 9548 15564
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 10140 15555 10192 15564
rect 10140 15521 10149 15555
rect 10149 15521 10183 15555
rect 10183 15521 10192 15555
rect 10140 15512 10192 15521
rect 1768 15351 1820 15360
rect 1768 15317 1777 15351
rect 1777 15317 1811 15351
rect 1811 15317 1820 15351
rect 1768 15308 1820 15317
rect 2320 15351 2372 15360
rect 2320 15317 2329 15351
rect 2329 15317 2363 15351
rect 2363 15317 2372 15351
rect 2320 15308 2372 15317
rect 4068 15351 4120 15360
rect 4068 15317 4077 15351
rect 4077 15317 4111 15351
rect 4111 15317 4120 15351
rect 4068 15308 4120 15317
rect 5816 15308 5868 15360
rect 7380 15308 7432 15360
rect 11796 15648 11848 15700
rect 10784 15580 10836 15632
rect 10692 15512 10744 15564
rect 11244 15512 11296 15564
rect 11888 15580 11940 15632
rect 12624 15648 12676 15700
rect 15476 15648 15528 15700
rect 19064 15691 19116 15700
rect 19064 15657 19073 15691
rect 19073 15657 19107 15691
rect 19107 15657 19116 15691
rect 19064 15648 19116 15657
rect 19248 15648 19300 15700
rect 18512 15623 18564 15632
rect 18512 15589 18521 15623
rect 18521 15589 18555 15623
rect 18555 15589 18564 15623
rect 18512 15580 18564 15589
rect 15844 15444 15896 15496
rect 18328 15555 18380 15564
rect 18328 15521 18337 15555
rect 18337 15521 18371 15555
rect 18371 15521 18380 15555
rect 18328 15512 18380 15521
rect 19984 15648 20036 15700
rect 20996 15648 21048 15700
rect 23848 15648 23900 15700
rect 22008 15580 22060 15632
rect 19340 15487 19392 15496
rect 19340 15453 19349 15487
rect 19349 15453 19383 15487
rect 19383 15453 19392 15487
rect 19340 15444 19392 15453
rect 10692 15376 10744 15428
rect 14924 15376 14976 15428
rect 12900 15351 12952 15360
rect 12900 15317 12909 15351
rect 12909 15317 12943 15351
rect 12943 15317 12952 15351
rect 12900 15308 12952 15317
rect 15108 15308 15160 15360
rect 15568 15376 15620 15428
rect 15384 15308 15436 15360
rect 15476 15351 15528 15360
rect 15476 15317 15485 15351
rect 15485 15317 15519 15351
rect 15519 15317 15528 15351
rect 15476 15308 15528 15317
rect 16764 15351 16816 15360
rect 16764 15317 16773 15351
rect 16773 15317 16807 15351
rect 16807 15317 16816 15351
rect 16764 15308 16816 15317
rect 21916 15555 21968 15564
rect 21916 15521 21925 15555
rect 21925 15521 21959 15555
rect 21959 15521 21968 15555
rect 21916 15512 21968 15521
rect 24308 15555 24360 15564
rect 24308 15521 24312 15555
rect 24312 15521 24346 15555
rect 24346 15521 24360 15555
rect 24308 15512 24360 15521
rect 24400 15555 24452 15564
rect 24400 15521 24409 15555
rect 24409 15521 24443 15555
rect 24443 15521 24452 15555
rect 24400 15512 24452 15521
rect 27528 15623 27580 15632
rect 27528 15589 27546 15623
rect 27546 15589 27580 15623
rect 28448 15691 28500 15700
rect 28448 15657 28457 15691
rect 28457 15657 28491 15691
rect 28491 15657 28500 15691
rect 28448 15648 28500 15657
rect 29000 15648 29052 15700
rect 30012 15648 30064 15700
rect 27528 15580 27580 15589
rect 24216 15444 24268 15496
rect 25964 15512 26016 15564
rect 27068 15512 27120 15564
rect 28632 15512 28684 15564
rect 19064 15308 19116 15360
rect 20720 15351 20772 15360
rect 20720 15317 20729 15351
rect 20729 15317 20763 15351
rect 20763 15317 20772 15351
rect 20720 15308 20772 15317
rect 20904 15351 20956 15360
rect 20904 15317 20913 15351
rect 20913 15317 20947 15351
rect 20947 15317 20956 15351
rect 20904 15308 20956 15317
rect 20996 15308 21048 15360
rect 23940 15308 23992 15360
rect 24124 15351 24176 15360
rect 24124 15317 24133 15351
rect 24133 15317 24167 15351
rect 24167 15317 24176 15351
rect 24124 15308 24176 15317
rect 26240 15308 26292 15360
rect 28816 15376 28868 15428
rect 29184 15376 29236 15428
rect 29552 15555 29604 15564
rect 29552 15521 29561 15555
rect 29561 15521 29595 15555
rect 29595 15521 29604 15555
rect 29552 15512 29604 15521
rect 30932 15351 30984 15360
rect 30932 15317 30941 15351
rect 30941 15317 30975 15351
rect 30975 15317 30984 15351
rect 30932 15308 30984 15317
rect 4250 15206 4302 15258
rect 4314 15206 4366 15258
rect 4378 15206 4430 15258
rect 4442 15206 4494 15258
rect 4506 15206 4558 15258
rect 11955 15206 12007 15258
rect 12019 15206 12071 15258
rect 12083 15206 12135 15258
rect 12147 15206 12199 15258
rect 12211 15206 12263 15258
rect 19660 15206 19712 15258
rect 19724 15206 19776 15258
rect 19788 15206 19840 15258
rect 19852 15206 19904 15258
rect 19916 15206 19968 15258
rect 27365 15206 27417 15258
rect 27429 15206 27481 15258
rect 27493 15206 27545 15258
rect 27557 15206 27609 15258
rect 27621 15206 27673 15258
rect 1768 15104 1820 15156
rect 9496 15104 9548 15156
rect 8208 15079 8260 15088
rect 8208 15045 8217 15079
rect 8217 15045 8251 15079
rect 8251 15045 8260 15079
rect 8208 15036 8260 15045
rect 13728 15104 13780 15156
rect 2688 14968 2740 15020
rect 2136 14943 2188 14952
rect 2136 14909 2145 14943
rect 2145 14909 2179 14943
rect 2179 14909 2188 14943
rect 2136 14900 2188 14909
rect 2320 14900 2372 14952
rect 6460 14968 6512 15020
rect 13084 14968 13136 15020
rect 15384 15104 15436 15156
rect 18788 15104 18840 15156
rect 20996 15104 21048 15156
rect 24400 15104 24452 15156
rect 28724 15147 28776 15156
rect 28724 15113 28733 15147
rect 28733 15113 28767 15147
rect 28767 15113 28776 15147
rect 28724 15104 28776 15113
rect 15292 15079 15344 15088
rect 15292 15045 15301 15079
rect 15301 15045 15335 15079
rect 15335 15045 15344 15079
rect 15292 15036 15344 15045
rect 4712 14832 4764 14884
rect 6092 14832 6144 14884
rect 9956 14900 10008 14952
rect 10784 14900 10836 14952
rect 11060 14900 11112 14952
rect 11888 14900 11940 14952
rect 15476 14968 15528 15020
rect 10140 14832 10192 14884
rect 10508 14832 10560 14884
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 6000 14807 6052 14816
rect 6000 14773 6009 14807
rect 6009 14773 6043 14807
rect 6043 14773 6052 14807
rect 6000 14764 6052 14773
rect 9680 14764 9732 14816
rect 13636 14764 13688 14816
rect 14188 14807 14240 14816
rect 14188 14773 14197 14807
rect 14197 14773 14231 14807
rect 14231 14773 14240 14807
rect 14188 14764 14240 14773
rect 14464 14807 14516 14816
rect 14464 14773 14473 14807
rect 14473 14773 14507 14807
rect 14507 14773 14516 14807
rect 14464 14764 14516 14773
rect 14924 14900 14976 14952
rect 16212 15011 16264 15020
rect 16212 14977 16221 15011
rect 16221 14977 16255 15011
rect 16255 14977 16264 15011
rect 16212 14968 16264 14977
rect 15568 14832 15620 14884
rect 15844 14943 15896 14952
rect 15844 14909 15853 14943
rect 15853 14909 15887 14943
rect 15887 14909 15896 14943
rect 15844 14900 15896 14909
rect 16764 14900 16816 14952
rect 17684 14943 17736 14952
rect 17684 14909 17693 14943
rect 17693 14909 17727 14943
rect 17727 14909 17736 14943
rect 17684 14900 17736 14909
rect 17868 14943 17920 14952
rect 17868 14909 17877 14943
rect 17877 14909 17911 14943
rect 17911 14909 17920 14943
rect 17868 14900 17920 14909
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 19064 15036 19116 15088
rect 19800 15036 19852 15088
rect 22744 15036 22796 15088
rect 29276 15104 29328 15156
rect 20536 14968 20588 15020
rect 23296 14968 23348 15020
rect 19064 14943 19116 14952
rect 19064 14909 19073 14943
rect 19073 14909 19107 14943
rect 19107 14909 19116 14943
rect 19064 14900 19116 14909
rect 19340 14900 19392 14952
rect 20996 14943 21048 14952
rect 20996 14909 21030 14943
rect 21030 14909 21048 14943
rect 20996 14900 21048 14909
rect 18236 14807 18288 14816
rect 18236 14773 18245 14807
rect 18245 14773 18279 14807
rect 18279 14773 18288 14807
rect 18236 14764 18288 14773
rect 21180 14832 21232 14884
rect 21364 14764 21416 14816
rect 22100 14807 22152 14816
rect 22100 14773 22109 14807
rect 22109 14773 22143 14807
rect 22143 14773 22152 14807
rect 22100 14764 22152 14773
rect 23940 14943 23992 14952
rect 23940 14909 23950 14943
rect 23950 14909 23984 14943
rect 23984 14909 23992 14943
rect 23940 14900 23992 14909
rect 24308 14900 24360 14952
rect 24584 14900 24636 14952
rect 25964 14900 26016 14952
rect 28724 14968 28776 15020
rect 29644 15036 29696 15088
rect 26240 14832 26292 14884
rect 26792 14832 26844 14884
rect 29184 14943 29236 14952
rect 29184 14909 29193 14943
rect 29193 14909 29227 14943
rect 29227 14909 29236 14943
rect 29184 14900 29236 14909
rect 29460 14943 29512 14952
rect 29460 14909 29469 14943
rect 29469 14909 29503 14943
rect 29503 14909 29512 14943
rect 29460 14900 29512 14909
rect 24308 14764 24360 14816
rect 29368 14807 29420 14816
rect 29368 14773 29377 14807
rect 29377 14773 29411 14807
rect 29411 14773 29420 14807
rect 29368 14764 29420 14773
rect 29644 14807 29696 14816
rect 29644 14773 29653 14807
rect 29653 14773 29687 14807
rect 29687 14773 29696 14807
rect 29644 14764 29696 14773
rect 8102 14662 8154 14714
rect 8166 14662 8218 14714
rect 8230 14662 8282 14714
rect 8294 14662 8346 14714
rect 8358 14662 8410 14714
rect 15807 14662 15859 14714
rect 15871 14662 15923 14714
rect 15935 14662 15987 14714
rect 15999 14662 16051 14714
rect 16063 14662 16115 14714
rect 23512 14662 23564 14714
rect 23576 14662 23628 14714
rect 23640 14662 23692 14714
rect 23704 14662 23756 14714
rect 23768 14662 23820 14714
rect 31217 14662 31269 14714
rect 31281 14662 31333 14714
rect 31345 14662 31397 14714
rect 31409 14662 31461 14714
rect 31473 14662 31525 14714
rect 1768 14560 1820 14612
rect 2228 14560 2280 14612
rect 5356 14560 5408 14612
rect 2320 14492 2372 14544
rect 4712 14492 4764 14544
rect 9680 14560 9732 14612
rect 10508 14603 10560 14612
rect 10508 14569 10517 14603
rect 10517 14569 10551 14603
rect 10551 14569 10560 14603
rect 10508 14560 10560 14569
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 1400 14288 1452 14340
rect 2688 14356 2740 14408
rect 5908 14467 5960 14476
rect 5908 14433 5917 14467
rect 5917 14433 5951 14467
rect 5951 14433 5960 14467
rect 5908 14424 5960 14433
rect 6460 14424 6512 14476
rect 6276 14356 6328 14408
rect 9772 14424 9824 14476
rect 9864 14356 9916 14408
rect 11060 14424 11112 14476
rect 11244 14467 11296 14476
rect 11244 14433 11278 14467
rect 11278 14433 11296 14467
rect 11244 14424 11296 14433
rect 13084 14467 13136 14476
rect 13084 14433 13093 14467
rect 13093 14433 13127 14467
rect 13127 14433 13136 14467
rect 13084 14424 13136 14433
rect 14188 14560 14240 14612
rect 18236 14560 18288 14612
rect 20444 14560 20496 14612
rect 14004 14492 14056 14544
rect 15016 14492 15068 14544
rect 12440 14356 12492 14408
rect 13360 14356 13412 14408
rect 14464 14424 14516 14476
rect 15200 14467 15252 14476
rect 15200 14433 15209 14467
rect 15209 14433 15243 14467
rect 15243 14433 15252 14467
rect 15200 14424 15252 14433
rect 16212 14424 16264 14476
rect 19340 14492 19392 14544
rect 19800 14467 19852 14476
rect 19800 14433 19823 14467
rect 19823 14433 19852 14467
rect 19800 14424 19852 14433
rect 17868 14356 17920 14408
rect 19064 14356 19116 14408
rect 21916 14560 21968 14612
rect 21640 14424 21692 14476
rect 22560 14424 22612 14476
rect 22928 14424 22980 14476
rect 23204 14535 23256 14544
rect 23204 14501 23213 14535
rect 23213 14501 23247 14535
rect 23247 14501 23256 14535
rect 23204 14492 23256 14501
rect 23664 14535 23716 14544
rect 23664 14501 23673 14535
rect 23673 14501 23707 14535
rect 23707 14501 23716 14535
rect 23664 14492 23716 14501
rect 26792 14603 26844 14612
rect 26792 14569 26801 14603
rect 26801 14569 26835 14603
rect 26835 14569 26844 14603
rect 26792 14560 26844 14569
rect 24952 14492 25004 14544
rect 29184 14560 29236 14612
rect 23940 14467 23992 14476
rect 23940 14433 23949 14467
rect 23949 14433 23983 14467
rect 23983 14433 23992 14467
rect 23940 14424 23992 14433
rect 24032 14467 24084 14476
rect 24032 14433 24042 14467
rect 24042 14433 24076 14467
rect 24076 14433 24084 14467
rect 24032 14424 24084 14433
rect 24216 14467 24268 14476
rect 24216 14433 24225 14467
rect 24225 14433 24259 14467
rect 24259 14433 24268 14467
rect 24216 14424 24268 14433
rect 4896 14220 4948 14272
rect 4988 14263 5040 14272
rect 4988 14229 4997 14263
rect 4997 14229 5031 14263
rect 5031 14229 5040 14263
rect 4988 14220 5040 14229
rect 6092 14220 6144 14272
rect 10140 14220 10192 14272
rect 11704 14220 11756 14272
rect 12348 14263 12400 14272
rect 12348 14229 12357 14263
rect 12357 14229 12391 14263
rect 12391 14229 12400 14263
rect 12348 14220 12400 14229
rect 13268 14220 13320 14272
rect 15476 14288 15528 14340
rect 14188 14220 14240 14272
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 15292 14220 15344 14272
rect 19432 14288 19484 14340
rect 17960 14263 18012 14272
rect 17960 14229 17969 14263
rect 17969 14229 18003 14263
rect 18003 14229 18012 14263
rect 17960 14220 18012 14229
rect 18880 14220 18932 14272
rect 21088 14220 21140 14272
rect 22284 14220 22336 14272
rect 22652 14263 22704 14272
rect 22652 14229 22661 14263
rect 22661 14229 22695 14263
rect 22695 14229 22704 14263
rect 22652 14220 22704 14229
rect 22836 14263 22888 14272
rect 22836 14229 22845 14263
rect 22845 14229 22879 14263
rect 22879 14229 22888 14263
rect 22836 14220 22888 14229
rect 23480 14356 23532 14408
rect 24584 14424 24636 14476
rect 26792 14424 26844 14476
rect 26608 14356 26660 14408
rect 27804 14424 27856 14476
rect 27712 14356 27764 14408
rect 28908 14492 28960 14544
rect 29552 14492 29604 14544
rect 29644 14492 29696 14544
rect 28080 14288 28132 14340
rect 23296 14263 23348 14272
rect 23296 14229 23305 14263
rect 23305 14229 23339 14263
rect 23339 14229 23348 14263
rect 23296 14220 23348 14229
rect 23940 14220 23992 14272
rect 24032 14220 24084 14272
rect 24676 14263 24728 14272
rect 24676 14229 24685 14263
rect 24685 14229 24719 14263
rect 24719 14229 24728 14263
rect 24676 14220 24728 14229
rect 24860 14263 24912 14272
rect 24860 14229 24869 14263
rect 24869 14229 24903 14263
rect 24903 14229 24912 14263
rect 24860 14220 24912 14229
rect 29276 14288 29328 14340
rect 29460 14220 29512 14272
rect 4250 14118 4302 14170
rect 4314 14118 4366 14170
rect 4378 14118 4430 14170
rect 4442 14118 4494 14170
rect 4506 14118 4558 14170
rect 11955 14118 12007 14170
rect 12019 14118 12071 14170
rect 12083 14118 12135 14170
rect 12147 14118 12199 14170
rect 12211 14118 12263 14170
rect 19660 14118 19712 14170
rect 19724 14118 19776 14170
rect 19788 14118 19840 14170
rect 19852 14118 19904 14170
rect 19916 14118 19968 14170
rect 27365 14118 27417 14170
rect 27429 14118 27481 14170
rect 27493 14118 27545 14170
rect 27557 14118 27609 14170
rect 27621 14118 27673 14170
rect 1584 14016 1636 14068
rect 1216 13923 1268 13932
rect 1216 13889 1225 13923
rect 1225 13889 1259 13923
rect 1259 13889 1268 13923
rect 2688 14016 2740 14068
rect 4988 14016 5040 14068
rect 5908 14016 5960 14068
rect 6920 14016 6972 14068
rect 7840 14016 7892 14068
rect 3976 13948 4028 14000
rect 1216 13880 1268 13889
rect 2228 13812 2280 13864
rect 4160 13744 4212 13796
rect 4896 13855 4948 13864
rect 4896 13821 4905 13855
rect 4905 13821 4939 13855
rect 4939 13821 4948 13855
rect 6092 13948 6144 14000
rect 4896 13812 4948 13821
rect 5448 13812 5500 13864
rect 6276 13880 6328 13932
rect 7564 13880 7616 13932
rect 5172 13676 5224 13728
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 7656 13855 7708 13864
rect 7656 13821 7665 13855
rect 7665 13821 7699 13855
rect 7699 13821 7708 13855
rect 7656 13812 7708 13821
rect 8024 13880 8076 13932
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 7840 13857 7892 13864
rect 7840 13823 7849 13857
rect 7849 13823 7883 13857
rect 7883 13823 7892 13857
rect 7840 13812 7892 13823
rect 8484 13744 8536 13796
rect 7472 13676 7524 13728
rect 11704 13812 11756 13864
rect 10140 13787 10192 13796
rect 10140 13753 10174 13787
rect 10174 13753 10192 13787
rect 10140 13744 10192 13753
rect 10784 13744 10836 13796
rect 10048 13676 10100 13728
rect 11244 13719 11296 13728
rect 11244 13685 11253 13719
rect 11253 13685 11287 13719
rect 11287 13685 11296 13719
rect 11244 13676 11296 13685
rect 11520 13719 11572 13728
rect 11520 13685 11529 13719
rect 11529 13685 11563 13719
rect 11563 13685 11572 13719
rect 11520 13676 11572 13685
rect 13268 14016 13320 14068
rect 13820 14059 13872 14068
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 15476 14016 15528 14068
rect 15200 13948 15252 14000
rect 17500 14016 17552 14068
rect 19984 14016 20036 14068
rect 20076 14016 20128 14068
rect 20996 14016 21048 14068
rect 21180 14016 21232 14068
rect 12440 13880 12492 13932
rect 14096 13880 14148 13932
rect 14280 13880 14332 13932
rect 14740 13880 14792 13932
rect 14832 13923 14884 13932
rect 14832 13889 14841 13923
rect 14841 13889 14875 13923
rect 14875 13889 14884 13923
rect 14832 13880 14884 13889
rect 14924 13880 14976 13932
rect 15292 13880 15344 13932
rect 18512 13948 18564 14000
rect 21732 14016 21784 14068
rect 22284 14016 22336 14068
rect 22652 14016 22704 14068
rect 22836 14016 22888 14068
rect 23296 14016 23348 14068
rect 23480 14016 23532 14068
rect 24860 14016 24912 14068
rect 26792 14059 26844 14068
rect 26792 14025 26801 14059
rect 26801 14025 26835 14059
rect 26835 14025 26844 14059
rect 26792 14016 26844 14025
rect 27712 14016 27764 14068
rect 29368 14059 29420 14068
rect 29368 14025 29377 14059
rect 29377 14025 29411 14059
rect 29411 14025 29420 14059
rect 29368 14016 29420 14025
rect 30932 14016 30984 14068
rect 22376 13948 22428 14000
rect 12164 13744 12216 13796
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 14004 13812 14056 13864
rect 13636 13787 13688 13796
rect 13636 13753 13645 13787
rect 13645 13753 13679 13787
rect 13679 13753 13688 13787
rect 13636 13744 13688 13753
rect 13728 13744 13780 13796
rect 15108 13787 15160 13796
rect 15108 13753 15126 13787
rect 15126 13753 15160 13787
rect 12808 13676 12860 13728
rect 13084 13719 13136 13728
rect 13084 13685 13093 13719
rect 13093 13685 13127 13719
rect 13127 13685 13136 13719
rect 13084 13676 13136 13685
rect 13176 13676 13228 13728
rect 14004 13719 14056 13728
rect 14004 13685 14013 13719
rect 14013 13685 14047 13719
rect 14047 13685 14056 13719
rect 14004 13676 14056 13685
rect 14832 13676 14884 13728
rect 15108 13744 15160 13753
rect 15200 13787 15252 13796
rect 15200 13753 15209 13787
rect 15209 13753 15243 13787
rect 15243 13753 15252 13787
rect 15200 13744 15252 13753
rect 15384 13744 15436 13796
rect 15568 13787 15620 13796
rect 15568 13753 15577 13787
rect 15577 13753 15611 13787
rect 15611 13753 15620 13787
rect 15568 13744 15620 13753
rect 16120 13812 16172 13864
rect 15936 13744 15988 13796
rect 16764 13812 16816 13864
rect 17776 13812 17828 13864
rect 16672 13744 16724 13796
rect 18052 13744 18104 13796
rect 18696 13787 18748 13796
rect 18696 13753 18705 13787
rect 18705 13753 18739 13787
rect 18739 13753 18748 13787
rect 18696 13744 18748 13753
rect 20444 13812 20496 13864
rect 19800 13744 19852 13796
rect 20352 13787 20404 13796
rect 20352 13753 20361 13787
rect 20361 13753 20395 13787
rect 20395 13753 20404 13787
rect 20352 13744 20404 13753
rect 20904 13812 20956 13864
rect 20996 13855 21048 13864
rect 20996 13821 21005 13855
rect 21005 13821 21039 13855
rect 21039 13821 21048 13855
rect 20996 13812 21048 13821
rect 21088 13855 21140 13864
rect 21088 13821 21097 13855
rect 21097 13821 21131 13855
rect 21131 13821 21140 13855
rect 21088 13812 21140 13821
rect 21364 13812 21416 13864
rect 21456 13855 21508 13864
rect 21456 13821 21465 13855
rect 21465 13821 21499 13855
rect 21499 13821 21508 13855
rect 21456 13812 21508 13821
rect 21548 13812 21600 13864
rect 20812 13787 20864 13796
rect 20812 13753 20821 13787
rect 20821 13753 20855 13787
rect 20855 13753 20864 13787
rect 20812 13744 20864 13753
rect 16396 13719 16448 13728
rect 16396 13685 16426 13719
rect 16426 13685 16448 13719
rect 16396 13676 16448 13685
rect 16948 13676 17000 13728
rect 17132 13719 17184 13728
rect 17132 13685 17141 13719
rect 17141 13685 17175 13719
rect 17175 13685 17184 13719
rect 17132 13676 17184 13685
rect 17316 13719 17368 13728
rect 17316 13685 17343 13719
rect 17343 13685 17368 13719
rect 17316 13676 17368 13685
rect 17592 13676 17644 13728
rect 18788 13676 18840 13728
rect 18880 13719 18932 13728
rect 18880 13685 18905 13719
rect 18905 13685 18932 13719
rect 18880 13676 18932 13685
rect 19248 13676 19300 13728
rect 19340 13676 19392 13728
rect 20168 13719 20220 13728
rect 20168 13685 20195 13719
rect 20195 13685 20220 13719
rect 20168 13676 20220 13685
rect 21180 13676 21232 13728
rect 21732 13855 21784 13864
rect 21732 13821 21741 13855
rect 21741 13821 21775 13855
rect 21775 13821 21784 13855
rect 21732 13812 21784 13821
rect 22468 13812 22520 13864
rect 23020 13812 23072 13864
rect 23572 13812 23624 13864
rect 22008 13744 22060 13796
rect 22560 13744 22612 13796
rect 23848 13787 23900 13796
rect 23848 13753 23857 13787
rect 23857 13753 23891 13787
rect 23891 13753 23900 13787
rect 23848 13744 23900 13753
rect 26608 13880 26660 13932
rect 28080 13948 28132 14000
rect 25964 13855 26016 13864
rect 25964 13821 25973 13855
rect 25973 13821 26007 13855
rect 26007 13821 26016 13855
rect 25964 13812 26016 13821
rect 22284 13719 22336 13728
rect 22284 13685 22293 13719
rect 22293 13685 22327 13719
rect 22327 13685 22336 13719
rect 22284 13676 22336 13685
rect 22376 13676 22428 13728
rect 23204 13676 23256 13728
rect 23388 13719 23440 13728
rect 23388 13685 23397 13719
rect 23397 13685 23431 13719
rect 23431 13685 23440 13719
rect 23388 13676 23440 13685
rect 24216 13719 24268 13728
rect 24216 13685 24225 13719
rect 24225 13685 24259 13719
rect 24259 13685 24268 13719
rect 24216 13676 24268 13685
rect 25044 13676 25096 13728
rect 26516 13812 26568 13864
rect 27804 13880 27856 13932
rect 29184 13880 29236 13932
rect 26792 13744 26844 13796
rect 26608 13676 26660 13728
rect 29276 13812 29328 13864
rect 28080 13744 28132 13796
rect 29460 13676 29512 13728
rect 8102 13574 8154 13626
rect 8166 13574 8218 13626
rect 8230 13574 8282 13626
rect 8294 13574 8346 13626
rect 8358 13574 8410 13626
rect 15807 13574 15859 13626
rect 15871 13574 15923 13626
rect 15935 13574 15987 13626
rect 15999 13574 16051 13626
rect 16063 13574 16115 13626
rect 23512 13574 23564 13626
rect 23576 13574 23628 13626
rect 23640 13574 23692 13626
rect 23704 13574 23756 13626
rect 23768 13574 23820 13626
rect 31217 13574 31269 13626
rect 31281 13574 31333 13626
rect 31345 13574 31397 13626
rect 31409 13574 31461 13626
rect 31473 13574 31525 13626
rect 1216 13472 1268 13524
rect 4160 13472 4212 13524
rect 4712 13472 4764 13524
rect 5172 13515 5224 13524
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 8024 13472 8076 13524
rect 9864 13515 9916 13524
rect 9864 13481 9873 13515
rect 9873 13481 9907 13515
rect 9907 13481 9916 13515
rect 9864 13472 9916 13481
rect 10140 13515 10192 13524
rect 10140 13481 10149 13515
rect 10149 13481 10183 13515
rect 10183 13481 10192 13515
rect 10140 13472 10192 13481
rect 11612 13472 11664 13524
rect 1400 13404 1452 13456
rect 1768 13336 1820 13388
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 4804 13379 4856 13388
rect 4804 13345 4813 13379
rect 4813 13345 4847 13379
rect 4847 13345 4856 13379
rect 4804 13336 4856 13345
rect 4988 13336 5040 13388
rect 3056 13243 3108 13252
rect 3056 13209 3065 13243
rect 3065 13209 3099 13243
rect 3099 13209 3108 13243
rect 3056 13200 3108 13209
rect 5448 13268 5500 13320
rect 7564 13336 7616 13388
rect 8484 13379 8536 13388
rect 8484 13345 8493 13379
rect 8493 13345 8527 13379
rect 8527 13345 8536 13379
rect 8484 13336 8536 13345
rect 12348 13472 12400 13524
rect 16580 13472 16632 13524
rect 16764 13515 16816 13524
rect 16764 13481 16773 13515
rect 16773 13481 16807 13515
rect 16807 13481 16816 13515
rect 16764 13472 16816 13481
rect 16856 13472 16908 13524
rect 12992 13404 13044 13456
rect 12164 13379 12216 13388
rect 7656 13268 7708 13320
rect 9312 13268 9364 13320
rect 9772 13268 9824 13320
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 13636 13404 13688 13456
rect 13728 13336 13780 13388
rect 7288 13200 7340 13252
rect 12072 13268 12124 13320
rect 12808 13200 12860 13252
rect 13084 13200 13136 13252
rect 14096 13200 14148 13252
rect 1124 13132 1176 13184
rect 4160 13132 4212 13184
rect 7564 13132 7616 13184
rect 9312 13132 9364 13184
rect 11612 13132 11664 13184
rect 11796 13132 11848 13184
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 14372 13336 14424 13388
rect 14832 13336 14884 13388
rect 15384 13404 15436 13456
rect 15752 13336 15804 13388
rect 16856 13336 16908 13388
rect 17132 13336 17184 13388
rect 17776 13404 17828 13456
rect 22836 13472 22888 13524
rect 23388 13472 23440 13524
rect 18328 13404 18380 13456
rect 18880 13404 18932 13456
rect 19156 13447 19208 13456
rect 19156 13413 19165 13447
rect 19165 13413 19199 13447
rect 19199 13413 19208 13447
rect 19156 13404 19208 13413
rect 18052 13379 18104 13388
rect 18052 13345 18066 13379
rect 18066 13345 18100 13379
rect 18100 13345 18104 13379
rect 18052 13336 18104 13345
rect 18604 13336 18656 13388
rect 14832 13175 14884 13184
rect 14832 13141 14841 13175
rect 14841 13141 14875 13175
rect 14875 13141 14884 13175
rect 14832 13132 14884 13141
rect 15200 13132 15252 13184
rect 15476 13132 15528 13184
rect 16396 13132 16448 13184
rect 16856 13132 16908 13184
rect 17224 13132 17276 13184
rect 17592 13132 17644 13184
rect 18052 13132 18104 13184
rect 18236 13175 18288 13184
rect 18236 13141 18245 13175
rect 18245 13141 18279 13175
rect 18279 13141 18288 13175
rect 18236 13132 18288 13141
rect 19340 13336 19392 13388
rect 19432 13379 19484 13388
rect 19432 13345 19441 13379
rect 19441 13345 19475 13379
rect 19475 13345 19484 13379
rect 19432 13336 19484 13345
rect 20168 13336 20220 13388
rect 20076 13268 20128 13320
rect 21640 13404 21692 13456
rect 20536 13379 20588 13388
rect 20536 13345 20545 13379
rect 20545 13345 20579 13379
rect 20579 13345 20588 13379
rect 20536 13336 20588 13345
rect 21180 13336 21232 13388
rect 21548 13336 21600 13388
rect 21824 13336 21876 13388
rect 22192 13336 22244 13388
rect 24400 13336 24452 13388
rect 25044 13336 25096 13388
rect 19156 13200 19208 13252
rect 20536 13200 20588 13252
rect 21364 13268 21416 13320
rect 21732 13268 21784 13320
rect 23480 13268 23532 13320
rect 24584 13268 24636 13320
rect 26608 13472 26660 13524
rect 26792 13515 26844 13524
rect 26792 13481 26801 13515
rect 26801 13481 26835 13515
rect 26835 13481 26844 13515
rect 26792 13472 26844 13481
rect 27712 13472 27764 13524
rect 28080 13447 28132 13456
rect 28080 13413 28098 13447
rect 28098 13413 28132 13447
rect 28080 13404 28132 13413
rect 29276 13404 29328 13456
rect 26516 13336 26568 13388
rect 25412 13268 25464 13320
rect 25688 13268 25740 13320
rect 25964 13268 26016 13320
rect 23296 13200 23348 13252
rect 19064 13132 19116 13184
rect 19432 13132 19484 13184
rect 20444 13132 20496 13184
rect 21640 13175 21692 13184
rect 21640 13141 21649 13175
rect 21649 13141 21683 13175
rect 21683 13141 21692 13175
rect 21640 13132 21692 13141
rect 25044 13132 25096 13184
rect 29092 13132 29144 13184
rect 4250 13030 4302 13082
rect 4314 13030 4366 13082
rect 4378 13030 4430 13082
rect 4442 13030 4494 13082
rect 4506 13030 4558 13082
rect 11955 13030 12007 13082
rect 12019 13030 12071 13082
rect 12083 13030 12135 13082
rect 12147 13030 12199 13082
rect 12211 13030 12263 13082
rect 19660 13030 19712 13082
rect 19724 13030 19776 13082
rect 19788 13030 19840 13082
rect 19852 13030 19904 13082
rect 19916 13030 19968 13082
rect 27365 13030 27417 13082
rect 27429 13030 27481 13082
rect 27493 13030 27545 13082
rect 27557 13030 27609 13082
rect 27621 13030 27673 13082
rect 4160 12928 4212 12980
rect 7288 12928 7340 12980
rect 7472 12928 7524 12980
rect 9312 12971 9364 12980
rect 9312 12937 9321 12971
rect 9321 12937 9355 12971
rect 9355 12937 9364 12971
rect 9312 12928 9364 12937
rect 1308 12767 1360 12776
rect 1308 12733 1317 12767
rect 1317 12733 1351 12767
rect 1351 12733 1360 12767
rect 1308 12724 1360 12733
rect 1400 12724 1452 12776
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 4160 12724 4212 12776
rect 4804 12792 4856 12844
rect 1124 12588 1176 12640
rect 3056 12631 3108 12640
rect 3056 12597 3065 12631
rect 3065 12597 3099 12631
rect 3099 12597 3108 12631
rect 3056 12588 3108 12597
rect 4252 12588 4304 12640
rect 6092 12767 6144 12776
rect 6092 12733 6101 12767
rect 6101 12733 6135 12767
rect 6135 12733 6144 12767
rect 6092 12724 6144 12733
rect 7932 12792 7984 12844
rect 10048 12928 10100 12980
rect 11796 12928 11848 12980
rect 13176 12971 13228 12980
rect 13176 12937 13185 12971
rect 13185 12937 13219 12971
rect 13219 12937 13228 12971
rect 13176 12928 13228 12937
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 14188 12928 14240 12980
rect 16488 12928 16540 12980
rect 16672 12971 16724 12980
rect 7656 12724 7708 12776
rect 10968 12792 11020 12844
rect 14648 12860 14700 12912
rect 14924 12860 14976 12912
rect 16212 12860 16264 12912
rect 16672 12937 16703 12971
rect 16703 12937 16724 12971
rect 16672 12928 16724 12937
rect 17684 12928 17736 12980
rect 19064 12928 19116 12980
rect 17500 12860 17552 12912
rect 17776 12860 17828 12912
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 9680 12767 9732 12776
rect 9680 12733 9689 12767
rect 9689 12733 9723 12767
rect 9723 12733 9732 12767
rect 9680 12724 9732 12733
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 13912 12767 13964 12776
rect 13912 12733 13921 12767
rect 13921 12733 13955 12767
rect 13955 12733 13964 12767
rect 13912 12724 13964 12733
rect 14188 12724 14240 12776
rect 15476 12724 15528 12776
rect 15752 12724 15804 12776
rect 7104 12656 7156 12708
rect 7196 12699 7248 12708
rect 7196 12665 7205 12699
rect 7205 12665 7239 12699
rect 7239 12665 7248 12699
rect 7196 12656 7248 12665
rect 9864 12656 9916 12708
rect 4988 12588 5040 12640
rect 7472 12588 7524 12640
rect 8024 12631 8076 12640
rect 8024 12597 8033 12631
rect 8033 12597 8067 12631
rect 8067 12597 8076 12631
rect 8024 12588 8076 12597
rect 11980 12631 12032 12640
rect 11980 12597 12015 12631
rect 12015 12597 12032 12631
rect 11980 12588 12032 12597
rect 12164 12631 12216 12640
rect 12164 12597 12173 12631
rect 12173 12597 12207 12631
rect 12207 12597 12216 12631
rect 12164 12588 12216 12597
rect 12256 12588 12308 12640
rect 13084 12588 13136 12640
rect 14740 12656 14792 12708
rect 17408 12792 17460 12844
rect 17040 12724 17092 12776
rect 13452 12588 13504 12640
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 17408 12588 17460 12640
rect 17776 12767 17828 12776
rect 17776 12733 17785 12767
rect 17785 12733 17819 12767
rect 17819 12733 17828 12767
rect 17776 12724 17828 12733
rect 17868 12767 17920 12776
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 17868 12724 17920 12733
rect 18604 12792 18656 12844
rect 19156 12792 19208 12844
rect 21824 12928 21876 12980
rect 18144 12767 18196 12776
rect 18144 12733 18153 12767
rect 18153 12733 18187 12767
rect 18187 12733 18196 12767
rect 18144 12724 18196 12733
rect 19248 12767 19300 12776
rect 19248 12733 19257 12767
rect 19257 12733 19291 12767
rect 19291 12733 19300 12767
rect 19248 12724 19300 12733
rect 19432 12767 19484 12776
rect 19432 12733 19441 12767
rect 19441 12733 19475 12767
rect 19475 12733 19484 12767
rect 19432 12724 19484 12733
rect 18788 12699 18840 12708
rect 18788 12665 18797 12699
rect 18797 12665 18831 12699
rect 18831 12665 18840 12699
rect 18788 12656 18840 12665
rect 20076 12724 20128 12776
rect 20168 12767 20220 12776
rect 20168 12733 20177 12767
rect 20177 12733 20211 12767
rect 20211 12733 20220 12767
rect 20168 12724 20220 12733
rect 20628 12792 20680 12844
rect 20260 12656 20312 12708
rect 20904 12767 20956 12776
rect 20904 12733 20913 12767
rect 20913 12733 20947 12767
rect 20947 12733 20956 12767
rect 20904 12724 20956 12733
rect 23388 12928 23440 12980
rect 24952 12928 25004 12980
rect 25044 12971 25096 12980
rect 25044 12937 25053 12971
rect 25053 12937 25087 12971
rect 25087 12937 25096 12971
rect 25044 12928 25096 12937
rect 30748 12971 30800 12980
rect 30748 12937 30757 12971
rect 30757 12937 30791 12971
rect 30791 12937 30800 12971
rect 30748 12928 30800 12937
rect 25688 12792 25740 12844
rect 29184 12792 29236 12844
rect 22560 12724 22612 12776
rect 23388 12724 23440 12776
rect 23848 12724 23900 12776
rect 24400 12767 24452 12776
rect 24400 12733 24409 12767
rect 24409 12733 24443 12767
rect 24443 12733 24452 12767
rect 24400 12724 24452 12733
rect 22744 12656 22796 12708
rect 25044 12724 25096 12776
rect 29000 12767 29052 12776
rect 29000 12733 29009 12767
rect 29009 12733 29043 12767
rect 29043 12733 29052 12767
rect 29000 12724 29052 12733
rect 29092 12724 29144 12776
rect 29460 12724 29512 12776
rect 26424 12699 26476 12708
rect 26424 12665 26442 12699
rect 26442 12665 26476 12699
rect 26424 12656 26476 12665
rect 18972 12588 19024 12640
rect 19248 12588 19300 12640
rect 20628 12588 20680 12640
rect 22836 12588 22888 12640
rect 23020 12588 23072 12640
rect 23388 12588 23440 12640
rect 25320 12631 25372 12640
rect 25320 12597 25329 12631
rect 25329 12597 25363 12631
rect 25363 12597 25372 12631
rect 25320 12588 25372 12597
rect 25412 12588 25464 12640
rect 26976 12656 27028 12708
rect 29276 12588 29328 12640
rect 29920 12588 29972 12640
rect 8102 12486 8154 12538
rect 8166 12486 8218 12538
rect 8230 12486 8282 12538
rect 8294 12486 8346 12538
rect 8358 12486 8410 12538
rect 15807 12486 15859 12538
rect 15871 12486 15923 12538
rect 15935 12486 15987 12538
rect 15999 12486 16051 12538
rect 16063 12486 16115 12538
rect 23512 12486 23564 12538
rect 23576 12486 23628 12538
rect 23640 12486 23692 12538
rect 23704 12486 23756 12538
rect 23768 12486 23820 12538
rect 31217 12486 31269 12538
rect 31281 12486 31333 12538
rect 31345 12486 31397 12538
rect 31409 12486 31461 12538
rect 31473 12486 31525 12538
rect 1400 12384 1452 12436
rect 4252 12384 4304 12436
rect 1584 12316 1636 12368
rect 3700 12248 3752 12300
rect 4528 12291 4580 12300
rect 4528 12257 4562 12291
rect 4562 12257 4580 12291
rect 4528 12248 4580 12257
rect 6552 12359 6604 12368
rect 6552 12325 6561 12359
rect 6561 12325 6595 12359
rect 6595 12325 6604 12359
rect 6552 12316 6604 12325
rect 6828 12427 6880 12436
rect 6828 12393 6837 12427
rect 6837 12393 6871 12427
rect 6871 12393 6880 12427
rect 6828 12384 6880 12393
rect 7104 12384 7156 12436
rect 8024 12384 8076 12436
rect 9680 12384 9732 12436
rect 6920 12316 6972 12368
rect 1308 12112 1360 12164
rect 6828 12248 6880 12300
rect 7472 12316 7524 12368
rect 7748 12316 7800 12368
rect 10048 12316 10100 12368
rect 9128 12248 9180 12300
rect 9588 12291 9640 12300
rect 9588 12257 9597 12291
rect 9597 12257 9631 12291
rect 9631 12257 9640 12291
rect 9588 12248 9640 12257
rect 9772 12248 9824 12300
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 11520 12384 11572 12436
rect 11888 12384 11940 12436
rect 12256 12427 12308 12436
rect 12256 12393 12265 12427
rect 12265 12393 12299 12427
rect 12299 12393 12308 12427
rect 12256 12384 12308 12393
rect 12624 12384 12676 12436
rect 15384 12384 15436 12436
rect 15476 12384 15528 12436
rect 12072 12316 12124 12368
rect 11888 12291 11940 12300
rect 11888 12257 11897 12291
rect 11897 12257 11931 12291
rect 11931 12257 11940 12291
rect 11888 12248 11940 12257
rect 12992 12359 13044 12368
rect 12992 12325 13001 12359
rect 13001 12325 13035 12359
rect 13035 12325 13044 12359
rect 12992 12316 13044 12325
rect 13084 12316 13136 12368
rect 13728 12316 13780 12368
rect 17040 12316 17092 12368
rect 17684 12384 17736 12436
rect 17776 12359 17828 12368
rect 17776 12325 17785 12359
rect 17785 12325 17819 12359
rect 17819 12325 17828 12359
rect 17776 12316 17828 12325
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 4160 12044 4212 12096
rect 7012 12180 7064 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 10968 12180 11020 12232
rect 7196 12112 7248 12164
rect 11612 12112 11664 12164
rect 15200 12248 15252 12300
rect 15292 12291 15344 12300
rect 15292 12257 15301 12291
rect 15301 12257 15335 12291
rect 15335 12257 15344 12291
rect 15292 12248 15344 12257
rect 13820 12180 13872 12232
rect 14924 12180 14976 12232
rect 15568 12291 15620 12300
rect 15568 12257 15577 12291
rect 15577 12257 15611 12291
rect 15611 12257 15620 12291
rect 15568 12248 15620 12257
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 15752 12248 15804 12300
rect 16396 12248 16448 12300
rect 16580 12248 16632 12300
rect 16764 12248 16816 12300
rect 16856 12248 16908 12300
rect 16488 12180 16540 12232
rect 17040 12180 17092 12232
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 8024 12044 8076 12096
rect 15200 12112 15252 12164
rect 15936 12155 15988 12164
rect 15936 12121 15945 12155
rect 15945 12121 15979 12155
rect 15979 12121 15988 12155
rect 15936 12112 15988 12121
rect 16028 12112 16080 12164
rect 17684 12291 17736 12300
rect 17684 12257 17693 12291
rect 17693 12257 17727 12291
rect 17727 12257 17736 12291
rect 17684 12248 17736 12257
rect 18144 12384 18196 12436
rect 18512 12384 18564 12436
rect 18788 12384 18840 12436
rect 19340 12384 19392 12436
rect 19524 12384 19576 12436
rect 21640 12384 21692 12436
rect 18236 12316 18288 12368
rect 19064 12316 19116 12368
rect 19248 12316 19300 12368
rect 19340 12291 19392 12300
rect 19340 12257 19349 12291
rect 19349 12257 19383 12291
rect 19383 12257 19392 12291
rect 19340 12248 19392 12257
rect 18144 12180 18196 12232
rect 19616 12291 19668 12300
rect 19616 12257 19625 12291
rect 19625 12257 19659 12291
rect 19659 12257 19668 12291
rect 19616 12248 19668 12257
rect 17868 12112 17920 12164
rect 18604 12112 18656 12164
rect 19892 12112 19944 12164
rect 20536 12316 20588 12368
rect 21456 12316 21508 12368
rect 23020 12359 23072 12368
rect 23020 12325 23029 12359
rect 23029 12325 23063 12359
rect 23063 12325 23072 12359
rect 23020 12316 23072 12325
rect 23112 12359 23164 12368
rect 23112 12325 23121 12359
rect 23121 12325 23155 12359
rect 23155 12325 23164 12359
rect 23112 12316 23164 12325
rect 23480 12384 23532 12436
rect 24400 12384 24452 12436
rect 24860 12384 24912 12436
rect 28632 12384 28684 12436
rect 20904 12180 20956 12232
rect 20076 12112 20128 12164
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 16580 12087 16632 12096
rect 16580 12053 16589 12087
rect 16589 12053 16623 12087
rect 16623 12053 16632 12087
rect 16580 12044 16632 12053
rect 16856 12087 16908 12096
rect 16856 12053 16865 12087
rect 16865 12053 16899 12087
rect 16899 12053 16908 12087
rect 16856 12044 16908 12053
rect 16948 12044 17000 12096
rect 18236 12044 18288 12096
rect 22376 12044 22428 12096
rect 22744 12291 22796 12300
rect 22744 12257 22753 12291
rect 22753 12257 22787 12291
rect 22787 12257 22796 12291
rect 22744 12248 22796 12257
rect 22836 12291 22888 12300
rect 22836 12257 22846 12291
rect 22846 12257 22880 12291
rect 22880 12257 22888 12291
rect 22836 12248 22888 12257
rect 23204 12291 23256 12300
rect 23204 12257 23218 12291
rect 23218 12257 23252 12291
rect 23252 12257 23256 12291
rect 23204 12248 23256 12257
rect 24032 12291 24084 12300
rect 24032 12257 24041 12291
rect 24041 12257 24075 12291
rect 24075 12257 24084 12291
rect 24032 12248 24084 12257
rect 26976 12316 27028 12368
rect 24676 12291 24728 12300
rect 24676 12257 24685 12291
rect 24685 12257 24719 12291
rect 24719 12257 24728 12291
rect 24676 12248 24728 12257
rect 22652 12112 22704 12164
rect 22836 12112 22888 12164
rect 23572 12112 23624 12164
rect 28172 12248 28224 12300
rect 29092 12316 29144 12368
rect 29276 12248 29328 12300
rect 29828 12291 29880 12300
rect 29828 12257 29837 12291
rect 29837 12257 29871 12291
rect 29871 12257 29880 12291
rect 29828 12248 29880 12257
rect 29920 12291 29972 12300
rect 29920 12257 29929 12291
rect 29929 12257 29963 12291
rect 29963 12257 29972 12291
rect 29920 12248 29972 12257
rect 30380 12044 30432 12096
rect 4250 11942 4302 11994
rect 4314 11942 4366 11994
rect 4378 11942 4430 11994
rect 4442 11942 4494 11994
rect 4506 11942 4558 11994
rect 11955 11942 12007 11994
rect 12019 11942 12071 11994
rect 12083 11942 12135 11994
rect 12147 11942 12199 11994
rect 12211 11942 12263 11994
rect 19660 11942 19712 11994
rect 19724 11942 19776 11994
rect 19788 11942 19840 11994
rect 19852 11942 19904 11994
rect 19916 11942 19968 11994
rect 27365 11942 27417 11994
rect 27429 11942 27481 11994
rect 27493 11942 27545 11994
rect 27557 11942 27609 11994
rect 27621 11942 27673 11994
rect 1400 11840 1452 11892
rect 1492 11840 1544 11892
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 1584 11636 1636 11688
rect 3332 11704 3384 11756
rect 4160 11840 4212 11892
rect 5264 11840 5316 11892
rect 7748 11840 7800 11892
rect 3700 11679 3752 11688
rect 3700 11645 3734 11679
rect 3734 11645 3752 11679
rect 3700 11636 3752 11645
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 6092 11772 6144 11824
rect 6920 11772 6972 11824
rect 7656 11772 7708 11824
rect 9588 11840 9640 11892
rect 9772 11840 9824 11892
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 6000 11636 6052 11645
rect 1032 11500 1084 11552
rect 1768 11500 1820 11552
rect 4252 11500 4304 11552
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 6644 11568 6696 11620
rect 7840 11679 7892 11688
rect 7840 11645 7849 11679
rect 7849 11645 7883 11679
rect 7883 11645 7892 11679
rect 7840 11636 7892 11645
rect 8024 11636 8076 11688
rect 7748 11611 7800 11620
rect 7748 11577 7757 11611
rect 7757 11577 7791 11611
rect 7791 11577 7800 11611
rect 7748 11568 7800 11577
rect 6828 11500 6880 11552
rect 9496 11636 9548 11688
rect 9772 11679 9824 11688
rect 9772 11645 9781 11679
rect 9781 11645 9815 11679
rect 9815 11645 9824 11679
rect 9772 11636 9824 11645
rect 14832 11840 14884 11892
rect 16764 11840 16816 11892
rect 19064 11840 19116 11892
rect 19616 11840 19668 11892
rect 11980 11772 12032 11824
rect 16488 11772 16540 11824
rect 16948 11772 17000 11824
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 11796 11636 11848 11688
rect 11888 11679 11940 11688
rect 11888 11645 11897 11679
rect 11897 11645 11931 11679
rect 11931 11645 11940 11679
rect 11888 11636 11940 11645
rect 11980 11679 12032 11688
rect 11980 11645 11989 11679
rect 11989 11645 12023 11679
rect 12023 11645 12032 11679
rect 11980 11636 12032 11645
rect 14096 11704 14148 11756
rect 10232 11611 10284 11620
rect 10232 11577 10266 11611
rect 10266 11577 10284 11611
rect 10232 11568 10284 11577
rect 11428 11568 11480 11620
rect 8116 11543 8168 11552
rect 8116 11509 8125 11543
rect 8125 11509 8159 11543
rect 8159 11509 8168 11543
rect 8116 11500 8168 11509
rect 8484 11500 8536 11552
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 11244 11500 11296 11552
rect 11520 11500 11572 11552
rect 12900 11568 12952 11620
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 13912 11679 13964 11688
rect 13912 11645 13921 11679
rect 13921 11645 13955 11679
rect 13955 11645 13964 11679
rect 13912 11636 13964 11645
rect 14004 11636 14056 11688
rect 14648 11636 14700 11688
rect 14280 11568 14332 11620
rect 14740 11568 14792 11620
rect 15016 11500 15068 11552
rect 16580 11704 16632 11756
rect 17224 11704 17276 11756
rect 18604 11704 18656 11756
rect 19156 11704 19208 11756
rect 15568 11568 15620 11620
rect 16948 11636 17000 11688
rect 18236 11636 18288 11688
rect 17408 11568 17460 11620
rect 17960 11568 18012 11620
rect 18420 11636 18472 11688
rect 18880 11679 18932 11688
rect 18880 11645 18889 11679
rect 18889 11645 18923 11679
rect 18923 11645 18932 11679
rect 18880 11636 18932 11645
rect 17868 11500 17920 11552
rect 18420 11500 18472 11552
rect 19708 11679 19760 11688
rect 19708 11645 19728 11679
rect 19728 11645 19760 11679
rect 19708 11636 19760 11645
rect 20352 11679 20404 11688
rect 20352 11645 20361 11679
rect 20361 11645 20395 11679
rect 20395 11645 20404 11679
rect 20352 11636 20404 11645
rect 20812 11840 20864 11892
rect 29000 11840 29052 11892
rect 29184 11840 29236 11892
rect 19800 11568 19852 11620
rect 19156 11500 19208 11552
rect 19616 11500 19668 11552
rect 20904 11636 20956 11688
rect 22008 11772 22060 11824
rect 22836 11772 22888 11824
rect 21640 11747 21692 11756
rect 21640 11713 21649 11747
rect 21649 11713 21683 11747
rect 21683 11713 21692 11747
rect 21640 11704 21692 11713
rect 23296 11772 23348 11824
rect 24032 11772 24084 11824
rect 23572 11747 23624 11756
rect 21456 11636 21508 11688
rect 22560 11679 22612 11688
rect 22560 11645 22569 11679
rect 22569 11645 22603 11679
rect 22603 11645 22612 11679
rect 22560 11636 22612 11645
rect 23572 11713 23581 11747
rect 23581 11713 23615 11747
rect 23615 11713 23624 11747
rect 23572 11704 23624 11713
rect 23480 11636 23532 11688
rect 23848 11704 23900 11756
rect 24768 11704 24820 11756
rect 28172 11704 28224 11756
rect 22284 11500 22336 11552
rect 22836 11500 22888 11552
rect 23940 11636 23992 11688
rect 24032 11568 24084 11620
rect 24584 11568 24636 11620
rect 24860 11500 24912 11552
rect 26240 11636 26292 11688
rect 26976 11636 27028 11688
rect 29276 11704 29328 11756
rect 25964 11568 26016 11620
rect 27252 11611 27304 11620
rect 27252 11577 27270 11611
rect 27270 11577 27304 11611
rect 27252 11568 27304 11577
rect 27988 11568 28040 11620
rect 29828 11636 29880 11688
rect 30288 11636 30340 11688
rect 30380 11568 30432 11620
rect 28448 11500 28500 11552
rect 29000 11500 29052 11552
rect 8102 11398 8154 11450
rect 8166 11398 8218 11450
rect 8230 11398 8282 11450
rect 8294 11398 8346 11450
rect 8358 11398 8410 11450
rect 15807 11398 15859 11450
rect 15871 11398 15923 11450
rect 15935 11398 15987 11450
rect 15999 11398 16051 11450
rect 16063 11398 16115 11450
rect 23512 11398 23564 11450
rect 23576 11398 23628 11450
rect 23640 11398 23692 11450
rect 23704 11398 23756 11450
rect 23768 11398 23820 11450
rect 31217 11398 31269 11450
rect 31281 11398 31333 11450
rect 31345 11398 31397 11450
rect 31409 11398 31461 11450
rect 31473 11398 31525 11450
rect 1676 11296 1728 11348
rect 3332 11296 3384 11348
rect 4252 11296 4304 11348
rect 6092 11296 6144 11348
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 7012 11296 7064 11348
rect 1400 11160 1452 11212
rect 3608 11203 3660 11212
rect 3608 11169 3642 11203
rect 3642 11169 3660 11203
rect 3608 11160 3660 11169
rect 5264 11203 5316 11212
rect 5264 11169 5273 11203
rect 5273 11169 5307 11203
rect 5307 11169 5316 11203
rect 5264 11160 5316 11169
rect 5724 11160 5776 11212
rect 2688 10999 2740 11008
rect 2688 10965 2697 10999
rect 2697 10965 2731 10999
rect 2731 10965 2740 10999
rect 2688 10956 2740 10965
rect 6184 11271 6236 11280
rect 6184 11237 6193 11271
rect 6193 11237 6227 11271
rect 6227 11237 6236 11271
rect 6184 11228 6236 11237
rect 8300 11228 8352 11280
rect 6828 11160 6880 11212
rect 8116 11160 8168 11212
rect 8576 11092 8628 11144
rect 11336 11228 11388 11280
rect 11612 11228 11664 11280
rect 14280 11296 14332 11348
rect 16028 11296 16080 11348
rect 9772 11092 9824 11144
rect 10140 11092 10192 11144
rect 9496 11024 9548 11076
rect 9588 11067 9640 11076
rect 9588 11033 9597 11067
rect 9597 11033 9631 11067
rect 9631 11033 9640 11067
rect 9588 11024 9640 11033
rect 10784 11203 10836 11212
rect 10784 11169 10793 11203
rect 10793 11169 10827 11203
rect 10827 11169 10836 11203
rect 10784 11160 10836 11169
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 12900 11160 12952 11212
rect 7196 10956 7248 11008
rect 9404 10956 9456 11008
rect 10048 10956 10100 11008
rect 10140 10999 10192 11008
rect 10140 10965 10149 10999
rect 10149 10965 10183 10999
rect 10183 10965 10192 10999
rect 10140 10956 10192 10965
rect 10232 10956 10284 11008
rect 11888 10956 11940 11008
rect 12072 10999 12124 11008
rect 12072 10965 12081 10999
rect 12081 10965 12115 10999
rect 12115 10965 12124 10999
rect 12072 10956 12124 10965
rect 16672 11296 16724 11348
rect 17224 11296 17276 11348
rect 14188 11203 14240 11212
rect 14188 11169 14197 11203
rect 14197 11169 14231 11203
rect 14231 11169 14240 11203
rect 14188 11160 14240 11169
rect 17500 11296 17552 11348
rect 17684 11296 17736 11348
rect 17776 11296 17828 11348
rect 17868 11296 17920 11348
rect 20076 11296 20128 11348
rect 13544 11092 13596 11144
rect 15844 11024 15896 11076
rect 16672 11203 16724 11212
rect 16672 11169 16681 11203
rect 16681 11169 16715 11203
rect 16715 11169 16724 11203
rect 16672 11160 16724 11169
rect 16856 11160 16908 11212
rect 17040 11203 17092 11212
rect 17040 11169 17049 11203
rect 17049 11169 17083 11203
rect 17083 11169 17092 11203
rect 17040 11160 17092 11169
rect 17408 11203 17460 11212
rect 17408 11169 17417 11203
rect 17417 11169 17451 11203
rect 17451 11169 17460 11203
rect 17408 11160 17460 11169
rect 18052 11228 18104 11280
rect 19156 11228 19208 11280
rect 17868 11203 17920 11212
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 18236 11160 18288 11212
rect 23204 11296 23256 11348
rect 24400 11296 24452 11348
rect 27252 11339 27304 11348
rect 27252 11305 27261 11339
rect 27261 11305 27295 11339
rect 27295 11305 27304 11339
rect 27252 11296 27304 11305
rect 28172 11296 28224 11348
rect 28448 11296 28500 11348
rect 21272 11228 21324 11280
rect 22192 11228 22244 11280
rect 20996 11160 21048 11212
rect 22008 11160 22060 11212
rect 22560 11160 22612 11212
rect 22744 11203 22796 11212
rect 22744 11169 22753 11203
rect 22753 11169 22787 11203
rect 22787 11169 22796 11203
rect 22744 11160 22796 11169
rect 26240 11228 26292 11280
rect 17500 11092 17552 11144
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 18972 11092 19024 11144
rect 19156 11092 19208 11144
rect 25504 11203 25556 11212
rect 25504 11169 25513 11203
rect 25513 11169 25547 11203
rect 25547 11169 25556 11203
rect 25504 11160 25556 11169
rect 28080 11228 28132 11280
rect 29276 11296 29328 11348
rect 26424 11092 26476 11144
rect 27252 11092 27304 11144
rect 14464 10956 14516 11008
rect 17040 11024 17092 11076
rect 20812 11024 20864 11076
rect 24676 11024 24728 11076
rect 27988 11024 28040 11076
rect 16028 10956 16080 11008
rect 16304 10956 16356 11008
rect 18328 10956 18380 11008
rect 18972 10956 19024 11008
rect 20076 10956 20128 11008
rect 21456 10956 21508 11008
rect 25596 10999 25648 11008
rect 25596 10965 25605 10999
rect 25605 10965 25639 10999
rect 25639 10965 25648 10999
rect 25596 10956 25648 10965
rect 26792 10956 26844 11008
rect 28448 10956 28500 11008
rect 30288 11160 30340 11212
rect 30656 11203 30708 11212
rect 30656 11169 30674 11203
rect 30674 11169 30708 11203
rect 30656 11160 30708 11169
rect 4250 10854 4302 10906
rect 4314 10854 4366 10906
rect 4378 10854 4430 10906
rect 4442 10854 4494 10906
rect 4506 10854 4558 10906
rect 11955 10854 12007 10906
rect 12019 10854 12071 10906
rect 12083 10854 12135 10906
rect 12147 10854 12199 10906
rect 12211 10854 12263 10906
rect 19660 10854 19712 10906
rect 19724 10854 19776 10906
rect 19788 10854 19840 10906
rect 19852 10854 19904 10906
rect 19916 10854 19968 10906
rect 27365 10854 27417 10906
rect 27429 10854 27481 10906
rect 27493 10854 27545 10906
rect 27557 10854 27609 10906
rect 27621 10854 27673 10906
rect 1768 10752 1820 10804
rect 5264 10752 5316 10804
rect 5632 10752 5684 10804
rect 1032 10616 1084 10668
rect 1400 10616 1452 10668
rect 1492 10480 1544 10532
rect 2688 10548 2740 10600
rect 4252 10591 4304 10600
rect 4252 10557 4261 10591
rect 4261 10557 4295 10591
rect 4295 10557 4304 10591
rect 4252 10548 4304 10557
rect 5448 10684 5500 10736
rect 7748 10684 7800 10736
rect 3516 10480 3568 10532
rect 7196 10548 7248 10600
rect 7748 10548 7800 10600
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 4160 10412 4212 10421
rect 4528 10412 4580 10464
rect 7104 10480 7156 10532
rect 7932 10412 7984 10464
rect 8576 10591 8628 10600
rect 8576 10557 8585 10591
rect 8585 10557 8619 10591
rect 8619 10557 8628 10591
rect 8576 10548 8628 10557
rect 9496 10752 9548 10804
rect 13176 10752 13228 10804
rect 14464 10752 14516 10804
rect 14740 10795 14792 10804
rect 14740 10761 14749 10795
rect 14749 10761 14783 10795
rect 14783 10761 14792 10795
rect 14740 10752 14792 10761
rect 14924 10752 14976 10804
rect 15660 10795 15712 10804
rect 15660 10761 15669 10795
rect 15669 10761 15703 10795
rect 15703 10761 15712 10795
rect 15660 10752 15712 10761
rect 16028 10752 16080 10804
rect 16396 10752 16448 10804
rect 16672 10752 16724 10804
rect 17040 10752 17092 10804
rect 17316 10752 17368 10804
rect 17684 10752 17736 10804
rect 18788 10752 18840 10804
rect 20352 10795 20404 10804
rect 20352 10761 20361 10795
rect 20361 10761 20395 10795
rect 20395 10761 20404 10795
rect 20352 10752 20404 10761
rect 22100 10752 22152 10804
rect 25688 10795 25740 10804
rect 25688 10761 25697 10795
rect 25697 10761 25731 10795
rect 25731 10761 25740 10795
rect 25688 10752 25740 10761
rect 25964 10795 26016 10804
rect 25964 10761 25973 10795
rect 25973 10761 26007 10795
rect 26007 10761 26016 10795
rect 25964 10752 26016 10761
rect 26424 10795 26476 10804
rect 26424 10761 26433 10795
rect 26433 10761 26467 10795
rect 26467 10761 26476 10795
rect 26424 10752 26476 10761
rect 27252 10795 27304 10804
rect 27252 10761 27261 10795
rect 27261 10761 27295 10795
rect 27295 10761 27304 10795
rect 27252 10752 27304 10761
rect 28080 10795 28132 10804
rect 28080 10761 28089 10795
rect 28089 10761 28123 10795
rect 28123 10761 28132 10795
rect 28080 10752 28132 10761
rect 28172 10752 28224 10804
rect 28816 10752 28868 10804
rect 29460 10795 29512 10804
rect 29460 10761 29469 10795
rect 29469 10761 29503 10795
rect 29503 10761 29512 10795
rect 29460 10752 29512 10761
rect 30656 10752 30708 10804
rect 10140 10616 10192 10668
rect 8668 10523 8720 10532
rect 8668 10489 8677 10523
rect 8677 10489 8711 10523
rect 8711 10489 8720 10523
rect 8668 10480 8720 10489
rect 9128 10548 9180 10600
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 10784 10591 10836 10600
rect 10784 10557 10793 10591
rect 10793 10557 10827 10591
rect 10827 10557 10836 10591
rect 10784 10548 10836 10557
rect 11888 10548 11940 10600
rect 13912 10684 13964 10736
rect 17132 10684 17184 10736
rect 8760 10412 8812 10464
rect 12532 10523 12584 10532
rect 12532 10489 12541 10523
rect 12541 10489 12575 10523
rect 12575 10489 12584 10523
rect 12532 10480 12584 10489
rect 12624 10480 12676 10532
rect 10232 10455 10284 10464
rect 10232 10421 10241 10455
rect 10241 10421 10275 10455
rect 10275 10421 10284 10455
rect 10232 10412 10284 10421
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 14096 10455 14148 10464
rect 14096 10421 14105 10455
rect 14105 10421 14139 10455
rect 14139 10421 14148 10455
rect 14096 10412 14148 10421
rect 14372 10480 14424 10532
rect 14556 10523 14608 10532
rect 14556 10489 14565 10523
rect 14565 10489 14599 10523
rect 14599 10489 14608 10523
rect 14556 10480 14608 10489
rect 14740 10523 14792 10532
rect 15844 10548 15896 10600
rect 15936 10591 15988 10600
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 16120 10616 16172 10668
rect 16856 10616 16908 10668
rect 17408 10616 17460 10668
rect 14740 10489 14765 10523
rect 14765 10489 14792 10523
rect 14740 10480 14792 10489
rect 15476 10523 15528 10532
rect 15476 10489 15485 10523
rect 15485 10489 15519 10523
rect 15519 10489 15528 10523
rect 15476 10480 15528 10489
rect 16396 10591 16448 10600
rect 16396 10557 16410 10591
rect 16410 10557 16444 10591
rect 16444 10557 16448 10591
rect 16396 10548 16448 10557
rect 16672 10523 16724 10532
rect 16672 10489 16681 10523
rect 16681 10489 16715 10523
rect 16715 10489 16724 10523
rect 16672 10480 16724 10489
rect 14924 10455 14976 10464
rect 14924 10421 14933 10455
rect 14933 10421 14967 10455
rect 14967 10421 14976 10455
rect 14924 10412 14976 10421
rect 15200 10455 15252 10464
rect 15200 10421 15225 10455
rect 15225 10421 15252 10455
rect 15200 10412 15252 10421
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 16304 10412 16356 10464
rect 17040 10455 17092 10464
rect 17040 10421 17049 10455
rect 17049 10421 17083 10455
rect 17083 10421 17092 10455
rect 17040 10412 17092 10421
rect 17224 10412 17276 10464
rect 17316 10412 17368 10464
rect 18144 10523 18196 10532
rect 18144 10489 18153 10523
rect 18153 10489 18187 10523
rect 18187 10489 18196 10523
rect 18144 10480 18196 10489
rect 17776 10412 17828 10464
rect 19248 10616 19300 10668
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 19800 10591 19852 10600
rect 19800 10557 19810 10591
rect 19810 10557 19844 10591
rect 19844 10557 19852 10591
rect 19800 10548 19852 10557
rect 20076 10591 20128 10600
rect 20076 10557 20085 10591
rect 20085 10557 20119 10591
rect 20119 10557 20128 10591
rect 20076 10548 20128 10557
rect 21272 10616 21324 10668
rect 22192 10616 22244 10668
rect 22836 10548 22888 10600
rect 25412 10548 25464 10600
rect 25964 10616 26016 10668
rect 21548 10480 21600 10532
rect 21732 10523 21784 10532
rect 21732 10489 21741 10523
rect 21741 10489 21775 10523
rect 21775 10489 21784 10523
rect 21732 10480 21784 10489
rect 18512 10455 18564 10464
rect 18512 10421 18521 10455
rect 18521 10421 18555 10455
rect 18555 10421 18564 10455
rect 18512 10412 18564 10421
rect 22192 10412 22244 10464
rect 23848 10412 23900 10464
rect 25504 10412 25556 10464
rect 25688 10412 25740 10464
rect 26424 10548 26476 10600
rect 27252 10616 27304 10668
rect 26792 10548 26844 10600
rect 28448 10591 28500 10600
rect 28448 10557 28457 10591
rect 28457 10557 28491 10591
rect 28491 10557 28500 10591
rect 28448 10548 28500 10557
rect 29092 10591 29144 10600
rect 29092 10557 29101 10591
rect 29101 10557 29135 10591
rect 29135 10557 29144 10591
rect 29092 10548 29144 10557
rect 29276 10548 29328 10600
rect 30380 10616 30432 10668
rect 31668 10548 31720 10600
rect 29000 10480 29052 10532
rect 29920 10480 29972 10532
rect 8102 10310 8154 10362
rect 8166 10310 8218 10362
rect 8230 10310 8282 10362
rect 8294 10310 8346 10362
rect 8358 10310 8410 10362
rect 15807 10310 15859 10362
rect 15871 10310 15923 10362
rect 15935 10310 15987 10362
rect 15999 10310 16051 10362
rect 16063 10310 16115 10362
rect 23512 10310 23564 10362
rect 23576 10310 23628 10362
rect 23640 10310 23692 10362
rect 23704 10310 23756 10362
rect 23768 10310 23820 10362
rect 31217 10310 31269 10362
rect 31281 10310 31333 10362
rect 31345 10310 31397 10362
rect 31409 10310 31461 10362
rect 31473 10310 31525 10362
rect 1400 10208 1452 10260
rect 1308 10140 1360 10192
rect 1492 10115 1544 10124
rect 1492 10081 1501 10115
rect 1501 10081 1535 10115
rect 1535 10081 1544 10115
rect 1492 10072 1544 10081
rect 1676 10072 1728 10124
rect 3608 10140 3660 10192
rect 3700 10183 3752 10192
rect 3700 10149 3709 10183
rect 3709 10149 3743 10183
rect 3743 10149 3752 10183
rect 3700 10140 3752 10149
rect 3792 10115 3844 10124
rect 3792 10081 3801 10115
rect 3801 10081 3835 10115
rect 3835 10081 3844 10115
rect 3792 10072 3844 10081
rect 4252 10140 4304 10192
rect 4068 10004 4120 10056
rect 4712 10115 4764 10124
rect 4712 10081 4721 10115
rect 4721 10081 4755 10115
rect 4755 10081 4764 10115
rect 4712 10072 4764 10081
rect 7472 10140 7524 10192
rect 7840 10140 7892 10192
rect 9588 10183 9640 10192
rect 9588 10149 9622 10183
rect 9622 10149 9640 10183
rect 9588 10140 9640 10149
rect 7748 10072 7800 10124
rect 4160 9936 4212 9988
rect 4988 9936 5040 9988
rect 1216 9868 1268 9920
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 8668 10004 8720 10056
rect 13912 10140 13964 10192
rect 11796 10072 11848 10124
rect 11980 10072 12032 10124
rect 13728 10072 13780 10124
rect 14188 10115 14240 10124
rect 14188 10081 14197 10115
rect 14197 10081 14231 10115
rect 14231 10081 14240 10115
rect 14188 10072 14240 10081
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 13268 9979 13320 9988
rect 13268 9945 13277 9979
rect 13277 9945 13311 9979
rect 13311 9945 13320 9979
rect 13268 9936 13320 9945
rect 14740 10004 14792 10056
rect 15292 10004 15344 10056
rect 15568 10115 15620 10124
rect 15568 10081 15577 10115
rect 15577 10081 15611 10115
rect 15611 10081 15620 10115
rect 15568 10072 15620 10081
rect 15752 10072 15804 10124
rect 16948 10072 17000 10124
rect 21272 10208 21324 10260
rect 22008 10208 22060 10260
rect 22100 10251 22152 10260
rect 22100 10217 22109 10251
rect 22109 10217 22143 10251
rect 22143 10217 22152 10251
rect 22100 10208 22152 10217
rect 22744 10208 22796 10260
rect 22836 10208 22888 10260
rect 23848 10251 23900 10260
rect 23848 10217 23857 10251
rect 23857 10217 23891 10251
rect 23891 10217 23900 10251
rect 23848 10208 23900 10217
rect 25688 10208 25740 10260
rect 26884 10251 26936 10260
rect 26884 10217 26893 10251
rect 26893 10217 26927 10251
rect 26927 10217 26936 10251
rect 26884 10208 26936 10217
rect 29276 10208 29328 10260
rect 30380 10208 30432 10260
rect 20444 10140 20496 10192
rect 21916 10140 21968 10192
rect 17960 10115 18012 10124
rect 17960 10081 17969 10115
rect 17969 10081 18003 10115
rect 18003 10081 18012 10115
rect 17960 10072 18012 10081
rect 7564 9911 7616 9920
rect 7564 9877 7573 9911
rect 7573 9877 7607 9911
rect 7607 9877 7616 9911
rect 7564 9868 7616 9877
rect 13544 9911 13596 9920
rect 13544 9877 13553 9911
rect 13553 9877 13587 9911
rect 13587 9877 13596 9911
rect 13544 9868 13596 9877
rect 13728 9911 13780 9920
rect 13728 9877 13737 9911
rect 13737 9877 13771 9911
rect 13771 9877 13780 9911
rect 13728 9868 13780 9877
rect 14096 9868 14148 9920
rect 14556 9868 14608 9920
rect 14648 9868 14700 9920
rect 14740 9911 14792 9920
rect 14740 9877 14749 9911
rect 14749 9877 14783 9911
rect 14783 9877 14792 9911
rect 14740 9868 14792 9877
rect 14832 9911 14884 9920
rect 14832 9877 14841 9911
rect 14841 9877 14875 9911
rect 14875 9877 14884 9911
rect 14832 9868 14884 9877
rect 15384 9868 15436 9920
rect 16580 9868 16632 9920
rect 18328 10115 18380 10124
rect 18328 10081 18337 10115
rect 18337 10081 18371 10115
rect 18371 10081 18380 10115
rect 18328 10072 18380 10081
rect 18236 10004 18288 10056
rect 18880 9936 18932 9988
rect 19984 10072 20036 10124
rect 20996 10115 21048 10124
rect 20996 10081 21005 10115
rect 21005 10081 21039 10115
rect 21039 10081 21048 10115
rect 20996 10072 21048 10081
rect 21640 10115 21692 10124
rect 21640 10081 21649 10115
rect 21649 10081 21683 10115
rect 21683 10081 21692 10115
rect 21640 10072 21692 10081
rect 21732 10115 21784 10124
rect 21732 10081 21741 10115
rect 21741 10081 21775 10115
rect 21775 10081 21784 10115
rect 21732 10072 21784 10081
rect 22192 10115 22244 10124
rect 22192 10081 22201 10115
rect 22201 10081 22235 10115
rect 22235 10081 22244 10115
rect 22192 10072 22244 10081
rect 22284 10115 22336 10124
rect 22284 10081 22293 10115
rect 22293 10081 22327 10115
rect 22327 10081 22336 10115
rect 22284 10072 22336 10081
rect 22560 10115 22612 10124
rect 22560 10081 22569 10115
rect 22569 10081 22603 10115
rect 22603 10081 22612 10115
rect 22560 10072 22612 10081
rect 25504 10183 25556 10192
rect 25504 10149 25513 10183
rect 25513 10149 25547 10183
rect 25547 10149 25556 10183
rect 25504 10140 25556 10149
rect 21548 9936 21600 9988
rect 23388 10004 23440 10056
rect 24492 10072 24544 10124
rect 25412 10115 25464 10124
rect 25412 10081 25421 10115
rect 25421 10081 25455 10115
rect 25455 10081 25464 10115
rect 25412 10072 25464 10081
rect 27988 10183 28040 10192
rect 27988 10149 28006 10183
rect 28006 10149 28040 10183
rect 28908 10183 28960 10192
rect 27988 10140 28040 10149
rect 28908 10149 28917 10183
rect 28917 10149 28951 10183
rect 28951 10149 28960 10183
rect 28908 10140 28960 10149
rect 28816 10115 28868 10124
rect 28816 10081 28825 10115
rect 28825 10081 28859 10115
rect 28859 10081 28868 10115
rect 28816 10072 28868 10081
rect 30288 10140 30340 10192
rect 29920 10072 29972 10124
rect 25596 10004 25648 10056
rect 29368 10047 29420 10056
rect 29368 10013 29377 10047
rect 29377 10013 29411 10047
rect 29411 10013 29420 10047
rect 29368 10004 29420 10013
rect 23204 9979 23256 9988
rect 23204 9945 23213 9979
rect 23213 9945 23247 9979
rect 23247 9945 23256 9979
rect 23204 9936 23256 9945
rect 24032 9936 24084 9988
rect 23848 9868 23900 9920
rect 24400 9868 24452 9920
rect 29184 9911 29236 9920
rect 29184 9877 29193 9911
rect 29193 9877 29227 9911
rect 29227 9877 29236 9911
rect 29184 9868 29236 9877
rect 4250 9766 4302 9818
rect 4314 9766 4366 9818
rect 4378 9766 4430 9818
rect 4442 9766 4494 9818
rect 4506 9766 4558 9818
rect 11955 9766 12007 9818
rect 12019 9766 12071 9818
rect 12083 9766 12135 9818
rect 12147 9766 12199 9818
rect 12211 9766 12263 9818
rect 19660 9766 19712 9818
rect 19724 9766 19776 9818
rect 19788 9766 19840 9818
rect 19852 9766 19904 9818
rect 19916 9766 19968 9818
rect 27365 9766 27417 9818
rect 27429 9766 27481 9818
rect 27493 9766 27545 9818
rect 27557 9766 27609 9818
rect 27621 9766 27673 9818
rect 1584 9664 1636 9716
rect 1768 9596 1820 9648
rect 3792 9707 3844 9716
rect 3792 9673 3801 9707
rect 3801 9673 3835 9707
rect 3835 9673 3844 9707
rect 3792 9664 3844 9673
rect 4068 9707 4120 9716
rect 4068 9673 4077 9707
rect 4077 9673 4111 9707
rect 4111 9673 4120 9707
rect 4068 9664 4120 9673
rect 1216 9528 1268 9580
rect 4712 9664 4764 9716
rect 8760 9664 8812 9716
rect 12532 9664 12584 9716
rect 13728 9664 13780 9716
rect 13912 9664 13964 9716
rect 14648 9707 14700 9716
rect 14648 9673 14657 9707
rect 14657 9673 14691 9707
rect 14691 9673 14700 9707
rect 14648 9664 14700 9673
rect 3608 9460 3660 9512
rect 3792 9460 3844 9512
rect 4988 9460 5040 9512
rect 7104 9460 7156 9512
rect 7472 9460 7524 9512
rect 7564 9460 7616 9512
rect 7840 9460 7892 9512
rect 10968 9460 11020 9512
rect 11612 9460 11664 9512
rect 11704 9460 11756 9512
rect 12256 9528 12308 9580
rect 13176 9528 13228 9580
rect 14832 9664 14884 9716
rect 14924 9664 14976 9716
rect 15108 9707 15160 9716
rect 15108 9673 15117 9707
rect 15117 9673 15151 9707
rect 15151 9673 15160 9707
rect 15108 9664 15160 9673
rect 16580 9707 16632 9716
rect 16580 9673 16589 9707
rect 16589 9673 16623 9707
rect 16623 9673 16632 9707
rect 16580 9664 16632 9673
rect 16856 9664 16908 9716
rect 17040 9664 17092 9716
rect 17132 9707 17184 9716
rect 17132 9673 17141 9707
rect 17141 9673 17175 9707
rect 17175 9673 17184 9707
rect 17132 9664 17184 9673
rect 17224 9664 17276 9716
rect 17592 9664 17644 9716
rect 15108 9528 15160 9580
rect 12348 9503 12400 9512
rect 1400 9324 1452 9376
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 3240 9324 3292 9376
rect 4160 9324 4212 9376
rect 6276 9367 6328 9376
rect 6276 9333 6285 9367
rect 6285 9333 6319 9367
rect 6319 9333 6328 9367
rect 6276 9324 6328 9333
rect 6736 9367 6788 9376
rect 6736 9333 6745 9367
rect 6745 9333 6779 9367
rect 6779 9333 6788 9367
rect 6736 9324 6788 9333
rect 7656 9324 7708 9376
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 8484 9324 8536 9376
rect 11888 9392 11940 9444
rect 11336 9324 11388 9376
rect 12348 9469 12357 9503
rect 12357 9469 12391 9503
rect 12391 9469 12400 9503
rect 12348 9460 12400 9469
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 13452 9460 13504 9512
rect 12072 9392 12124 9444
rect 14832 9503 14884 9512
rect 14832 9469 14841 9503
rect 14841 9469 14875 9503
rect 14875 9469 14884 9503
rect 14832 9460 14884 9469
rect 15200 9392 15252 9444
rect 15384 9503 15436 9512
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 15384 9460 15436 9469
rect 15660 9460 15712 9512
rect 15752 9392 15804 9444
rect 16396 9503 16448 9512
rect 16396 9469 16429 9503
rect 16429 9469 16448 9503
rect 16396 9460 16448 9469
rect 16120 9392 16172 9444
rect 14740 9324 14792 9376
rect 14832 9324 14884 9376
rect 16948 9460 17000 9512
rect 17132 9460 17184 9512
rect 16856 9324 16908 9376
rect 17316 9324 17368 9376
rect 18236 9596 18288 9648
rect 18512 9596 18564 9648
rect 19524 9596 19576 9648
rect 19708 9596 19760 9648
rect 20536 9664 20588 9716
rect 17776 9503 17828 9506
rect 17776 9469 17785 9503
rect 17785 9469 17819 9503
rect 17819 9469 17828 9503
rect 17776 9454 17828 9469
rect 19340 9503 19392 9512
rect 19340 9469 19349 9503
rect 19349 9469 19383 9503
rect 19383 9469 19392 9503
rect 19340 9460 19392 9469
rect 18328 9392 18380 9444
rect 19524 9392 19576 9444
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 20812 9596 20864 9648
rect 21272 9664 21324 9716
rect 21640 9664 21692 9716
rect 22560 9664 22612 9716
rect 28908 9664 28960 9716
rect 29092 9639 29144 9648
rect 29092 9605 29101 9639
rect 29101 9605 29135 9639
rect 29135 9605 29144 9639
rect 29092 9596 29144 9605
rect 20444 9503 20496 9512
rect 20444 9469 20453 9503
rect 20453 9469 20487 9503
rect 20487 9469 20496 9503
rect 20444 9460 20496 9469
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 20352 9392 20404 9444
rect 20904 9503 20956 9512
rect 20904 9469 20913 9503
rect 20913 9469 20947 9503
rect 20947 9469 20956 9503
rect 20904 9460 20956 9469
rect 22192 9503 22244 9512
rect 22192 9469 22201 9503
rect 22201 9469 22235 9503
rect 22235 9469 22244 9503
rect 22192 9460 22244 9469
rect 21088 9392 21140 9444
rect 22100 9392 22152 9444
rect 22468 9460 22520 9512
rect 22560 9503 22612 9512
rect 22560 9469 22569 9503
rect 22569 9469 22603 9503
rect 22603 9469 22612 9503
rect 22560 9460 22612 9469
rect 24124 9503 24176 9512
rect 24124 9469 24133 9503
rect 24133 9469 24167 9503
rect 24167 9469 24176 9503
rect 24124 9460 24176 9469
rect 25688 9571 25740 9580
rect 25688 9537 25697 9571
rect 25697 9537 25731 9571
rect 25731 9537 25740 9571
rect 25688 9528 25740 9537
rect 24492 9503 24544 9512
rect 24492 9469 24501 9503
rect 24501 9469 24535 9503
rect 24535 9469 24544 9503
rect 24492 9460 24544 9469
rect 24676 9460 24728 9512
rect 24584 9392 24636 9444
rect 22284 9324 22336 9376
rect 22376 9367 22428 9376
rect 22376 9333 22385 9367
rect 22385 9333 22419 9367
rect 22419 9333 22428 9367
rect 22376 9324 22428 9333
rect 27896 9460 27948 9512
rect 26792 9392 26844 9444
rect 29460 9503 29512 9512
rect 29460 9469 29469 9503
rect 29469 9469 29503 9503
rect 29503 9469 29512 9503
rect 29460 9460 29512 9469
rect 30288 9707 30340 9716
rect 30288 9673 30297 9707
rect 30297 9673 30331 9707
rect 30331 9673 30340 9707
rect 30288 9664 30340 9673
rect 30288 9460 30340 9512
rect 29184 9324 29236 9376
rect 8102 9222 8154 9274
rect 8166 9222 8218 9274
rect 8230 9222 8282 9274
rect 8294 9222 8346 9274
rect 8358 9222 8410 9274
rect 15807 9222 15859 9274
rect 15871 9222 15923 9274
rect 15935 9222 15987 9274
rect 15999 9222 16051 9274
rect 16063 9222 16115 9274
rect 23512 9222 23564 9274
rect 23576 9222 23628 9274
rect 23640 9222 23692 9274
rect 23704 9222 23756 9274
rect 23768 9222 23820 9274
rect 31217 9222 31269 9274
rect 31281 9222 31333 9274
rect 31345 9222 31397 9274
rect 31409 9222 31461 9274
rect 31473 9222 31525 9274
rect 1400 9120 1452 9172
rect 2136 9120 2188 9172
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 3608 9120 3660 9172
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 6276 9120 6328 9172
rect 6644 9052 6696 9104
rect 6736 9052 6788 9104
rect 2596 9027 2648 9036
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 2596 8993 2605 9027
rect 2605 8993 2639 9027
rect 2639 8993 2648 9027
rect 2596 8984 2648 8993
rect 2412 8916 2464 8968
rect 3792 8916 3844 8968
rect 7840 9052 7892 9104
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 12716 9120 12768 9172
rect 14188 9120 14240 9172
rect 14556 9120 14608 9172
rect 14924 9120 14976 9172
rect 15384 9120 15436 9172
rect 16120 9120 16172 9172
rect 7472 8916 7524 8968
rect 11612 8984 11664 9036
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 13084 8984 13136 9036
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 14556 8984 14608 9036
rect 16120 8984 16172 9036
rect 16672 9120 16724 9172
rect 4160 8780 4212 8832
rect 7012 8823 7064 8832
rect 7012 8789 7021 8823
rect 7021 8789 7055 8823
rect 7055 8789 7064 8823
rect 7012 8780 7064 8789
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 8392 8780 8444 8832
rect 8576 8780 8628 8832
rect 11520 8780 11572 8832
rect 15476 8916 15528 8968
rect 15660 8916 15712 8968
rect 13452 8891 13504 8900
rect 13452 8857 13461 8891
rect 13461 8857 13495 8891
rect 13495 8857 13504 8891
rect 13452 8848 13504 8857
rect 13544 8848 13596 8900
rect 15200 8848 15252 8900
rect 16304 8848 16356 8900
rect 19708 9120 19760 9172
rect 20536 9163 20588 9172
rect 20536 9129 20545 9163
rect 20545 9129 20579 9163
rect 20579 9129 20588 9163
rect 20536 9120 20588 9129
rect 22100 9120 22152 9172
rect 24860 9120 24912 9172
rect 16948 8984 17000 9036
rect 17592 9052 17644 9104
rect 17040 8916 17092 8968
rect 18052 9027 18104 9036
rect 18052 8993 18061 9027
rect 18061 8993 18095 9027
rect 18095 8993 18104 9027
rect 18052 8984 18104 8993
rect 18144 8984 18196 9036
rect 18328 9052 18380 9104
rect 18512 9095 18564 9104
rect 18512 9061 18539 9095
rect 18539 9061 18564 9095
rect 18512 9052 18564 9061
rect 18696 9095 18748 9104
rect 18696 9061 18705 9095
rect 18705 9061 18739 9095
rect 18739 9061 18748 9095
rect 18696 9052 18748 9061
rect 19984 9052 20036 9104
rect 24124 9052 24176 9104
rect 29368 9120 29420 9172
rect 30932 9163 30984 9172
rect 30932 9129 30941 9163
rect 30941 9129 30975 9163
rect 30975 9129 30984 9163
rect 30932 9120 30984 9129
rect 17960 8916 18012 8968
rect 18328 8916 18380 8968
rect 18696 8916 18748 8968
rect 16580 8848 16632 8900
rect 20628 8984 20680 9036
rect 20444 8916 20496 8968
rect 22100 9027 22152 9036
rect 22100 8993 22109 9027
rect 22109 8993 22143 9027
rect 22143 8993 22152 9027
rect 22100 8984 22152 8993
rect 12716 8780 12768 8832
rect 14280 8780 14332 8832
rect 14924 8780 14976 8832
rect 17040 8780 17092 8832
rect 17408 8780 17460 8832
rect 17592 8780 17644 8832
rect 17868 8823 17920 8832
rect 17868 8789 17877 8823
rect 17877 8789 17911 8823
rect 17911 8789 17920 8823
rect 17868 8780 17920 8789
rect 18512 8823 18564 8832
rect 18512 8789 18521 8823
rect 18521 8789 18555 8823
rect 18555 8789 18564 8823
rect 18512 8780 18564 8789
rect 19064 8780 19116 8832
rect 22008 8848 22060 8900
rect 22560 8984 22612 9036
rect 23480 8984 23532 9036
rect 23940 8984 23992 9036
rect 24400 8984 24452 9036
rect 26516 8984 26568 9036
rect 22468 8959 22520 8968
rect 22468 8925 22477 8959
rect 22477 8925 22511 8959
rect 22511 8925 22520 8959
rect 22468 8916 22520 8925
rect 27896 9027 27948 9036
rect 27896 8993 27905 9027
rect 27905 8993 27939 9027
rect 27939 8993 27948 9027
rect 27896 8984 27948 8993
rect 28724 8984 28776 9036
rect 23664 8848 23716 8900
rect 19892 8780 19944 8832
rect 22284 8780 22336 8832
rect 24124 8780 24176 8832
rect 25320 8823 25372 8832
rect 25320 8789 25329 8823
rect 25329 8789 25363 8823
rect 25363 8789 25372 8823
rect 25320 8780 25372 8789
rect 28448 8823 28500 8832
rect 28448 8789 28457 8823
rect 28457 8789 28491 8823
rect 28491 8789 28500 8823
rect 28448 8780 28500 8789
rect 28724 8823 28776 8832
rect 28724 8789 28733 8823
rect 28733 8789 28767 8823
rect 28767 8789 28776 8823
rect 28724 8780 28776 8789
rect 29092 9027 29144 9036
rect 29092 8993 29101 9027
rect 29101 8993 29135 9027
rect 29135 8993 29144 9027
rect 29092 8984 29144 8993
rect 29184 8984 29236 9036
rect 29184 8780 29236 8832
rect 4250 8678 4302 8730
rect 4314 8678 4366 8730
rect 4378 8678 4430 8730
rect 4442 8678 4494 8730
rect 4506 8678 4558 8730
rect 11955 8678 12007 8730
rect 12019 8678 12071 8730
rect 12083 8678 12135 8730
rect 12147 8678 12199 8730
rect 12211 8678 12263 8730
rect 19660 8678 19712 8730
rect 19724 8678 19776 8730
rect 19788 8678 19840 8730
rect 19852 8678 19904 8730
rect 19916 8678 19968 8730
rect 27365 8678 27417 8730
rect 27429 8678 27481 8730
rect 27493 8678 27545 8730
rect 27557 8678 27609 8730
rect 27621 8678 27673 8730
rect 1584 8576 1636 8628
rect 2412 8619 2464 8628
rect 1400 8440 1452 8492
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 2596 8576 2648 8628
rect 5724 8576 5776 8628
rect 7012 8576 7064 8628
rect 3700 8236 3752 8288
rect 4160 8236 4212 8288
rect 6368 8415 6420 8424
rect 6368 8381 6377 8415
rect 6377 8381 6411 8415
rect 6411 8381 6420 8415
rect 6368 8372 6420 8381
rect 5724 8304 5776 8356
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 7840 8440 7892 8492
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 10968 8372 11020 8424
rect 10232 8304 10284 8356
rect 12900 8576 12952 8628
rect 12992 8619 13044 8628
rect 12992 8585 13001 8619
rect 13001 8585 13035 8619
rect 13035 8585 13044 8619
rect 12992 8576 13044 8585
rect 13268 8576 13320 8628
rect 14556 8619 14608 8628
rect 14556 8585 14565 8619
rect 14565 8585 14599 8619
rect 14599 8585 14608 8619
rect 14556 8576 14608 8585
rect 15016 8576 15068 8628
rect 15844 8619 15896 8628
rect 15844 8585 15853 8619
rect 15853 8585 15887 8619
rect 15887 8585 15896 8619
rect 15844 8576 15896 8585
rect 16396 8576 16448 8628
rect 16764 8576 16816 8628
rect 17132 8576 17184 8628
rect 11888 8508 11940 8560
rect 13360 8508 13412 8560
rect 14188 8508 14240 8560
rect 16120 8508 16172 8560
rect 12348 8372 12400 8424
rect 12532 8372 12584 8424
rect 12716 8415 12768 8424
rect 12716 8381 12725 8415
rect 12725 8381 12759 8415
rect 12759 8381 12768 8415
rect 12716 8372 12768 8381
rect 13360 8372 13412 8424
rect 17776 8576 17828 8628
rect 18236 8576 18288 8628
rect 19984 8619 20036 8628
rect 19984 8585 19993 8619
rect 19993 8585 20027 8619
rect 20027 8585 20036 8619
rect 19984 8576 20036 8585
rect 21088 8576 21140 8628
rect 21732 8576 21784 8628
rect 22008 8576 22060 8628
rect 23480 8619 23532 8628
rect 23480 8585 23489 8619
rect 23489 8585 23523 8619
rect 23523 8585 23532 8619
rect 23480 8576 23532 8585
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 25320 8576 25372 8628
rect 26516 8619 26568 8628
rect 26516 8585 26525 8619
rect 26525 8585 26559 8619
rect 26559 8585 26568 8619
rect 26516 8576 26568 8585
rect 28448 8576 28500 8628
rect 29736 8576 29788 8628
rect 22652 8508 22704 8560
rect 17592 8440 17644 8492
rect 19524 8440 19576 8492
rect 19616 8440 19668 8492
rect 19892 8440 19944 8492
rect 20168 8440 20220 8492
rect 30012 8508 30064 8560
rect 13820 8415 13872 8424
rect 13820 8381 13829 8415
rect 13829 8381 13863 8415
rect 13863 8381 13872 8415
rect 13820 8372 13872 8381
rect 14188 8372 14240 8424
rect 14556 8372 14608 8424
rect 15384 8415 15436 8424
rect 15384 8381 15393 8415
rect 15393 8381 15427 8415
rect 15427 8381 15436 8415
rect 15384 8372 15436 8381
rect 15476 8415 15528 8424
rect 15476 8381 15485 8415
rect 15485 8381 15519 8415
rect 15519 8381 15528 8415
rect 15476 8372 15528 8381
rect 15844 8372 15896 8424
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 16948 8372 17000 8424
rect 16396 8304 16448 8356
rect 17316 8372 17368 8424
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 17960 8372 18012 8424
rect 19064 8372 19116 8424
rect 19156 8415 19208 8424
rect 19156 8381 19165 8415
rect 19165 8381 19199 8415
rect 19199 8381 19208 8415
rect 19156 8372 19208 8381
rect 19248 8415 19300 8424
rect 19248 8381 19257 8415
rect 19257 8381 19291 8415
rect 19291 8381 19300 8415
rect 19248 8372 19300 8381
rect 19800 8372 19852 8424
rect 22468 8372 22520 8424
rect 22928 8372 22980 8424
rect 23112 8372 23164 8424
rect 27896 8483 27948 8492
rect 27896 8449 27905 8483
rect 27905 8449 27939 8483
rect 27939 8449 27948 8483
rect 27896 8440 27948 8449
rect 28724 8440 28776 8492
rect 24124 8415 24176 8424
rect 24124 8381 24133 8415
rect 24133 8381 24167 8415
rect 24167 8381 24176 8415
rect 24124 8372 24176 8381
rect 24400 8372 24452 8424
rect 7380 8279 7432 8288
rect 7380 8245 7389 8279
rect 7389 8245 7423 8279
rect 7423 8245 7432 8279
rect 7380 8236 7432 8245
rect 7840 8236 7892 8288
rect 12992 8236 13044 8288
rect 14556 8279 14608 8288
rect 14556 8245 14581 8279
rect 14581 8245 14608 8279
rect 14556 8236 14608 8245
rect 15660 8236 15712 8288
rect 16028 8236 16080 8288
rect 16764 8236 16816 8288
rect 17040 8236 17092 8288
rect 18972 8236 19024 8288
rect 22100 8347 22152 8356
rect 22100 8313 22118 8347
rect 22118 8313 22152 8347
rect 22100 8304 22152 8313
rect 24492 8279 24544 8288
rect 24492 8245 24501 8279
rect 24501 8245 24535 8279
rect 24535 8245 24544 8279
rect 24492 8236 24544 8245
rect 25780 8304 25832 8356
rect 28540 8304 28592 8356
rect 29184 8415 29236 8424
rect 29184 8381 29193 8415
rect 29193 8381 29227 8415
rect 29227 8381 29236 8415
rect 29184 8372 29236 8381
rect 29736 8415 29788 8424
rect 29736 8381 29745 8415
rect 29745 8381 29779 8415
rect 29779 8381 29788 8415
rect 29736 8372 29788 8381
rect 30472 8372 30524 8424
rect 29000 8304 29052 8356
rect 29736 8236 29788 8288
rect 30196 8279 30248 8288
rect 30196 8245 30205 8279
rect 30205 8245 30239 8279
rect 30239 8245 30248 8279
rect 30196 8236 30248 8245
rect 30380 8236 30432 8288
rect 30748 8279 30800 8288
rect 30748 8245 30757 8279
rect 30757 8245 30791 8279
rect 30791 8245 30800 8279
rect 30748 8236 30800 8245
rect 8102 8134 8154 8186
rect 8166 8134 8218 8186
rect 8230 8134 8282 8186
rect 8294 8134 8346 8186
rect 8358 8134 8410 8186
rect 15807 8134 15859 8186
rect 15871 8134 15923 8186
rect 15935 8134 15987 8186
rect 15999 8134 16051 8186
rect 16063 8134 16115 8186
rect 23512 8134 23564 8186
rect 23576 8134 23628 8186
rect 23640 8134 23692 8186
rect 23704 8134 23756 8186
rect 23768 8134 23820 8186
rect 31217 8134 31269 8186
rect 31281 8134 31333 8186
rect 31345 8134 31397 8186
rect 31409 8134 31461 8186
rect 31473 8134 31525 8186
rect 1952 7828 2004 7880
rect 2504 7939 2556 7948
rect 2504 7905 2538 7939
rect 2538 7905 2556 7939
rect 2504 7896 2556 7905
rect 3792 7964 3844 8016
rect 5724 7964 5776 8016
rect 6368 8032 6420 8084
rect 3700 7939 3752 7948
rect 3700 7905 3709 7939
rect 3709 7905 3743 7939
rect 3743 7905 3752 7939
rect 3700 7896 3752 7905
rect 6092 7896 6144 7948
rect 7380 7964 7432 8016
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 8852 8032 8904 8084
rect 12992 8032 13044 8084
rect 10324 7896 10376 7948
rect 12532 7896 12584 7948
rect 13268 8007 13320 8016
rect 13268 7973 13277 8007
rect 13277 7973 13311 8007
rect 13311 7973 13320 8007
rect 13268 7964 13320 7973
rect 13360 7964 13412 8016
rect 13452 8007 13504 8016
rect 13452 7973 13477 8007
rect 13477 7973 13504 8007
rect 13820 8032 13872 8084
rect 15108 8032 15160 8084
rect 15200 8032 15252 8084
rect 13452 7964 13504 7973
rect 15292 7964 15344 8016
rect 16396 8032 16448 8084
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 16764 8032 16816 8084
rect 17040 8032 17092 8084
rect 17684 8032 17736 8084
rect 17868 8032 17920 8084
rect 15568 7896 15620 7948
rect 16396 7896 16448 7948
rect 5724 7828 5776 7880
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 7840 7871 7892 7880
rect 6552 7828 6604 7837
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 8852 7828 8904 7880
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 5632 7692 5684 7744
rect 5724 7692 5776 7744
rect 6276 7692 6328 7744
rect 11244 7692 11296 7744
rect 12624 7692 12676 7744
rect 12808 7735 12860 7744
rect 12808 7701 12817 7735
rect 12817 7701 12851 7735
rect 12851 7701 12860 7735
rect 12808 7692 12860 7701
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 12992 7692 13044 7744
rect 14096 7760 14148 7812
rect 14280 7828 14332 7880
rect 14740 7828 14792 7880
rect 13820 7692 13872 7744
rect 18144 7939 18196 7948
rect 18144 7905 18153 7939
rect 18153 7905 18187 7939
rect 18187 7905 18196 7939
rect 18144 7896 18196 7905
rect 17684 7828 17736 7880
rect 17224 7760 17276 7812
rect 18512 7939 18564 7948
rect 18512 7905 18521 7939
rect 18521 7905 18555 7939
rect 18555 7905 18564 7939
rect 18512 7896 18564 7905
rect 18788 7896 18840 7948
rect 19248 8032 19300 8084
rect 19616 8032 19668 8084
rect 19800 8032 19852 8084
rect 20536 8032 20588 8084
rect 18972 8007 19024 8016
rect 18972 7973 18981 8007
rect 18981 7973 19015 8007
rect 19015 7973 19024 8007
rect 18972 7964 19024 7973
rect 19708 8007 19760 8016
rect 19708 7973 19717 8007
rect 19717 7973 19751 8007
rect 19751 7973 19760 8007
rect 19708 7964 19760 7973
rect 19248 7828 19300 7880
rect 19984 7828 20036 7880
rect 18696 7692 18748 7744
rect 18788 7735 18840 7744
rect 18788 7701 18797 7735
rect 18797 7701 18831 7735
rect 18831 7701 18840 7735
rect 21640 8032 21692 8084
rect 21732 8032 21784 8084
rect 22100 8032 22152 8084
rect 22560 8075 22612 8084
rect 22560 8041 22569 8075
rect 22569 8041 22603 8075
rect 22603 8041 22612 8075
rect 22560 8032 22612 8041
rect 24492 8032 24544 8084
rect 27896 8032 27948 8084
rect 28540 8032 28592 8084
rect 30288 8032 30340 8084
rect 30932 8075 30984 8084
rect 30932 8041 30941 8075
rect 30941 8041 30975 8075
rect 30975 8041 30984 8075
rect 30932 8032 30984 8041
rect 21824 7964 21876 8016
rect 22192 7896 22244 7948
rect 22652 7896 22704 7948
rect 25964 7896 26016 7948
rect 27804 7939 27856 7948
rect 27804 7905 27822 7939
rect 27822 7905 27856 7939
rect 27804 7896 27856 7905
rect 30196 7964 30248 8016
rect 30564 7964 30616 8016
rect 21272 7760 21324 7812
rect 22928 7828 22980 7880
rect 25412 7871 25464 7880
rect 25412 7837 25421 7871
rect 25421 7837 25455 7871
rect 25455 7837 25464 7871
rect 25412 7828 25464 7837
rect 18788 7692 18840 7701
rect 20168 7692 20220 7744
rect 21640 7692 21692 7744
rect 22284 7692 22336 7744
rect 26700 7803 26752 7812
rect 26700 7769 26709 7803
rect 26709 7769 26743 7803
rect 26743 7769 26752 7803
rect 26700 7760 26752 7769
rect 28448 7760 28500 7812
rect 29000 7896 29052 7948
rect 29368 7896 29420 7948
rect 24676 7692 24728 7744
rect 28632 7735 28684 7744
rect 28632 7701 28641 7735
rect 28641 7701 28675 7735
rect 28675 7701 28684 7735
rect 28632 7692 28684 7701
rect 29184 7735 29236 7744
rect 29184 7701 29193 7735
rect 29193 7701 29227 7735
rect 29227 7701 29236 7735
rect 29184 7692 29236 7701
rect 30748 7760 30800 7812
rect 4250 7590 4302 7642
rect 4314 7590 4366 7642
rect 4378 7590 4430 7642
rect 4442 7590 4494 7642
rect 4506 7590 4558 7642
rect 11955 7590 12007 7642
rect 12019 7590 12071 7642
rect 12083 7590 12135 7642
rect 12147 7590 12199 7642
rect 12211 7590 12263 7642
rect 19660 7590 19712 7642
rect 19724 7590 19776 7642
rect 19788 7590 19840 7642
rect 19852 7590 19904 7642
rect 19916 7590 19968 7642
rect 27365 7590 27417 7642
rect 27429 7590 27481 7642
rect 27493 7590 27545 7642
rect 27557 7590 27609 7642
rect 27621 7590 27673 7642
rect 6184 7420 6236 7472
rect 6552 7352 6604 7404
rect 1952 7284 2004 7336
rect 5724 7284 5776 7336
rect 6000 7327 6052 7336
rect 6000 7293 6009 7327
rect 6009 7293 6043 7327
rect 6043 7293 6052 7327
rect 6000 7284 6052 7293
rect 6092 7327 6144 7336
rect 6092 7293 6101 7327
rect 6101 7293 6135 7327
rect 6135 7293 6144 7327
rect 6092 7284 6144 7293
rect 6276 7284 6328 7336
rect 6460 7327 6512 7336
rect 6460 7293 6469 7327
rect 6469 7293 6503 7327
rect 6503 7293 6512 7327
rect 6460 7284 6512 7293
rect 8024 7420 8076 7472
rect 11520 7488 11572 7540
rect 12900 7488 12952 7540
rect 12992 7488 13044 7540
rect 13912 7488 13964 7540
rect 14740 7488 14792 7540
rect 15568 7488 15620 7540
rect 16212 7488 16264 7540
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 8760 7352 8812 7404
rect 1400 7259 1452 7268
rect 1400 7225 1434 7259
rect 1434 7225 1452 7259
rect 1400 7216 1452 7225
rect 5632 7216 5684 7268
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 7196 7216 7248 7268
rect 8024 7216 8076 7268
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 8668 7148 8720 7200
rect 12440 7284 12492 7336
rect 10968 7216 11020 7268
rect 11244 7216 11296 7268
rect 13452 7284 13504 7336
rect 15200 7420 15252 7472
rect 16304 7420 16356 7472
rect 16396 7420 16448 7472
rect 18328 7420 18380 7472
rect 14556 7352 14608 7404
rect 21456 7488 21508 7540
rect 21732 7488 21784 7540
rect 21824 7488 21876 7540
rect 22192 7531 22244 7540
rect 22192 7497 22201 7531
rect 22201 7497 22235 7531
rect 22235 7497 22244 7531
rect 22192 7488 22244 7497
rect 21272 7420 21324 7472
rect 27804 7488 27856 7540
rect 30288 7531 30340 7540
rect 30288 7497 30297 7531
rect 30297 7497 30331 7531
rect 30331 7497 30340 7531
rect 30288 7488 30340 7497
rect 30748 7488 30800 7540
rect 24676 7463 24728 7472
rect 24676 7429 24685 7463
rect 24685 7429 24719 7463
rect 24719 7429 24728 7463
rect 24676 7420 24728 7429
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 11612 7191 11664 7200
rect 11612 7157 11637 7191
rect 11637 7157 11664 7191
rect 11612 7148 11664 7157
rect 12716 7148 12768 7200
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 16488 7284 16540 7336
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 17224 7327 17276 7336
rect 17224 7293 17233 7327
rect 17233 7293 17267 7327
rect 17267 7293 17276 7327
rect 17224 7284 17276 7293
rect 17316 7327 17368 7336
rect 17316 7293 17325 7327
rect 17325 7293 17359 7327
rect 17359 7293 17368 7327
rect 17316 7284 17368 7293
rect 17684 7284 17736 7336
rect 21916 7352 21968 7404
rect 21180 7329 21232 7336
rect 21180 7295 21189 7329
rect 21189 7295 21223 7329
rect 21223 7295 21232 7329
rect 21180 7284 21232 7295
rect 21456 7327 21508 7336
rect 21456 7293 21465 7327
rect 21465 7293 21499 7327
rect 21499 7293 21508 7327
rect 21456 7284 21508 7293
rect 21548 7327 21600 7336
rect 21548 7293 21557 7327
rect 21557 7293 21591 7327
rect 21591 7293 21600 7327
rect 21548 7284 21600 7293
rect 21824 7284 21876 7336
rect 22376 7327 22428 7336
rect 22376 7293 22385 7327
rect 22385 7293 22419 7327
rect 22419 7293 22428 7327
rect 22376 7284 22428 7293
rect 25964 7284 26016 7336
rect 27896 7352 27948 7404
rect 28908 7352 28960 7404
rect 28448 7284 28500 7336
rect 22928 7259 22980 7268
rect 22928 7225 22937 7259
rect 22937 7225 22971 7259
rect 22971 7225 22980 7259
rect 22928 7216 22980 7225
rect 27528 7216 27580 7268
rect 29736 7284 29788 7336
rect 30472 7327 30524 7336
rect 30472 7293 30473 7327
rect 30473 7293 30507 7327
rect 30507 7293 30524 7327
rect 30472 7284 30524 7293
rect 30564 7327 30616 7336
rect 30564 7293 30573 7327
rect 30573 7293 30607 7327
rect 30607 7293 30616 7327
rect 30564 7284 30616 7293
rect 30748 7216 30800 7268
rect 19248 7148 19300 7200
rect 20812 7148 20864 7200
rect 21548 7148 21600 7200
rect 23204 7148 23256 7200
rect 24400 7148 24452 7200
rect 26056 7148 26108 7200
rect 28540 7148 28592 7200
rect 29276 7191 29328 7200
rect 29276 7157 29285 7191
rect 29285 7157 29319 7191
rect 29319 7157 29328 7191
rect 29276 7148 29328 7157
rect 29828 7148 29880 7200
rect 30656 7191 30708 7200
rect 30656 7157 30665 7191
rect 30665 7157 30699 7191
rect 30699 7157 30708 7191
rect 30656 7148 30708 7157
rect 8102 7046 8154 7098
rect 8166 7046 8218 7098
rect 8230 7046 8282 7098
rect 8294 7046 8346 7098
rect 8358 7046 8410 7098
rect 15807 7046 15859 7098
rect 15871 7046 15923 7098
rect 15935 7046 15987 7098
rect 15999 7046 16051 7098
rect 16063 7046 16115 7098
rect 23512 7046 23564 7098
rect 23576 7046 23628 7098
rect 23640 7046 23692 7098
rect 23704 7046 23756 7098
rect 23768 7046 23820 7098
rect 31217 7046 31269 7098
rect 31281 7046 31333 7098
rect 31345 7046 31397 7098
rect 31409 7046 31461 7098
rect 31473 7046 31525 7098
rect 5540 6944 5592 6996
rect 5632 6876 5684 6928
rect 1952 6808 2004 6860
rect 2228 6808 2280 6860
rect 6552 6876 6604 6928
rect 7196 6876 7248 6928
rect 7288 6919 7340 6928
rect 7288 6885 7297 6919
rect 7297 6885 7331 6919
rect 7331 6885 7340 6919
rect 7288 6876 7340 6885
rect 8024 6876 8076 6928
rect 8668 6987 8720 6996
rect 8668 6953 8677 6987
rect 8677 6953 8711 6987
rect 8711 6953 8720 6987
rect 8668 6944 8720 6953
rect 12532 6919 12584 6928
rect 12532 6885 12541 6919
rect 12541 6885 12575 6919
rect 12575 6885 12584 6919
rect 12532 6876 12584 6885
rect 13452 6944 13504 6996
rect 13912 6944 13964 6996
rect 14648 6944 14700 6996
rect 15292 6944 15344 6996
rect 13268 6876 13320 6928
rect 14280 6876 14332 6928
rect 15660 6876 15712 6928
rect 16488 6944 16540 6996
rect 16764 6944 16816 6996
rect 17224 6944 17276 6996
rect 6184 6808 6236 6860
rect 17132 6876 17184 6928
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 6920 6740 6972 6792
rect 7748 6808 7800 6860
rect 8668 6808 8720 6860
rect 10508 6808 10560 6860
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 3608 6604 3660 6656
rect 8852 6672 8904 6724
rect 8484 6604 8536 6656
rect 8944 6604 8996 6656
rect 10324 6604 10376 6656
rect 10968 6783 11020 6792
rect 10968 6749 10977 6783
rect 10977 6749 11011 6783
rect 11011 6749 11020 6783
rect 10968 6740 11020 6749
rect 12256 6672 12308 6724
rect 13820 6851 13872 6860
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 14004 6808 14056 6860
rect 14740 6808 14792 6860
rect 15292 6851 15344 6860
rect 15292 6817 15301 6851
rect 15301 6817 15335 6851
rect 15335 6817 15344 6851
rect 15292 6808 15344 6817
rect 12716 6740 12768 6792
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 12716 6647 12768 6656
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 14832 6740 14884 6792
rect 15936 6808 15988 6860
rect 16120 6808 16172 6860
rect 17316 6876 17368 6928
rect 18328 6944 18380 6996
rect 17500 6808 17552 6860
rect 17776 6808 17828 6860
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 20536 6944 20588 6996
rect 21548 6944 21600 6996
rect 27528 6987 27580 6996
rect 27528 6953 27537 6987
rect 27537 6953 27571 6987
rect 27571 6953 27580 6987
rect 27528 6944 27580 6953
rect 27712 6944 27764 6996
rect 27896 6944 27948 6996
rect 29184 6944 29236 6996
rect 30564 6944 30616 6996
rect 30656 6944 30708 6996
rect 19708 6919 19760 6928
rect 19708 6885 19717 6919
rect 19717 6885 19751 6919
rect 19751 6885 19760 6919
rect 19708 6876 19760 6885
rect 23848 6876 23900 6928
rect 24400 6876 24452 6928
rect 25964 6876 26016 6928
rect 28632 6876 28684 6928
rect 14556 6672 14608 6724
rect 12716 6604 12768 6613
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 13360 6604 13412 6613
rect 13452 6647 13504 6656
rect 13452 6613 13461 6647
rect 13461 6613 13495 6647
rect 13495 6613 13504 6647
rect 13452 6604 13504 6613
rect 14188 6604 14240 6656
rect 15108 6647 15160 6656
rect 15108 6613 15117 6647
rect 15117 6613 15151 6647
rect 15151 6613 15160 6647
rect 15108 6604 15160 6613
rect 16764 6740 16816 6792
rect 18880 6783 18932 6792
rect 18880 6749 18889 6783
rect 18889 6749 18923 6783
rect 18923 6749 18932 6783
rect 18880 6740 18932 6749
rect 16304 6604 16356 6656
rect 16764 6647 16816 6656
rect 16764 6613 16773 6647
rect 16773 6613 16807 6647
rect 16807 6613 16816 6647
rect 16764 6604 16816 6613
rect 21456 6740 21508 6792
rect 22284 6851 22336 6860
rect 22284 6817 22293 6851
rect 22293 6817 22327 6851
rect 22327 6817 22336 6851
rect 22284 6808 22336 6817
rect 17684 6604 17736 6656
rect 19064 6672 19116 6724
rect 17868 6604 17920 6656
rect 17960 6604 18012 6656
rect 20168 6672 20220 6724
rect 21180 6672 21232 6724
rect 22100 6740 22152 6792
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 22376 6672 22428 6724
rect 23940 6851 23992 6860
rect 23940 6817 23958 6851
rect 23958 6817 23992 6851
rect 23940 6808 23992 6817
rect 26240 6851 26292 6860
rect 26240 6817 26249 6851
rect 26249 6817 26283 6851
rect 26283 6817 26292 6851
rect 26240 6808 26292 6817
rect 27804 6808 27856 6860
rect 28724 6851 28776 6860
rect 28724 6817 28733 6851
rect 28733 6817 28767 6851
rect 28767 6817 28776 6851
rect 28724 6808 28776 6817
rect 28908 6808 28960 6860
rect 29736 6851 29788 6860
rect 29736 6817 29745 6851
rect 29745 6817 29779 6851
rect 29779 6817 29788 6851
rect 29736 6808 29788 6817
rect 29828 6851 29880 6860
rect 29828 6817 29837 6851
rect 29837 6817 29871 6851
rect 29871 6817 29880 6851
rect 29828 6808 29880 6817
rect 22652 6604 22704 6656
rect 22836 6647 22888 6656
rect 22836 6613 22845 6647
rect 22845 6613 22879 6647
rect 22879 6613 22888 6647
rect 22836 6604 22888 6613
rect 22928 6604 22980 6656
rect 27160 6604 27212 6656
rect 28172 6647 28224 6656
rect 28172 6613 28181 6647
rect 28181 6613 28215 6647
rect 28215 6613 28224 6647
rect 28172 6604 28224 6613
rect 28816 6647 28868 6656
rect 28816 6613 28825 6647
rect 28825 6613 28859 6647
rect 28859 6613 28868 6647
rect 28816 6604 28868 6613
rect 29736 6604 29788 6656
rect 30656 6647 30708 6656
rect 30656 6613 30665 6647
rect 30665 6613 30699 6647
rect 30699 6613 30708 6647
rect 30656 6604 30708 6613
rect 30932 6604 30984 6656
rect 4250 6502 4302 6554
rect 4314 6502 4366 6554
rect 4378 6502 4430 6554
rect 4442 6502 4494 6554
rect 4506 6502 4558 6554
rect 11955 6502 12007 6554
rect 12019 6502 12071 6554
rect 12083 6502 12135 6554
rect 12147 6502 12199 6554
rect 12211 6502 12263 6554
rect 19660 6502 19712 6554
rect 19724 6502 19776 6554
rect 19788 6502 19840 6554
rect 19852 6502 19904 6554
rect 19916 6502 19968 6554
rect 27365 6502 27417 6554
rect 27429 6502 27481 6554
rect 27493 6502 27545 6554
rect 27557 6502 27609 6554
rect 27621 6502 27673 6554
rect 6000 6400 6052 6452
rect 1032 6196 1084 6248
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 2596 6196 2648 6205
rect 2964 6264 3016 6316
rect 6276 6400 6328 6452
rect 8484 6443 8536 6452
rect 8484 6409 8493 6443
rect 8493 6409 8527 6443
rect 8527 6409 8536 6443
rect 8484 6400 8536 6409
rect 9772 6400 9824 6452
rect 10508 6443 10560 6452
rect 10508 6409 10517 6443
rect 10517 6409 10551 6443
rect 10551 6409 10560 6443
rect 10508 6400 10560 6409
rect 12716 6400 12768 6452
rect 13360 6400 13412 6452
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 14372 6400 14424 6452
rect 14464 6400 14516 6452
rect 14832 6400 14884 6452
rect 15292 6400 15344 6452
rect 3056 6196 3108 6248
rect 3608 6196 3660 6248
rect 4436 6239 4488 6248
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 5080 6196 5132 6248
rect 8760 6264 8812 6316
rect 10600 6264 10652 6316
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 4896 6128 4948 6180
rect 6552 6196 6604 6248
rect 8852 6196 8904 6248
rect 8944 6239 8996 6248
rect 8944 6205 8953 6239
rect 8953 6205 8987 6239
rect 8987 6205 8996 6239
rect 8944 6196 8996 6205
rect 9680 6128 9732 6180
rect 2412 6060 2464 6112
rect 3148 6060 3200 6112
rect 4160 6060 4212 6112
rect 8944 6060 8996 6112
rect 9036 6103 9088 6112
rect 9036 6069 9045 6103
rect 9045 6069 9079 6103
rect 9079 6069 9088 6103
rect 9036 6060 9088 6069
rect 10324 6196 10376 6248
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 10692 6239 10744 6248
rect 10692 6205 10701 6239
rect 10701 6205 10735 6239
rect 10735 6205 10744 6239
rect 10692 6196 10744 6205
rect 11612 6196 11664 6248
rect 10324 6060 10376 6112
rect 12716 6171 12768 6180
rect 12716 6137 12725 6171
rect 12725 6137 12759 6171
rect 12759 6137 12768 6171
rect 12716 6128 12768 6137
rect 13360 6196 13412 6248
rect 15936 6375 15988 6384
rect 15936 6341 15945 6375
rect 15945 6341 15979 6375
rect 15979 6341 15988 6375
rect 15936 6332 15988 6341
rect 16120 6332 16172 6384
rect 16856 6332 16908 6384
rect 21456 6400 21508 6452
rect 22100 6443 22152 6452
rect 22100 6409 22109 6443
rect 22109 6409 22143 6443
rect 22143 6409 22152 6443
rect 22100 6400 22152 6409
rect 22284 6400 22336 6452
rect 13820 6239 13872 6248
rect 13820 6205 13829 6239
rect 13829 6205 13863 6239
rect 13863 6205 13872 6239
rect 13820 6196 13872 6205
rect 13912 6239 13964 6248
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 14924 6196 14976 6248
rect 15200 6196 15252 6248
rect 15568 6239 15620 6248
rect 15568 6205 15593 6239
rect 15593 6205 15620 6239
rect 15568 6196 15620 6205
rect 17868 6264 17920 6316
rect 18788 6264 18840 6316
rect 19340 6264 19392 6316
rect 13636 6060 13688 6112
rect 14372 6171 14424 6180
rect 14372 6137 14381 6171
rect 14381 6137 14415 6171
rect 14415 6137 14424 6171
rect 14372 6128 14424 6137
rect 18512 6196 18564 6248
rect 18880 6239 18932 6248
rect 18880 6205 18889 6239
rect 18889 6205 18923 6239
rect 18923 6205 18932 6239
rect 18880 6196 18932 6205
rect 20168 6196 20220 6248
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 21364 6196 21416 6248
rect 21916 6239 21968 6248
rect 21916 6205 21925 6239
rect 21925 6205 21959 6239
rect 21959 6205 21968 6239
rect 21916 6196 21968 6205
rect 22652 6375 22704 6384
rect 22652 6341 22661 6375
rect 22661 6341 22695 6375
rect 22695 6341 22704 6375
rect 22652 6332 22704 6341
rect 24216 6443 24268 6452
rect 24216 6409 24225 6443
rect 24225 6409 24259 6443
rect 24259 6409 24268 6443
rect 24216 6400 24268 6409
rect 28632 6400 28684 6452
rect 31024 6443 31076 6452
rect 31024 6409 31033 6443
rect 31033 6409 31067 6443
rect 31067 6409 31076 6443
rect 31024 6400 31076 6409
rect 26240 6332 26292 6384
rect 28816 6332 28868 6384
rect 23940 6264 23992 6316
rect 16856 6128 16908 6180
rect 17500 6128 17552 6180
rect 17776 6128 17828 6180
rect 21180 6171 21232 6180
rect 21180 6137 21189 6171
rect 21189 6137 21223 6171
rect 21223 6137 21232 6171
rect 21180 6128 21232 6137
rect 18144 6060 18196 6112
rect 19524 6060 19576 6112
rect 23756 6196 23808 6248
rect 24216 6196 24268 6248
rect 22376 6103 22428 6112
rect 22376 6069 22385 6103
rect 22385 6069 22419 6103
rect 22419 6069 22428 6103
rect 22376 6060 22428 6069
rect 22652 6060 22704 6112
rect 24492 6060 24544 6112
rect 25136 6196 25188 6248
rect 25780 6196 25832 6248
rect 26056 6196 26108 6248
rect 26332 6239 26384 6248
rect 26332 6205 26341 6239
rect 26341 6205 26375 6239
rect 26375 6205 26384 6239
rect 26332 6196 26384 6205
rect 27160 6196 27212 6248
rect 27436 6196 27488 6248
rect 27620 6239 27672 6248
rect 27620 6205 27629 6239
rect 27629 6205 27663 6239
rect 27663 6205 27672 6239
rect 27620 6196 27672 6205
rect 28172 6239 28224 6248
rect 28172 6205 28181 6239
rect 28181 6205 28215 6239
rect 28215 6205 28224 6239
rect 28540 6264 28592 6316
rect 29184 6264 29236 6316
rect 28448 6241 28500 6248
rect 28172 6196 28224 6205
rect 28448 6207 28457 6241
rect 28457 6207 28491 6241
rect 28491 6207 28500 6241
rect 28448 6196 28500 6207
rect 29644 6239 29696 6248
rect 29644 6205 29653 6239
rect 29653 6205 29687 6239
rect 29687 6205 29696 6239
rect 29644 6196 29696 6205
rect 29736 6196 29788 6248
rect 30380 6196 30432 6248
rect 27436 6060 27488 6112
rect 29368 6103 29420 6112
rect 29368 6069 29377 6103
rect 29377 6069 29411 6103
rect 29411 6069 29420 6103
rect 29368 6060 29420 6069
rect 8102 5958 8154 6010
rect 8166 5958 8218 6010
rect 8230 5958 8282 6010
rect 8294 5958 8346 6010
rect 8358 5958 8410 6010
rect 15807 5958 15859 6010
rect 15871 5958 15923 6010
rect 15935 5958 15987 6010
rect 15999 5958 16051 6010
rect 16063 5958 16115 6010
rect 23512 5958 23564 6010
rect 23576 5958 23628 6010
rect 23640 5958 23692 6010
rect 23704 5958 23756 6010
rect 23768 5958 23820 6010
rect 31217 5958 31269 6010
rect 31281 5958 31333 6010
rect 31345 5958 31397 6010
rect 31409 5958 31461 6010
rect 31473 5958 31525 6010
rect 2596 5856 2648 5908
rect 2688 5788 2740 5840
rect 4436 5856 4488 5908
rect 4620 5899 4672 5908
rect 4620 5865 4629 5899
rect 4629 5865 4663 5899
rect 4663 5865 4672 5899
rect 4620 5856 4672 5865
rect 4896 5899 4948 5908
rect 4896 5865 4905 5899
rect 4905 5865 4939 5899
rect 4939 5865 4948 5899
rect 4896 5856 4948 5865
rect 1400 5763 1452 5772
rect 1400 5729 1423 5763
rect 1423 5729 1452 5763
rect 1400 5720 1452 5729
rect 2964 5720 3016 5772
rect 3148 5763 3200 5772
rect 3148 5729 3157 5763
rect 3157 5729 3191 5763
rect 3191 5729 3200 5763
rect 3148 5720 3200 5729
rect 4160 5788 4212 5840
rect 8944 5856 8996 5908
rect 9588 5856 9640 5908
rect 10324 5899 10376 5908
rect 10324 5865 10333 5899
rect 10333 5865 10367 5899
rect 10367 5865 10376 5899
rect 10324 5856 10376 5865
rect 11612 5788 11664 5840
rect 12348 5856 12400 5908
rect 12716 5856 12768 5908
rect 14280 5856 14332 5908
rect 15108 5856 15160 5908
rect 3516 5763 3568 5772
rect 3516 5729 3550 5763
rect 3550 5729 3568 5763
rect 3516 5720 3568 5729
rect 4988 5763 5040 5772
rect 4988 5729 4997 5763
rect 4997 5729 5031 5763
rect 5031 5729 5040 5763
rect 4988 5720 5040 5729
rect 5080 5720 5132 5772
rect 5448 5720 5500 5772
rect 5724 5720 5776 5772
rect 7748 5720 7800 5772
rect 8208 5720 8260 5772
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 9956 5763 10008 5772
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 9956 5720 10008 5729
rect 10416 5763 10468 5772
rect 10416 5729 10425 5763
rect 10425 5729 10459 5763
rect 10459 5729 10468 5763
rect 10416 5720 10468 5729
rect 14096 5831 14148 5840
rect 14096 5797 14105 5831
rect 14105 5797 14139 5831
rect 14139 5797 14148 5831
rect 14096 5788 14148 5797
rect 19984 5856 20036 5908
rect 19248 5831 19300 5840
rect 12256 5720 12308 5772
rect 14924 5763 14976 5772
rect 14924 5729 14933 5763
rect 14933 5729 14967 5763
rect 14967 5729 14976 5763
rect 14924 5720 14976 5729
rect 15568 5720 15620 5772
rect 16488 5763 16540 5772
rect 2412 5584 2464 5636
rect 10692 5652 10744 5704
rect 16488 5729 16497 5763
rect 16497 5729 16531 5763
rect 16531 5729 16540 5763
rect 16488 5720 16540 5729
rect 16856 5763 16908 5772
rect 16856 5729 16865 5763
rect 16865 5729 16899 5763
rect 16899 5729 16908 5763
rect 16856 5720 16908 5729
rect 16948 5720 17000 5772
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 9496 5584 9548 5636
rect 7288 5516 7340 5568
rect 9036 5516 9088 5568
rect 9312 5516 9364 5568
rect 17316 5720 17368 5772
rect 18880 5720 18932 5772
rect 19248 5797 19275 5831
rect 19275 5797 19300 5831
rect 19248 5788 19300 5797
rect 19800 5788 19852 5840
rect 19892 5831 19944 5840
rect 19892 5797 19901 5831
rect 19901 5797 19935 5831
rect 19935 5797 19944 5831
rect 19892 5788 19944 5797
rect 23572 5856 23624 5908
rect 24492 5856 24544 5908
rect 25320 5856 25372 5908
rect 26332 5856 26384 5908
rect 27804 5856 27856 5908
rect 28448 5856 28500 5908
rect 29184 5856 29236 5908
rect 30564 5856 30616 5908
rect 17500 5652 17552 5704
rect 21456 5788 21508 5840
rect 21364 5720 21416 5772
rect 21548 5763 21600 5772
rect 21548 5729 21582 5763
rect 21582 5729 21600 5763
rect 21548 5720 21600 5729
rect 21732 5788 21784 5840
rect 22376 5788 22428 5840
rect 23204 5788 23256 5840
rect 12440 5516 12492 5568
rect 12900 5516 12952 5568
rect 13268 5516 13320 5568
rect 17500 5516 17552 5568
rect 17868 5559 17920 5568
rect 17868 5525 17877 5559
rect 17877 5525 17911 5559
rect 17911 5525 17920 5559
rect 17868 5516 17920 5525
rect 18512 5584 18564 5636
rect 18788 5516 18840 5568
rect 19064 5516 19116 5568
rect 19616 5584 19668 5636
rect 19984 5559 20036 5568
rect 19984 5525 19993 5559
rect 19993 5525 20027 5559
rect 20027 5525 20036 5559
rect 19984 5516 20036 5525
rect 20444 5559 20496 5568
rect 20444 5525 20453 5559
rect 20453 5525 20487 5559
rect 20487 5525 20496 5559
rect 20444 5516 20496 5525
rect 23020 5695 23072 5704
rect 23020 5661 23029 5695
rect 23029 5661 23063 5695
rect 23063 5661 23072 5695
rect 23020 5652 23072 5661
rect 23296 5763 23348 5772
rect 23296 5729 23305 5763
rect 23305 5729 23339 5763
rect 23339 5729 23348 5763
rect 23296 5720 23348 5729
rect 23940 5720 23992 5772
rect 25136 5788 25188 5840
rect 26056 5788 26108 5840
rect 26240 5788 26292 5840
rect 23480 5652 23532 5704
rect 24308 5652 24360 5704
rect 24952 5652 25004 5704
rect 27988 5788 28040 5840
rect 25320 5652 25372 5704
rect 27160 5720 27212 5772
rect 29644 5788 29696 5840
rect 28540 5720 28592 5772
rect 29092 5720 29144 5772
rect 29184 5763 29236 5772
rect 29184 5729 29193 5763
rect 29193 5729 29227 5763
rect 29227 5729 29236 5763
rect 29184 5720 29236 5729
rect 29368 5720 29420 5772
rect 30656 5720 30708 5772
rect 30748 5763 30800 5772
rect 30748 5729 30757 5763
rect 30757 5729 30791 5763
rect 30791 5729 30800 5763
rect 30748 5720 30800 5729
rect 30932 5899 30984 5908
rect 30932 5865 30941 5899
rect 30941 5865 30975 5899
rect 30975 5865 30984 5899
rect 30932 5856 30984 5865
rect 22652 5559 22704 5568
rect 22652 5525 22661 5559
rect 22661 5525 22695 5559
rect 22695 5525 22704 5559
rect 22652 5516 22704 5525
rect 22836 5584 22888 5636
rect 22928 5584 22980 5636
rect 29368 5627 29420 5636
rect 29368 5593 29377 5627
rect 29377 5593 29411 5627
rect 29411 5593 29420 5627
rect 29368 5584 29420 5593
rect 25044 5516 25096 5568
rect 4250 5414 4302 5466
rect 4314 5414 4366 5466
rect 4378 5414 4430 5466
rect 4442 5414 4494 5466
rect 4506 5414 4558 5466
rect 11955 5414 12007 5466
rect 12019 5414 12071 5466
rect 12083 5414 12135 5466
rect 12147 5414 12199 5466
rect 12211 5414 12263 5466
rect 19660 5414 19712 5466
rect 19724 5414 19776 5466
rect 19788 5414 19840 5466
rect 19852 5414 19904 5466
rect 19916 5414 19968 5466
rect 27365 5414 27417 5466
rect 27429 5414 27481 5466
rect 27493 5414 27545 5466
rect 27557 5414 27609 5466
rect 27621 5414 27673 5466
rect 2228 5312 2280 5364
rect 2412 5312 2464 5364
rect 2596 5312 2648 5364
rect 4988 5312 5040 5364
rect 1676 5151 1728 5160
rect 1676 5117 1685 5151
rect 1685 5117 1719 5151
rect 1719 5117 1728 5151
rect 1676 5108 1728 5117
rect 1952 5108 2004 5160
rect 4896 5244 4948 5296
rect 5080 5287 5132 5296
rect 5080 5253 5089 5287
rect 5089 5253 5123 5287
rect 5123 5253 5132 5287
rect 5080 5244 5132 5253
rect 3148 5108 3200 5160
rect 4160 5108 4212 5160
rect 5448 5312 5500 5364
rect 9220 5312 9272 5364
rect 9956 5312 10008 5364
rect 3516 5040 3568 5092
rect 7748 5244 7800 5296
rect 8208 5244 8260 5296
rect 9496 5244 9548 5296
rect 7288 5108 7340 5160
rect 1400 4972 1452 5024
rect 5080 4972 5132 5024
rect 9312 5151 9364 5160
rect 9312 5117 9321 5151
rect 9321 5117 9355 5151
rect 9355 5117 9364 5151
rect 9312 5108 9364 5117
rect 9772 5151 9824 5160
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 9772 5108 9824 5117
rect 10324 5312 10376 5364
rect 10416 5312 10468 5364
rect 12348 5312 12400 5364
rect 14096 5312 14148 5364
rect 15384 5312 15436 5364
rect 15936 5355 15988 5364
rect 15936 5321 15945 5355
rect 15945 5321 15979 5355
rect 15979 5321 15988 5355
rect 15936 5312 15988 5321
rect 16304 5312 16356 5364
rect 13084 5244 13136 5296
rect 10600 5219 10652 5228
rect 10600 5185 10609 5219
rect 10609 5185 10643 5219
rect 10643 5185 10652 5219
rect 10600 5176 10652 5185
rect 15568 5244 15620 5296
rect 16488 5244 16540 5296
rect 18788 5312 18840 5364
rect 19524 5312 19576 5364
rect 19984 5312 20036 5364
rect 20260 5355 20312 5364
rect 20260 5321 20269 5355
rect 20269 5321 20303 5355
rect 20303 5321 20312 5355
rect 20260 5312 20312 5321
rect 20444 5312 20496 5364
rect 20720 5355 20772 5364
rect 20720 5321 20729 5355
rect 20729 5321 20763 5355
rect 20763 5321 20772 5355
rect 20720 5312 20772 5321
rect 20812 5312 20864 5364
rect 13452 5108 13504 5160
rect 15384 5108 15436 5160
rect 7380 4972 7432 5024
rect 7748 4972 7800 5024
rect 10416 4972 10468 5024
rect 12164 5040 12216 5092
rect 12992 5083 13044 5092
rect 12992 5049 13001 5083
rect 13001 5049 13035 5083
rect 13035 5049 13044 5083
rect 12992 5040 13044 5049
rect 11244 4972 11296 5024
rect 15016 5083 15068 5092
rect 15016 5049 15025 5083
rect 15025 5049 15059 5083
rect 15059 5049 15068 5083
rect 15016 5040 15068 5049
rect 15660 5108 15712 5160
rect 16212 5108 16264 5160
rect 18420 5176 18472 5228
rect 19524 5176 19576 5228
rect 17500 5151 17552 5160
rect 17500 5117 17509 5151
rect 17509 5117 17543 5151
rect 17543 5117 17552 5151
rect 17500 5108 17552 5117
rect 14740 4972 14792 5024
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 15476 4972 15528 4981
rect 16396 5040 16448 5092
rect 16856 5040 16908 5092
rect 16580 4972 16632 5024
rect 16948 4972 17000 5024
rect 19156 5108 19208 5160
rect 18880 5083 18932 5092
rect 18880 5049 18907 5083
rect 18907 5049 18932 5083
rect 18880 5040 18932 5049
rect 19984 5151 20036 5160
rect 19984 5117 19993 5151
rect 19993 5117 20027 5151
rect 20027 5117 20036 5151
rect 19984 5108 20036 5117
rect 20996 5244 21048 5296
rect 22928 5244 22980 5296
rect 23112 5244 23164 5296
rect 23572 5312 23624 5364
rect 24860 5312 24912 5364
rect 25044 5312 25096 5364
rect 28724 5355 28776 5364
rect 28724 5321 28733 5355
rect 28733 5321 28767 5355
rect 28767 5321 28776 5355
rect 28724 5312 28776 5321
rect 28908 5244 28960 5296
rect 30380 5244 30432 5296
rect 20628 5176 20680 5228
rect 22652 5176 22704 5228
rect 25412 5176 25464 5228
rect 20260 5108 20312 5160
rect 20996 5151 21048 5160
rect 20996 5117 21005 5151
rect 21005 5117 21039 5151
rect 21039 5117 21048 5151
rect 20996 5108 21048 5117
rect 21640 5108 21692 5160
rect 23112 5108 23164 5160
rect 24952 5151 25004 5160
rect 24952 5117 24970 5151
rect 24970 5117 25004 5151
rect 24952 5108 25004 5117
rect 27160 5108 27212 5160
rect 27988 5108 28040 5160
rect 28632 5108 28684 5160
rect 28908 5108 28960 5160
rect 29276 5151 29328 5160
rect 29276 5117 29310 5151
rect 29310 5117 29328 5151
rect 29276 5108 29328 5117
rect 30564 5355 30616 5364
rect 30564 5321 30573 5355
rect 30573 5321 30607 5355
rect 30607 5321 30616 5355
rect 30564 5312 30616 5321
rect 18696 5015 18748 5024
rect 18696 4981 18705 5015
rect 18705 4981 18739 5015
rect 18739 4981 18748 5015
rect 18696 4972 18748 4981
rect 20812 4972 20864 5024
rect 22836 5083 22888 5092
rect 22836 5049 22845 5083
rect 22845 5049 22879 5083
rect 22879 5049 22888 5083
rect 22836 5040 22888 5049
rect 23848 5040 23900 5092
rect 24860 5040 24912 5092
rect 23112 4972 23164 5024
rect 23204 4972 23256 5024
rect 23480 4972 23532 5024
rect 8102 4870 8154 4922
rect 8166 4870 8218 4922
rect 8230 4870 8282 4922
rect 8294 4870 8346 4922
rect 8358 4870 8410 4922
rect 15807 4870 15859 4922
rect 15871 4870 15923 4922
rect 15935 4870 15987 4922
rect 15999 4870 16051 4922
rect 16063 4870 16115 4922
rect 23512 4870 23564 4922
rect 23576 4870 23628 4922
rect 23640 4870 23692 4922
rect 23704 4870 23756 4922
rect 23768 4870 23820 4922
rect 31217 4870 31269 4922
rect 31281 4870 31333 4922
rect 31345 4870 31397 4922
rect 31409 4870 31461 4922
rect 31473 4870 31525 4922
rect 1400 4768 1452 4820
rect 1676 4768 1728 4820
rect 1952 4768 2004 4820
rect 3056 4768 3108 4820
rect 1216 4675 1268 4684
rect 1216 4641 1225 4675
rect 1225 4641 1259 4675
rect 1259 4641 1268 4675
rect 1216 4632 1268 4641
rect 2688 4700 2740 4752
rect 7196 4811 7248 4820
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 11336 4768 11388 4820
rect 6920 4700 6972 4752
rect 3516 4607 3568 4616
rect 3516 4573 3525 4607
rect 3525 4573 3559 4607
rect 3559 4573 3568 4607
rect 3516 4564 3568 4573
rect 7380 4700 7432 4752
rect 9496 4743 9548 4752
rect 9496 4709 9530 4743
rect 9530 4709 9548 4743
rect 9496 4700 9548 4709
rect 10692 4700 10744 4752
rect 9128 4632 9180 4684
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 11796 4632 11848 4684
rect 12164 4743 12216 4752
rect 12164 4709 12173 4743
rect 12173 4709 12207 4743
rect 12207 4709 12216 4743
rect 12164 4700 12216 4709
rect 13268 4768 13320 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 13820 4768 13872 4820
rect 14188 4768 14240 4820
rect 940 4471 992 4480
rect 940 4437 949 4471
rect 949 4437 983 4471
rect 983 4437 992 4471
rect 940 4428 992 4437
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 3424 4471 3476 4480
rect 3424 4437 3433 4471
rect 3433 4437 3467 4471
rect 3467 4437 3476 4471
rect 3424 4428 3476 4437
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 4896 4539 4948 4548
rect 4896 4505 4905 4539
rect 4905 4505 4939 4539
rect 4939 4505 4948 4539
rect 4896 4496 4948 4505
rect 9404 4428 9456 4480
rect 11428 4471 11480 4480
rect 11428 4437 11437 4471
rect 11437 4437 11471 4471
rect 11471 4437 11480 4471
rect 11428 4428 11480 4437
rect 11612 4539 11664 4548
rect 11612 4505 11621 4539
rect 11621 4505 11655 4539
rect 11655 4505 11664 4539
rect 11612 4496 11664 4505
rect 13084 4564 13136 4616
rect 13452 4675 13504 4684
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 13452 4632 13504 4641
rect 13636 4632 13688 4684
rect 14280 4632 14332 4684
rect 13360 4564 13412 4616
rect 14740 4700 14792 4752
rect 15384 4700 15436 4752
rect 15660 4700 15712 4752
rect 14648 4564 14700 4616
rect 14832 4564 14884 4616
rect 15200 4564 15252 4616
rect 16304 4768 16356 4820
rect 16764 4700 16816 4752
rect 18604 4811 18656 4820
rect 18604 4777 18613 4811
rect 18613 4777 18647 4811
rect 18647 4777 18656 4811
rect 18604 4768 18656 4777
rect 18972 4811 19024 4820
rect 18972 4777 18981 4811
rect 18981 4777 19015 4811
rect 19015 4777 19024 4811
rect 18972 4768 19024 4777
rect 19156 4768 19208 4820
rect 19432 4768 19484 4820
rect 20168 4768 20220 4820
rect 18052 4675 18104 4684
rect 18052 4641 18061 4675
rect 18061 4641 18095 4675
rect 18095 4641 18104 4675
rect 18052 4632 18104 4641
rect 18696 4632 18748 4684
rect 19340 4632 19392 4684
rect 20260 4743 20312 4752
rect 20260 4709 20269 4743
rect 20269 4709 20303 4743
rect 20303 4709 20312 4743
rect 20260 4700 20312 4709
rect 20352 4632 20404 4684
rect 21088 4675 21140 4684
rect 21088 4641 21097 4675
rect 21097 4641 21131 4675
rect 21131 4641 21140 4675
rect 21088 4632 21140 4641
rect 21364 4632 21416 4684
rect 22192 4700 22244 4752
rect 23020 4811 23072 4820
rect 23020 4777 23029 4811
rect 23029 4777 23063 4811
rect 23063 4777 23072 4811
rect 23020 4768 23072 4777
rect 23112 4768 23164 4820
rect 28264 4700 28316 4752
rect 28724 4700 28776 4752
rect 24768 4632 24820 4684
rect 27712 4675 27764 4684
rect 27712 4641 27730 4675
rect 27730 4641 27764 4675
rect 27712 4632 27764 4641
rect 28908 4675 28960 4684
rect 28908 4641 28917 4675
rect 28917 4641 28951 4675
rect 28951 4641 28960 4675
rect 28908 4632 28960 4641
rect 29092 4743 29144 4752
rect 29092 4709 29101 4743
rect 29101 4709 29135 4743
rect 29135 4709 29144 4743
rect 29092 4700 29144 4709
rect 30564 4675 30616 4684
rect 30564 4641 30582 4675
rect 30582 4641 30616 4675
rect 30564 4632 30616 4641
rect 30748 4632 30800 4684
rect 20168 4564 20220 4616
rect 20260 4564 20312 4616
rect 27988 4607 28040 4616
rect 27988 4573 27997 4607
rect 27997 4573 28031 4607
rect 28031 4573 28040 4607
rect 27988 4564 28040 4573
rect 29828 4564 29880 4616
rect 11980 4428 12032 4480
rect 19984 4496 20036 4548
rect 14004 4428 14056 4480
rect 15476 4428 15528 4480
rect 15844 4428 15896 4480
rect 16488 4428 16540 4480
rect 16948 4471 17000 4480
rect 16948 4437 16957 4471
rect 16957 4437 16991 4471
rect 16991 4437 17000 4471
rect 16948 4428 17000 4437
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 18328 4428 18380 4437
rect 18420 4428 18472 4480
rect 19340 4471 19392 4480
rect 19340 4437 19349 4471
rect 19349 4437 19383 4471
rect 19383 4437 19392 4471
rect 19340 4428 19392 4437
rect 20628 4471 20680 4480
rect 20628 4437 20637 4471
rect 20637 4437 20671 4471
rect 20671 4437 20680 4471
rect 20628 4428 20680 4437
rect 20720 4471 20772 4480
rect 20720 4437 20729 4471
rect 20729 4437 20763 4471
rect 20763 4437 20772 4471
rect 20720 4428 20772 4437
rect 20812 4471 20864 4480
rect 20812 4437 20821 4471
rect 20821 4437 20855 4471
rect 20855 4437 20864 4471
rect 20812 4428 20864 4437
rect 4250 4326 4302 4378
rect 4314 4326 4366 4378
rect 4378 4326 4430 4378
rect 4442 4326 4494 4378
rect 4506 4326 4558 4378
rect 11955 4326 12007 4378
rect 12019 4326 12071 4378
rect 12083 4326 12135 4378
rect 12147 4326 12199 4378
rect 12211 4326 12263 4378
rect 19660 4326 19712 4378
rect 19724 4326 19776 4378
rect 19788 4326 19840 4378
rect 19852 4326 19904 4378
rect 19916 4326 19968 4378
rect 27365 4326 27417 4378
rect 27429 4326 27481 4378
rect 27493 4326 27545 4378
rect 27557 4326 27609 4378
rect 27621 4326 27673 4378
rect 1216 4224 1268 4276
rect 1492 4224 1544 4276
rect 1952 4156 2004 4208
rect 3424 4224 3476 4276
rect 11520 4224 11572 4276
rect 11888 4224 11940 4276
rect 13636 4224 13688 4276
rect 14004 4224 14056 4276
rect 14832 4224 14884 4276
rect 15200 4224 15252 4276
rect 15292 4267 15344 4276
rect 15292 4233 15301 4267
rect 15301 4233 15335 4267
rect 15335 4233 15344 4267
rect 15292 4224 15344 4233
rect 15660 4224 15712 4276
rect 16580 4224 16632 4276
rect 16764 4267 16816 4276
rect 16764 4233 16773 4267
rect 16773 4233 16807 4267
rect 16807 4233 16816 4267
rect 16764 4224 16816 4233
rect 17408 4224 17460 4276
rect 18052 4267 18104 4276
rect 18052 4233 18061 4267
rect 18061 4233 18095 4267
rect 18095 4233 18104 4267
rect 18052 4224 18104 4233
rect 18328 4224 18380 4276
rect 20168 4224 20220 4276
rect 20260 4224 20312 4276
rect 20720 4224 20772 4276
rect 21732 4267 21784 4276
rect 21732 4233 21741 4267
rect 21741 4233 21775 4267
rect 21775 4233 21784 4267
rect 21732 4224 21784 4233
rect 22652 4224 22704 4276
rect 2320 4088 2372 4140
rect 940 4020 992 4072
rect 1860 4063 1912 4072
rect 1860 4029 1869 4063
rect 1869 4029 1903 4063
rect 1903 4029 1912 4063
rect 1860 4020 1912 4029
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 2228 4063 2280 4072
rect 2228 4029 2237 4063
rect 2237 4029 2271 4063
rect 2271 4029 2280 4063
rect 2228 4020 2280 4029
rect 3516 4020 3568 4072
rect 7288 4020 7340 4072
rect 9312 4020 9364 4072
rect 9404 4020 9456 4072
rect 10692 4088 10744 4140
rect 14372 4156 14424 4208
rect 2504 3952 2556 4004
rect 5448 3952 5500 4004
rect 11336 4020 11388 4072
rect 2044 3884 2096 3936
rect 11520 3995 11572 4004
rect 11520 3961 11529 3995
rect 11529 3961 11563 3995
rect 11563 3961 11572 3995
rect 11520 3952 11572 3961
rect 11796 3952 11848 4004
rect 12532 3952 12584 4004
rect 12624 3952 12676 4004
rect 9128 3884 9180 3936
rect 13820 3884 13872 3936
rect 14280 3995 14332 4004
rect 14280 3961 14289 3995
rect 14289 3961 14323 3995
rect 14323 3961 14332 3995
rect 14280 3952 14332 3961
rect 14648 3952 14700 4004
rect 14832 4020 14884 4072
rect 15568 4020 15620 4072
rect 15844 4020 15896 4072
rect 19616 4088 19668 4140
rect 20076 4088 20128 4140
rect 17500 4063 17552 4072
rect 17500 4029 17509 4063
rect 17509 4029 17543 4063
rect 17543 4029 17552 4063
rect 17500 4020 17552 4029
rect 22836 4224 22888 4276
rect 22928 4224 22980 4276
rect 23112 4224 23164 4276
rect 24124 4224 24176 4276
rect 22652 4088 22704 4140
rect 23112 4088 23164 4140
rect 24032 4088 24084 4140
rect 16856 3952 16908 4004
rect 16948 3995 17000 4004
rect 16948 3961 16957 3995
rect 16957 3961 16991 3995
rect 16991 3961 17000 3995
rect 16948 3952 17000 3961
rect 17316 3952 17368 4004
rect 17960 3952 18012 4004
rect 16580 3927 16632 3936
rect 16580 3893 16589 3927
rect 16589 3893 16623 3927
rect 16623 3893 16632 3927
rect 16580 3884 16632 3893
rect 17040 3884 17092 3936
rect 21456 3952 21508 4004
rect 22376 3952 22428 4004
rect 21824 3884 21876 3936
rect 22560 3927 22612 3936
rect 22560 3893 22569 3927
rect 22569 3893 22603 3927
rect 22603 3893 22612 3927
rect 22560 3884 22612 3893
rect 22928 3995 22980 4004
rect 22928 3961 22937 3995
rect 22937 3961 22971 3995
rect 22971 3961 22980 3995
rect 22928 3952 22980 3961
rect 23296 3952 23348 4004
rect 23204 3927 23256 3936
rect 23204 3893 23221 3927
rect 23221 3893 23256 3927
rect 23204 3884 23256 3893
rect 23940 4020 23992 4072
rect 24768 4267 24820 4276
rect 24768 4233 24777 4267
rect 24777 4233 24811 4267
rect 24811 4233 24820 4267
rect 24768 4224 24820 4233
rect 29828 4224 29880 4276
rect 26056 4020 26108 4072
rect 27988 4063 28040 4072
rect 27988 4029 27997 4063
rect 27997 4029 28031 4063
rect 28031 4029 28040 4063
rect 27988 4020 28040 4029
rect 24584 3952 24636 4004
rect 26332 3952 26384 4004
rect 27252 3952 27304 4004
rect 28264 3952 28316 4004
rect 24492 3927 24544 3936
rect 24492 3893 24519 3927
rect 24519 3893 24544 3927
rect 24492 3884 24544 3893
rect 26608 3927 26660 3936
rect 26608 3893 26617 3927
rect 26617 3893 26651 3927
rect 26651 3893 26660 3927
rect 26608 3884 26660 3893
rect 27804 3884 27856 3936
rect 29644 4020 29696 4072
rect 30564 4088 30616 4140
rect 29644 3927 29696 3936
rect 29644 3893 29653 3927
rect 29653 3893 29687 3927
rect 29687 3893 29696 3927
rect 29644 3884 29696 3893
rect 29920 3927 29972 3936
rect 29920 3893 29929 3927
rect 29929 3893 29963 3927
rect 29963 3893 29972 3927
rect 29920 3884 29972 3893
rect 30472 3927 30524 3936
rect 30472 3893 30481 3927
rect 30481 3893 30515 3927
rect 30515 3893 30524 3927
rect 30472 3884 30524 3893
rect 8102 3782 8154 3834
rect 8166 3782 8218 3834
rect 8230 3782 8282 3834
rect 8294 3782 8346 3834
rect 8358 3782 8410 3834
rect 15807 3782 15859 3834
rect 15871 3782 15923 3834
rect 15935 3782 15987 3834
rect 15999 3782 16051 3834
rect 16063 3782 16115 3834
rect 23512 3782 23564 3834
rect 23576 3782 23628 3834
rect 23640 3782 23692 3834
rect 23704 3782 23756 3834
rect 23768 3782 23820 3834
rect 31217 3782 31269 3834
rect 31281 3782 31333 3834
rect 31345 3782 31397 3834
rect 31409 3782 31461 3834
rect 31473 3782 31525 3834
rect 940 3680 992 3732
rect 1860 3680 1912 3732
rect 2504 3723 2556 3732
rect 2504 3689 2513 3723
rect 2513 3689 2547 3723
rect 2547 3689 2556 3723
rect 2504 3680 2556 3689
rect 2044 3587 2096 3596
rect 2044 3553 2053 3587
rect 2053 3553 2087 3587
rect 2087 3553 2096 3587
rect 2044 3544 2096 3553
rect 2320 3587 2372 3596
rect 2320 3553 2329 3587
rect 2329 3553 2363 3587
rect 2363 3553 2372 3587
rect 2320 3544 2372 3553
rect 3516 3680 3568 3732
rect 2136 3476 2188 3528
rect 3056 3587 3108 3596
rect 3056 3553 3090 3587
rect 3090 3553 3108 3587
rect 3056 3544 3108 3553
rect 7288 3612 7340 3664
rect 6828 3587 6880 3596
rect 6828 3553 6862 3587
rect 6862 3553 6880 3587
rect 6828 3544 6880 3553
rect 8116 3544 8168 3596
rect 11612 3612 11664 3664
rect 13912 3680 13964 3732
rect 14832 3723 14884 3732
rect 12624 3544 12676 3596
rect 12716 3544 12768 3596
rect 13452 3655 13504 3664
rect 13452 3621 13461 3655
rect 13461 3621 13495 3655
rect 13495 3621 13504 3655
rect 13452 3612 13504 3621
rect 13268 3544 13320 3596
rect 14832 3689 14859 3723
rect 14859 3689 14884 3723
rect 14832 3680 14884 3689
rect 15108 3723 15160 3732
rect 15108 3689 15117 3723
rect 15117 3689 15151 3723
rect 15151 3689 15160 3723
rect 15108 3680 15160 3689
rect 16488 3723 16540 3732
rect 14188 3655 14240 3664
rect 14188 3621 14197 3655
rect 14197 3621 14231 3655
rect 14231 3621 14240 3655
rect 14188 3612 14240 3621
rect 14648 3612 14700 3664
rect 7932 3476 7984 3528
rect 13452 3476 13504 3528
rect 14464 3476 14516 3528
rect 14924 3544 14976 3596
rect 16488 3689 16513 3723
rect 16513 3689 16540 3723
rect 16488 3680 16540 3689
rect 16212 3612 16264 3664
rect 16304 3655 16356 3664
rect 16304 3621 16313 3655
rect 16313 3621 16347 3655
rect 16347 3621 16356 3655
rect 16304 3612 16356 3621
rect 16672 3723 16724 3732
rect 16672 3689 16681 3723
rect 16681 3689 16715 3723
rect 16715 3689 16724 3723
rect 16672 3680 16724 3689
rect 17224 3723 17276 3732
rect 17224 3689 17249 3723
rect 17249 3689 17276 3723
rect 17224 3680 17276 3689
rect 17132 3612 17184 3664
rect 17500 3680 17552 3732
rect 18880 3723 18932 3732
rect 18880 3689 18889 3723
rect 18889 3689 18923 3723
rect 18923 3689 18932 3723
rect 18880 3680 18932 3689
rect 19340 3723 19392 3732
rect 19340 3689 19349 3723
rect 19349 3689 19383 3723
rect 19383 3689 19392 3723
rect 19340 3680 19392 3689
rect 19616 3680 19668 3732
rect 19064 3655 19116 3664
rect 19064 3621 19075 3655
rect 19075 3621 19116 3655
rect 19064 3612 19116 3621
rect 19156 3612 19208 3664
rect 19984 3612 20036 3664
rect 20628 3680 20680 3732
rect 21272 3723 21324 3732
rect 21272 3689 21281 3723
rect 21281 3689 21315 3723
rect 21315 3689 21324 3723
rect 21272 3680 21324 3689
rect 21916 3723 21968 3732
rect 21916 3689 21943 3723
rect 21943 3689 21968 3723
rect 21916 3680 21968 3689
rect 22652 3680 22704 3732
rect 23204 3680 23256 3732
rect 3056 3340 3108 3392
rect 11980 3340 12032 3392
rect 12808 3340 12860 3392
rect 13728 3408 13780 3460
rect 13820 3408 13872 3460
rect 13544 3340 13596 3392
rect 13636 3383 13688 3392
rect 13636 3349 13645 3383
rect 13645 3349 13679 3383
rect 13679 3349 13688 3383
rect 13636 3340 13688 3349
rect 14556 3451 14608 3460
rect 14556 3417 14565 3451
rect 14565 3417 14599 3451
rect 14599 3417 14608 3451
rect 14556 3408 14608 3417
rect 19064 3476 19116 3528
rect 18420 3408 18472 3460
rect 21548 3612 21600 3664
rect 22008 3612 22060 3664
rect 19524 3476 19576 3528
rect 15200 3340 15252 3392
rect 16764 3340 16816 3392
rect 18052 3340 18104 3392
rect 18972 3340 19024 3392
rect 19064 3383 19116 3392
rect 19064 3349 19073 3383
rect 19073 3349 19107 3383
rect 19107 3349 19116 3383
rect 19064 3340 19116 3349
rect 19248 3340 19300 3392
rect 20720 3340 20772 3392
rect 21732 3340 21784 3392
rect 24400 3680 24452 3732
rect 24584 3723 24636 3732
rect 24584 3689 24593 3723
rect 24593 3689 24627 3723
rect 24627 3689 24636 3723
rect 24584 3680 24636 3689
rect 27252 3723 27304 3732
rect 27252 3689 27261 3723
rect 27261 3689 27295 3723
rect 27295 3689 27304 3723
rect 27252 3680 27304 3689
rect 27712 3680 27764 3732
rect 24492 3612 24544 3664
rect 25596 3612 25648 3664
rect 28264 3680 28316 3732
rect 28908 3680 28960 3732
rect 29644 3680 29696 3732
rect 25412 3544 25464 3596
rect 27160 3587 27212 3596
rect 27160 3553 27169 3587
rect 27169 3553 27203 3587
rect 27203 3553 27212 3587
rect 27160 3544 27212 3553
rect 27252 3544 27304 3596
rect 27988 3544 28040 3596
rect 29092 3587 29144 3596
rect 29092 3553 29101 3587
rect 29101 3553 29135 3587
rect 29135 3553 29144 3587
rect 29092 3544 29144 3553
rect 29920 3612 29972 3664
rect 25228 3340 25280 3392
rect 26056 3476 26108 3528
rect 30932 3383 30984 3392
rect 30932 3349 30941 3383
rect 30941 3349 30975 3383
rect 30975 3349 30984 3383
rect 30932 3340 30984 3349
rect 4250 3238 4302 3290
rect 4314 3238 4366 3290
rect 4378 3238 4430 3290
rect 4442 3238 4494 3290
rect 4506 3238 4558 3290
rect 11955 3238 12007 3290
rect 12019 3238 12071 3290
rect 12083 3238 12135 3290
rect 12147 3238 12199 3290
rect 12211 3238 12263 3290
rect 19660 3238 19712 3290
rect 19724 3238 19776 3290
rect 19788 3238 19840 3290
rect 19852 3238 19904 3290
rect 19916 3238 19968 3290
rect 27365 3238 27417 3290
rect 27429 3238 27481 3290
rect 27493 3238 27545 3290
rect 27557 3238 27609 3290
rect 27621 3238 27673 3290
rect 3056 3136 3108 3188
rect 7196 3136 7248 3188
rect 8116 3136 8168 3188
rect 11520 3136 11572 3188
rect 12716 3136 12768 3188
rect 12808 3136 12860 3188
rect 11244 3068 11296 3120
rect 13176 3179 13228 3188
rect 13176 3145 13185 3179
rect 13185 3145 13219 3179
rect 13219 3145 13228 3179
rect 13176 3136 13228 3145
rect 13360 3136 13412 3188
rect 14464 3136 14516 3188
rect 14924 3179 14976 3188
rect 14924 3145 14933 3179
rect 14933 3145 14967 3179
rect 14967 3145 14976 3179
rect 14924 3136 14976 3145
rect 16948 3136 17000 3188
rect 19064 3136 19116 3188
rect 20812 3136 20864 3188
rect 21456 3136 21508 3188
rect 21548 3179 21600 3188
rect 21548 3145 21557 3179
rect 21557 3145 21591 3179
rect 21591 3145 21600 3179
rect 21548 3136 21600 3145
rect 23296 3179 23348 3188
rect 23296 3145 23305 3179
rect 23305 3145 23339 3179
rect 23339 3145 23348 3179
rect 23296 3136 23348 3145
rect 23388 3136 23440 3188
rect 25412 3068 25464 3120
rect 27252 3068 27304 3120
rect 29092 3179 29144 3188
rect 29092 3145 29101 3179
rect 29101 3145 29135 3179
rect 29135 3145 29144 3179
rect 29092 3136 29144 3145
rect 30472 3136 30524 3188
rect 30932 3136 30984 3188
rect 7932 3000 7984 3052
rect 1860 2977 1912 2984
rect 1860 2943 1869 2977
rect 1869 2943 1903 2977
rect 1903 2943 1912 2977
rect 1860 2932 1912 2943
rect 2136 2975 2188 2984
rect 2136 2941 2145 2975
rect 2145 2941 2179 2975
rect 2179 2941 2188 2975
rect 2136 2932 2188 2941
rect 2504 2932 2556 2984
rect 9404 2932 9456 2984
rect 12440 2932 12492 2984
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 15476 2932 15528 2984
rect 20076 2975 20128 2984
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 21180 2932 21232 2984
rect 21916 2975 21968 2984
rect 21916 2941 21925 2975
rect 21925 2941 21959 2975
rect 21959 2941 21968 2975
rect 21916 2932 21968 2941
rect 25136 2932 25188 2984
rect 3976 2864 4028 2916
rect 5448 2864 5500 2916
rect 7104 2907 7156 2916
rect 7104 2873 7116 2907
rect 7116 2873 7156 2907
rect 7104 2864 7156 2873
rect 9864 2907 9916 2916
rect 9864 2873 9898 2907
rect 9898 2873 9916 2907
rect 9864 2864 9916 2873
rect 10416 2864 10468 2916
rect 11060 2864 11112 2916
rect 12808 2907 12860 2916
rect 12808 2873 12817 2907
rect 12817 2873 12851 2907
rect 12851 2873 12860 2907
rect 12808 2864 12860 2873
rect 12900 2864 12952 2916
rect 13268 2864 13320 2916
rect 14372 2864 14424 2916
rect 16212 2864 16264 2916
rect 19432 2864 19484 2916
rect 20260 2864 20312 2916
rect 24032 2864 24084 2916
rect 24952 2907 25004 2916
rect 24952 2873 24970 2907
rect 24970 2873 25004 2907
rect 25688 2932 25740 2984
rect 24952 2864 25004 2873
rect 2412 2839 2464 2848
rect 2412 2805 2421 2839
rect 2421 2805 2455 2839
rect 2455 2805 2464 2839
rect 2412 2796 2464 2805
rect 2688 2839 2740 2848
rect 2688 2805 2697 2839
rect 2697 2805 2731 2839
rect 2731 2805 2740 2839
rect 2688 2796 2740 2805
rect 5264 2839 5316 2848
rect 5264 2805 5273 2839
rect 5273 2805 5307 2839
rect 5307 2805 5316 2839
rect 5264 2796 5316 2805
rect 22560 2796 22612 2848
rect 25320 2796 25372 2848
rect 25596 2796 25648 2848
rect 26332 2932 26384 2984
rect 26700 2864 26752 2916
rect 26148 2796 26200 2848
rect 26608 2796 26660 2848
rect 27988 2932 28040 2984
rect 27528 2864 27580 2916
rect 29828 2975 29880 2984
rect 29828 2941 29837 2975
rect 29837 2941 29871 2975
rect 29871 2941 29880 2975
rect 29828 2932 29880 2941
rect 31576 2932 31628 2984
rect 8102 2694 8154 2746
rect 8166 2694 8218 2746
rect 8230 2694 8282 2746
rect 8294 2694 8346 2746
rect 8358 2694 8410 2746
rect 15807 2694 15859 2746
rect 15871 2694 15923 2746
rect 15935 2694 15987 2746
rect 15999 2694 16051 2746
rect 16063 2694 16115 2746
rect 23512 2694 23564 2746
rect 23576 2694 23628 2746
rect 23640 2694 23692 2746
rect 23704 2694 23756 2746
rect 23768 2694 23820 2746
rect 31217 2694 31269 2746
rect 31281 2694 31333 2746
rect 31345 2694 31397 2746
rect 31409 2694 31461 2746
rect 31473 2694 31525 2746
rect 2412 2635 2464 2644
rect 2412 2601 2421 2635
rect 2421 2601 2455 2635
rect 2455 2601 2464 2635
rect 2412 2592 2464 2601
rect 2688 2524 2740 2576
rect 3976 2592 4028 2644
rect 11612 2592 11664 2644
rect 13084 2592 13136 2644
rect 14648 2592 14700 2644
rect 16304 2592 16356 2644
rect 17960 2635 18012 2644
rect 17960 2601 17969 2635
rect 17969 2601 18003 2635
rect 18003 2601 18012 2635
rect 17960 2592 18012 2601
rect 19524 2635 19576 2644
rect 19524 2601 19533 2635
rect 19533 2601 19567 2635
rect 19567 2601 19576 2635
rect 19524 2592 19576 2601
rect 20260 2635 20312 2644
rect 20260 2601 20269 2635
rect 20269 2601 20303 2635
rect 20303 2601 20312 2635
rect 20260 2592 20312 2601
rect 24032 2635 24084 2644
rect 24032 2601 24041 2635
rect 24041 2601 24075 2635
rect 24075 2601 24084 2635
rect 24032 2592 24084 2601
rect 2780 2456 2832 2508
rect 5356 2524 5408 2576
rect 7012 2524 7064 2576
rect 3332 2320 3384 2372
rect 7932 2499 7984 2508
rect 7932 2465 7941 2499
rect 7941 2465 7975 2499
rect 7975 2465 7984 2499
rect 7932 2456 7984 2465
rect 8208 2499 8260 2508
rect 8208 2465 8242 2499
rect 8242 2465 8260 2499
rect 8208 2456 8260 2465
rect 9404 2499 9456 2508
rect 9404 2465 9413 2499
rect 9413 2465 9447 2499
rect 9447 2465 9456 2499
rect 9404 2456 9456 2465
rect 9680 2499 9732 2508
rect 9680 2465 9714 2499
rect 9714 2465 9732 2499
rect 9680 2456 9732 2465
rect 11520 2456 11572 2508
rect 11704 2456 11756 2508
rect 13636 2524 13688 2576
rect 13176 2456 13228 2508
rect 13728 2456 13780 2508
rect 15476 2524 15528 2576
rect 16212 2388 16264 2440
rect 16856 2499 16908 2508
rect 16856 2465 16890 2499
rect 16890 2465 16908 2499
rect 16856 2456 16908 2465
rect 21916 2524 21968 2576
rect 25596 2592 25648 2644
rect 26608 2635 26660 2644
rect 26608 2601 26617 2635
rect 26617 2601 26651 2635
rect 26651 2601 26660 2635
rect 26608 2592 26660 2601
rect 26700 2592 26752 2644
rect 27160 2592 27212 2644
rect 27528 2635 27580 2644
rect 27528 2601 27537 2635
rect 27537 2601 27571 2635
rect 27571 2601 27580 2635
rect 27528 2592 27580 2601
rect 26148 2567 26200 2576
rect 18236 2456 18288 2508
rect 20168 2499 20220 2508
rect 20168 2465 20177 2499
rect 20177 2465 20211 2499
rect 20211 2465 20220 2499
rect 20168 2456 20220 2465
rect 22836 2499 22888 2508
rect 26148 2533 26157 2567
rect 26157 2533 26191 2567
rect 26191 2533 26200 2567
rect 26148 2524 26200 2533
rect 22836 2465 22854 2499
rect 22854 2465 22888 2499
rect 22836 2456 22888 2465
rect 24124 2499 24176 2508
rect 24124 2465 24133 2499
rect 24133 2465 24167 2499
rect 24167 2465 24176 2499
rect 24124 2456 24176 2465
rect 25320 2456 25372 2508
rect 25596 2456 25648 2508
rect 27252 2456 27304 2508
rect 4620 2252 4672 2304
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 7288 2295 7340 2304
rect 7288 2261 7297 2295
rect 7297 2261 7331 2295
rect 7331 2261 7340 2295
rect 7288 2252 7340 2261
rect 25688 2388 25740 2440
rect 26332 2320 26384 2372
rect 14188 2252 14240 2304
rect 15568 2252 15620 2304
rect 24492 2252 24544 2304
rect 24952 2252 25004 2304
rect 25412 2252 25464 2304
rect 25596 2295 25648 2304
rect 25596 2261 25605 2295
rect 25605 2261 25639 2295
rect 25639 2261 25648 2295
rect 25596 2252 25648 2261
rect 31024 2295 31076 2304
rect 31024 2261 31033 2295
rect 31033 2261 31067 2295
rect 31067 2261 31076 2295
rect 31024 2252 31076 2261
rect 4250 2150 4302 2202
rect 4314 2150 4366 2202
rect 4378 2150 4430 2202
rect 4442 2150 4494 2202
rect 4506 2150 4558 2202
rect 11955 2150 12007 2202
rect 12019 2150 12071 2202
rect 12083 2150 12135 2202
rect 12147 2150 12199 2202
rect 12211 2150 12263 2202
rect 19660 2150 19712 2202
rect 19724 2150 19776 2202
rect 19788 2150 19840 2202
rect 19852 2150 19904 2202
rect 19916 2150 19968 2202
rect 27365 2150 27417 2202
rect 27429 2150 27481 2202
rect 27493 2150 27545 2202
rect 27557 2150 27609 2202
rect 27621 2150 27673 2202
rect 2688 2091 2740 2100
rect 2688 2057 2697 2091
rect 2697 2057 2731 2091
rect 2731 2057 2740 2091
rect 2688 2048 2740 2057
rect 3332 2091 3384 2100
rect 3332 2057 3341 2091
rect 3341 2057 3375 2091
rect 3375 2057 3384 2091
rect 3332 2048 3384 2057
rect 7196 2091 7248 2100
rect 7196 2057 7205 2091
rect 7205 2057 7239 2091
rect 7239 2057 7248 2091
rect 7196 2048 7248 2057
rect 7840 2048 7892 2100
rect 8208 2048 8260 2100
rect 9680 2048 9732 2100
rect 4712 1980 4764 2032
rect 2780 1887 2832 1896
rect 2780 1853 2789 1887
rect 2789 1853 2823 1887
rect 2823 1853 2832 1887
rect 2780 1844 2832 1853
rect 4620 1887 4672 1896
rect 4620 1853 4629 1887
rect 4629 1853 4663 1887
rect 4663 1853 4672 1887
rect 4620 1844 4672 1853
rect 5172 1887 5224 1896
rect 5172 1853 5173 1887
rect 5173 1853 5207 1887
rect 5207 1853 5224 1887
rect 5172 1844 5224 1853
rect 5448 1887 5500 1896
rect 5448 1853 5457 1887
rect 5457 1853 5491 1887
rect 5491 1853 5500 1887
rect 5448 1844 5500 1853
rect 6828 1980 6880 2032
rect 7012 1980 7064 2032
rect 7288 1980 7340 2032
rect 6828 1887 6880 1896
rect 6828 1853 6837 1887
rect 6837 1853 6871 1887
rect 6871 1853 6880 1887
rect 6828 1844 6880 1853
rect 8116 1844 8168 1896
rect 9496 1887 9548 1896
rect 9496 1853 9505 1887
rect 9505 1853 9539 1887
rect 9539 1853 9548 1887
rect 9496 1844 9548 1853
rect 11152 2048 11204 2100
rect 11520 2048 11572 2100
rect 12992 2048 13044 2100
rect 16120 2091 16172 2100
rect 16120 2057 16129 2091
rect 16129 2057 16163 2091
rect 16163 2057 16172 2091
rect 16120 2048 16172 2057
rect 17960 2048 18012 2100
rect 18236 2048 18288 2100
rect 20168 2048 20220 2100
rect 22008 2048 22060 2100
rect 22376 2048 22428 2100
rect 24124 2048 24176 2100
rect 24492 2091 24544 2100
rect 24492 2057 24501 2091
rect 24501 2057 24535 2091
rect 24535 2057 24544 2091
rect 24492 2048 24544 2057
rect 16856 1912 16908 1964
rect 9864 1844 9916 1896
rect 11612 1844 11664 1896
rect 10600 1776 10652 1828
rect 15200 1887 15252 1896
rect 15200 1853 15209 1887
rect 15209 1853 15243 1887
rect 15243 1853 15252 1887
rect 15200 1844 15252 1853
rect 15476 1889 15528 1896
rect 15476 1855 15485 1889
rect 15485 1855 15519 1889
rect 15519 1855 15528 1889
rect 15476 1844 15528 1855
rect 15660 1844 15712 1896
rect 16304 1887 16356 1896
rect 16304 1853 16313 1887
rect 16313 1853 16347 1887
rect 16347 1853 16356 1887
rect 16304 1844 16356 1853
rect 9404 1751 9456 1760
rect 9404 1717 9413 1751
rect 9413 1717 9447 1751
rect 9447 1717 9456 1751
rect 9404 1708 9456 1717
rect 9680 1751 9732 1760
rect 9680 1717 9689 1751
rect 9689 1717 9723 1751
rect 9723 1717 9732 1751
rect 9680 1708 9732 1717
rect 12348 1751 12400 1760
rect 12348 1717 12357 1751
rect 12357 1717 12391 1751
rect 12391 1717 12400 1751
rect 12348 1708 12400 1717
rect 12624 1751 12676 1760
rect 12624 1717 12633 1751
rect 12633 1717 12667 1751
rect 12667 1717 12676 1751
rect 12624 1708 12676 1717
rect 14464 1751 14516 1760
rect 14464 1717 14473 1751
rect 14473 1717 14507 1751
rect 14507 1717 14516 1751
rect 14464 1708 14516 1717
rect 14556 1708 14608 1760
rect 16856 1751 16908 1760
rect 16856 1717 16865 1751
rect 16865 1717 16899 1751
rect 16899 1717 16908 1751
rect 17960 1887 18012 1896
rect 17960 1853 17969 1887
rect 17969 1853 18003 1887
rect 18003 1853 18012 1887
rect 17960 1844 18012 1853
rect 18696 1912 18748 1964
rect 20076 1912 20128 1964
rect 24492 1912 24544 1964
rect 17592 1776 17644 1828
rect 19064 1844 19116 1896
rect 16856 1708 16908 1717
rect 18788 1708 18840 1760
rect 19432 1776 19484 1828
rect 20444 1776 20496 1828
rect 22836 1844 22888 1896
rect 25136 1912 25188 1964
rect 31024 1887 31076 1896
rect 31024 1853 31033 1887
rect 31033 1853 31067 1887
rect 31067 1853 31076 1887
rect 31024 1844 31076 1853
rect 19524 1708 19576 1760
rect 22008 1708 22060 1760
rect 22100 1708 22152 1760
rect 24216 1708 24268 1760
rect 8102 1606 8154 1658
rect 8166 1606 8218 1658
rect 8230 1606 8282 1658
rect 8294 1606 8346 1658
rect 8358 1606 8410 1658
rect 15807 1606 15859 1658
rect 15871 1606 15923 1658
rect 15935 1606 15987 1658
rect 15999 1606 16051 1658
rect 16063 1606 16115 1658
rect 23512 1606 23564 1658
rect 23576 1606 23628 1658
rect 23640 1606 23692 1658
rect 23704 1606 23756 1658
rect 23768 1606 23820 1658
rect 31217 1606 31269 1658
rect 31281 1606 31333 1658
rect 31345 1606 31397 1658
rect 31409 1606 31461 1658
rect 31473 1606 31525 1658
rect 7196 1504 7248 1556
rect 7288 1504 7340 1556
rect 7840 1504 7892 1556
rect 8484 1436 8536 1488
rect 8024 1300 8076 1352
rect 9496 1504 9548 1556
rect 9404 1436 9456 1488
rect 9680 1411 9732 1420
rect 9680 1377 9689 1411
rect 9689 1377 9723 1411
rect 9723 1377 9732 1411
rect 9680 1368 9732 1377
rect 10600 1368 10652 1420
rect 11060 1479 11112 1488
rect 11060 1445 11069 1479
rect 11069 1445 11103 1479
rect 11103 1445 11112 1479
rect 11060 1436 11112 1445
rect 11152 1436 11204 1488
rect 11612 1504 11664 1556
rect 12808 1504 12860 1556
rect 13176 1504 13228 1556
rect 14556 1504 14608 1556
rect 12624 1368 12676 1420
rect 13176 1368 13228 1420
rect 14464 1436 14516 1488
rect 14740 1504 14792 1556
rect 15200 1436 15252 1488
rect 15476 1504 15528 1556
rect 15660 1504 15712 1556
rect 16304 1504 16356 1556
rect 16396 1547 16448 1556
rect 16396 1513 16405 1547
rect 16405 1513 16439 1547
rect 16439 1513 16448 1547
rect 16396 1504 16448 1513
rect 16856 1504 16908 1556
rect 17592 1504 17644 1556
rect 17776 1504 17828 1556
rect 17960 1547 18012 1556
rect 17960 1513 17969 1547
rect 17969 1513 18003 1547
rect 18003 1513 18012 1547
rect 17960 1504 18012 1513
rect 18052 1504 18104 1556
rect 18512 1547 18564 1556
rect 18512 1513 18521 1547
rect 18521 1513 18555 1547
rect 18555 1513 18564 1547
rect 18512 1504 18564 1513
rect 18788 1547 18840 1556
rect 18788 1513 18797 1547
rect 18797 1513 18831 1547
rect 18831 1513 18840 1547
rect 18788 1504 18840 1513
rect 19064 1547 19116 1556
rect 19064 1513 19073 1547
rect 19073 1513 19107 1547
rect 19107 1513 19116 1547
rect 19064 1504 19116 1513
rect 19432 1504 19484 1556
rect 20076 1504 20128 1556
rect 20260 1504 20312 1556
rect 13728 1300 13780 1352
rect 14372 1232 14424 1284
rect 16304 1368 16356 1420
rect 17500 1411 17552 1420
rect 17500 1377 17509 1411
rect 17509 1377 17543 1411
rect 17543 1377 17552 1411
rect 17500 1368 17552 1377
rect 18236 1411 18288 1420
rect 18236 1377 18245 1411
rect 18245 1377 18279 1411
rect 18279 1377 18288 1411
rect 18236 1368 18288 1377
rect 22008 1504 22060 1556
rect 22468 1547 22520 1556
rect 22468 1513 22477 1547
rect 22477 1513 22511 1547
rect 22511 1513 22520 1547
rect 22468 1504 22520 1513
rect 22836 1504 22888 1556
rect 23848 1504 23900 1556
rect 25412 1547 25464 1556
rect 25412 1513 25421 1547
rect 25421 1513 25455 1547
rect 25455 1513 25464 1547
rect 25412 1504 25464 1513
rect 19524 1411 19576 1420
rect 19524 1377 19533 1411
rect 19533 1377 19567 1411
rect 19567 1377 19576 1411
rect 19524 1368 19576 1377
rect 17592 1232 17644 1284
rect 20168 1300 20220 1352
rect 20444 1411 20496 1420
rect 20444 1377 20453 1411
rect 20453 1377 20487 1411
rect 20487 1377 20496 1411
rect 20444 1368 20496 1377
rect 24216 1436 24268 1488
rect 20076 1232 20128 1284
rect 21824 1411 21876 1420
rect 21824 1377 21833 1411
rect 21833 1377 21867 1411
rect 21867 1377 21876 1411
rect 21824 1368 21876 1377
rect 21732 1300 21784 1352
rect 22928 1411 22980 1420
rect 22928 1377 22937 1411
rect 22937 1377 22971 1411
rect 22971 1377 22980 1411
rect 22928 1368 22980 1377
rect 23572 1411 23624 1420
rect 23572 1377 23581 1411
rect 23581 1377 23615 1411
rect 23615 1377 23624 1411
rect 23572 1368 23624 1377
rect 24584 1368 24636 1420
rect 25136 1411 25188 1420
rect 25136 1377 25145 1411
rect 25145 1377 25179 1411
rect 25179 1377 25188 1411
rect 25136 1368 25188 1377
rect 11612 1164 11664 1216
rect 14188 1207 14240 1216
rect 14188 1173 14197 1207
rect 14197 1173 14231 1207
rect 14231 1173 14240 1207
rect 14188 1164 14240 1173
rect 14648 1164 14700 1216
rect 14740 1164 14792 1216
rect 21272 1164 21324 1216
rect 22100 1164 22152 1216
rect 4250 1062 4302 1114
rect 4314 1062 4366 1114
rect 4378 1062 4430 1114
rect 4442 1062 4494 1114
rect 4506 1062 4558 1114
rect 11955 1062 12007 1114
rect 12019 1062 12071 1114
rect 12083 1062 12135 1114
rect 12147 1062 12199 1114
rect 12211 1062 12263 1114
rect 19660 1062 19712 1114
rect 19724 1062 19776 1114
rect 19788 1062 19840 1114
rect 19852 1062 19904 1114
rect 19916 1062 19968 1114
rect 27365 1062 27417 1114
rect 27429 1062 27481 1114
rect 27493 1062 27545 1114
rect 27557 1062 27609 1114
rect 27621 1062 27673 1114
rect 8024 960 8076 1012
rect 8484 1003 8536 1012
rect 8484 969 8493 1003
rect 8493 969 8527 1003
rect 8527 969 8536 1003
rect 8484 960 8536 969
rect 9404 1003 9456 1012
rect 9404 969 9413 1003
rect 9413 969 9447 1003
rect 9447 969 9456 1003
rect 9404 960 9456 969
rect 9680 960 9732 1012
rect 11060 960 11112 1012
rect 11704 892 11756 944
rect 9864 824 9916 876
rect 7840 756 7892 808
rect 10600 756 10652 808
rect 12624 960 12676 1012
rect 14188 960 14240 1012
rect 14464 1003 14516 1012
rect 14464 969 14473 1003
rect 14473 969 14507 1003
rect 14507 969 14516 1003
rect 14464 960 14516 969
rect 15016 960 15068 1012
rect 17132 960 17184 1012
rect 19984 960 20036 1012
rect 20444 960 20496 1012
rect 21824 960 21876 1012
rect 22100 960 22152 1012
rect 22468 960 22520 1012
rect 14740 935 14792 944
rect 14740 901 14749 935
rect 14749 901 14783 935
rect 14783 901 14792 935
rect 14740 892 14792 901
rect 12348 799 12400 808
rect 12348 765 12357 799
rect 12357 765 12391 799
rect 12391 765 12400 799
rect 12348 756 12400 765
rect 13176 799 13228 808
rect 13176 765 13185 799
rect 13185 765 13219 799
rect 13219 765 13228 799
rect 13176 756 13228 765
rect 13728 756 13780 808
rect 14648 799 14700 808
rect 14648 765 14657 799
rect 14657 765 14691 799
rect 14691 765 14700 799
rect 14648 756 14700 765
rect 18696 867 18748 876
rect 15660 731 15712 740
rect 15660 697 15669 731
rect 15669 697 15703 731
rect 15703 697 15712 731
rect 15660 688 15712 697
rect 16212 756 16264 808
rect 18696 833 18705 867
rect 18705 833 18739 867
rect 18739 833 18748 867
rect 18696 824 18748 833
rect 16764 688 16816 740
rect 17868 799 17920 808
rect 17868 765 17877 799
rect 17877 765 17911 799
rect 17911 765 17920 799
rect 17868 756 17920 765
rect 19524 756 19576 808
rect 21272 799 21324 808
rect 21272 765 21281 799
rect 21281 765 21315 799
rect 21315 765 21324 799
rect 21272 756 21324 765
rect 21732 799 21784 808
rect 21732 765 21741 799
rect 21741 765 21775 799
rect 21775 765 21784 799
rect 21732 756 21784 765
rect 21916 824 21968 876
rect 22928 756 22980 808
rect 23572 960 23624 1012
rect 23848 892 23900 944
rect 24216 1003 24268 1012
rect 24216 969 24225 1003
rect 24225 969 24259 1003
rect 24259 969 24268 1003
rect 24216 960 24268 969
rect 24492 1003 24544 1012
rect 24492 969 24501 1003
rect 24501 969 24535 1003
rect 24535 969 24544 1003
rect 24492 960 24544 969
rect 24584 799 24636 808
rect 24584 765 24593 799
rect 24593 765 24627 799
rect 24627 765 24636 799
rect 24584 756 24636 765
rect 31024 799 31076 808
rect 31024 765 31033 799
rect 31033 765 31067 799
rect 31067 765 31076 799
rect 31024 756 31076 765
rect 8102 518 8154 570
rect 8166 518 8218 570
rect 8230 518 8282 570
rect 8294 518 8346 570
rect 8358 518 8410 570
rect 15807 518 15859 570
rect 15871 518 15923 570
rect 15935 518 15987 570
rect 15999 518 16051 570
rect 16063 518 16115 570
rect 23512 518 23564 570
rect 23576 518 23628 570
rect 23640 518 23692 570
rect 23704 518 23756 570
rect 23768 518 23820 570
rect 31217 518 31269 570
rect 31281 518 31333 570
rect 31345 518 31397 570
rect 31409 518 31461 570
rect 31473 518 31525 570
rect 16120 348 16172 400
rect 16304 348 16356 400
<< metal2 >>
rect 1122 19816 1178 19825
rect 1122 19751 1178 19760
rect 754 19136 810 19145
rect 754 19071 810 19080
rect 768 18834 796 19071
rect 756 18828 808 18834
rect 756 18770 808 18776
rect 1136 18766 1164 19751
rect 6458 19600 6514 20000
rect 7102 19600 7158 20000
rect 7746 19600 7802 20000
rect 17406 19600 17462 20000
rect 18050 19600 18106 20000
rect 18694 19600 18750 20000
rect 18800 19638 19012 19666
rect 6472 18834 6500 19600
rect 7116 18834 7144 19600
rect 7760 18834 7788 19600
rect 8102 19068 8410 19077
rect 8102 19066 8108 19068
rect 8164 19066 8188 19068
rect 8244 19066 8268 19068
rect 8324 19066 8348 19068
rect 8404 19066 8410 19068
rect 8164 19014 8166 19066
rect 8346 19014 8348 19066
rect 8102 19012 8108 19014
rect 8164 19012 8188 19014
rect 8244 19012 8268 19014
rect 8324 19012 8348 19014
rect 8404 19012 8410 19014
rect 8102 19003 8410 19012
rect 15807 19068 16115 19077
rect 15807 19066 15813 19068
rect 15869 19066 15893 19068
rect 15949 19066 15973 19068
rect 16029 19066 16053 19068
rect 16109 19066 16115 19068
rect 15869 19014 15871 19066
rect 16051 19014 16053 19066
rect 15807 19012 15813 19014
rect 15869 19012 15893 19014
rect 15949 19012 15973 19014
rect 16029 19012 16053 19014
rect 16109 19012 16115 19014
rect 15807 19003 16115 19012
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 1124 18760 1176 18766
rect 1124 18702 1176 18708
rect 848 18624 900 18630
rect 848 18566 900 18572
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 860 18465 888 18566
rect 4250 18524 4558 18533
rect 4250 18522 4256 18524
rect 4312 18522 4336 18524
rect 4392 18522 4416 18524
rect 4472 18522 4496 18524
rect 4552 18522 4558 18524
rect 4312 18470 4314 18522
rect 4494 18470 4496 18522
rect 4250 18468 4256 18470
rect 4312 18468 4336 18470
rect 4392 18468 4416 18470
rect 4472 18468 4496 18470
rect 4552 18468 4558 18470
rect 846 18456 902 18465
rect 4250 18459 4558 18468
rect 846 18391 902 18400
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 848 18216 900 18222
rect 848 18158 900 18164
rect 860 17785 888 18158
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7116 17882 7144 18022
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 846 17776 902 17785
rect 846 17711 902 17720
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 4250 17436 4558 17445
rect 4250 17434 4256 17436
rect 4312 17434 4336 17436
rect 4392 17434 4416 17436
rect 4472 17434 4496 17436
rect 4552 17434 4558 17436
rect 4312 17382 4314 17434
rect 4494 17382 4496 17434
rect 4250 17380 4256 17382
rect 4312 17380 4336 17382
rect 4392 17380 4416 17382
rect 4472 17380 4496 17382
rect 4552 17380 4558 17382
rect 4250 17371 4558 17380
rect 6472 17338 6500 17478
rect 7024 17338 7052 17478
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 6000 17264 6052 17270
rect 6052 17224 6224 17252
rect 6000 17206 6052 17212
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 848 17128 900 17134
rect 846 17096 848 17105
rect 900 17096 902 17105
rect 846 17031 902 17040
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5460 16794 5488 16934
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 16250 1992 16390
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15570 1532 15846
rect 1964 15706 1992 16186
rect 2424 16182 2452 16594
rect 2412 16176 2464 16182
rect 2412 16118 2464 16124
rect 2424 15910 2452 16118
rect 3252 16046 3280 16594
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 3528 16046 3556 16390
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 4172 15910 4200 16390
rect 4250 16348 4558 16357
rect 4250 16346 4256 16348
rect 4312 16346 4336 16348
rect 4392 16346 4416 16348
rect 4472 16346 4496 16348
rect 4552 16346 4558 16348
rect 4312 16294 4314 16346
rect 4494 16294 4496 16346
rect 4250 16292 4256 16294
rect 4312 16292 4336 16294
rect 4392 16292 4416 16294
rect 4472 16292 4496 16294
rect 4552 16292 4558 16294
rect 4250 16283 4558 16292
rect 5644 16046 5672 17138
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5736 16658 5764 16934
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 2700 15706 2728 15846
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 4172 15586 4200 15846
rect 4172 15570 4292 15586
rect 1492 15564 1544 15570
rect 4172 15564 4304 15570
rect 4172 15558 4252 15564
rect 1492 15506 1544 15512
rect 4252 15506 4304 15512
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1780 15162 1808 15302
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1780 14618 1808 15098
rect 2148 14958 2176 15370
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2332 14958 2360 15302
rect 2700 15026 2728 15438
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2240 14618 2268 14758
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1400 14340 1452 14346
rect 1400 14282 1452 14288
rect 1216 13932 1268 13938
rect 1216 13874 1268 13880
rect 1228 13530 1256 13874
rect 1216 13524 1268 13530
rect 1216 13466 1268 13472
rect 1412 13462 1440 14282
rect 1596 14074 1624 14350
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1400 13456 1452 13462
rect 1400 13398 1452 13404
rect 1124 13184 1176 13190
rect 1124 13126 1176 13132
rect 1136 12646 1164 13126
rect 1412 12782 1440 13398
rect 1308 12776 1360 12782
rect 1308 12718 1360 12724
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1124 12640 1176 12646
rect 1124 12582 1176 12588
rect 1136 12434 1164 12582
rect 1044 12406 1164 12434
rect 1044 11558 1072 12406
rect 1320 12170 1348 12718
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1308 12164 1360 12170
rect 1308 12106 1360 12112
rect 1412 11898 1440 12378
rect 1596 12374 1624 14010
rect 2240 13870 2268 14554
rect 2332 14550 2360 14894
rect 2320 14544 2372 14550
rect 2320 14486 2372 14492
rect 2700 14414 2728 14962
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2700 14074 2728 14350
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1688 12782 1716 13262
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1584 12368 1636 12374
rect 1584 12310 1636 12316
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11898 1532 12038
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1492 11892 1544 11898
rect 1492 11834 1544 11840
rect 1032 11552 1084 11558
rect 1032 11494 1084 11500
rect 1044 10674 1072 11494
rect 1412 11218 1440 11834
rect 1596 11694 1624 12310
rect 1688 11762 1716 12718
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1688 11354 1716 11698
rect 1780 11558 1808 13330
rect 3054 13288 3110 13297
rect 3054 13223 3056 13232
rect 3108 13223 3110 13232
rect 3056 13194 3108 13200
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 12345 3096 12582
rect 3054 12336 3110 12345
rect 3054 12271 3110 12280
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10674 1440 11154
rect 1032 10668 1084 10674
rect 1032 10610 1084 10616
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1044 6254 1072 10610
rect 1412 10266 1440 10610
rect 1492 10532 1544 10538
rect 1492 10474 1544 10480
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1308 10192 1360 10198
rect 1308 10134 1360 10140
rect 1216 9920 1268 9926
rect 1216 9862 1268 9868
rect 1228 9586 1256 9862
rect 1216 9580 1268 9586
rect 1216 9522 1268 9528
rect 1032 6248 1084 6254
rect 1032 6190 1084 6196
rect 1216 4684 1268 4690
rect 1216 4626 1268 4632
rect 940 4480 992 4486
rect 940 4422 992 4428
rect 952 4078 980 4422
rect 1228 4282 1256 4626
rect 1216 4276 1268 4282
rect 1216 4218 1268 4224
rect 940 4072 992 4078
rect 940 4014 992 4020
rect 952 3738 980 4014
rect 940 3732 992 3738
rect 940 3674 992 3680
rect 1320 400 1348 10134
rect 1504 10130 1532 10474
rect 1688 10130 1716 11290
rect 1780 10810 1808 11494
rect 3344 11354 3372 11698
rect 3712 11694 3740 12242
rect 3988 12209 4016 13942
rect 4080 13433 4108 15302
rect 4250 15260 4558 15269
rect 4250 15258 4256 15260
rect 4312 15258 4336 15260
rect 4392 15258 4416 15260
rect 4472 15258 4496 15260
rect 4552 15258 4558 15260
rect 4312 15206 4314 15258
rect 4494 15206 4496 15258
rect 4250 15204 4256 15206
rect 4312 15204 4336 15206
rect 4392 15204 4416 15206
rect 4472 15204 4496 15206
rect 4552 15204 4558 15206
rect 4250 15195 4558 15204
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4724 14550 4752 14826
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4250 14172 4558 14181
rect 4250 14170 4256 14172
rect 4312 14170 4336 14172
rect 4392 14170 4416 14172
rect 4472 14170 4496 14172
rect 4552 14170 4558 14172
rect 4312 14118 4314 14170
rect 4494 14118 4496 14170
rect 4250 14116 4256 14118
rect 4312 14116 4336 14118
rect 4392 14116 4416 14118
rect 4472 14116 4496 14118
rect 4552 14116 4558 14118
rect 4250 14107 4558 14116
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 4172 13530 4200 13738
rect 4724 13530 4752 14486
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4908 13870 4936 14214
rect 5000 14074 5028 14214
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5184 13530 5212 13670
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 4066 13424 4122 13433
rect 4066 13359 4122 13368
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4172 12986 4200 13126
rect 4250 13084 4558 13093
rect 4250 13082 4256 13084
rect 4312 13082 4336 13084
rect 4392 13082 4416 13084
rect 4472 13082 4496 13084
rect 4552 13082 4558 13084
rect 4312 13030 4314 13082
rect 4494 13030 4496 13082
rect 4250 13028 4256 13030
rect 4312 13028 4336 13030
rect 4392 13028 4416 13030
rect 4472 13028 4496 13030
rect 4552 13028 4558 13030
rect 4250 13019 4558 13028
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4816 12850 4844 13330
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 3974 12200 4030 12209
rect 4172 12186 4200 12718
rect 5000 12646 5028 13330
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4264 12442 4292 12582
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4540 12186 4568 12242
rect 4172 12158 4660 12186
rect 3974 12135 4030 12144
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4172 11898 4200 12038
rect 4250 11996 4558 12005
rect 4250 11994 4256 11996
rect 4312 11994 4336 11996
rect 4392 11994 4416 11996
rect 4472 11994 4496 11996
rect 4552 11994 4558 11996
rect 4312 11942 4314 11994
rect 4494 11942 4496 11994
rect 4250 11940 4256 11942
rect 4312 11940 4336 11942
rect 4392 11940 4416 11942
rect 4472 11940 4496 11942
rect 4552 11940 4558 11942
rect 4250 11931 4558 11940
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 9722 1624 9862
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1596 9602 1624 9658
rect 1780 9654 1808 10746
rect 2700 10606 2728 10950
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 1768 9648 1820 9654
rect 1596 9574 1716 9602
rect 1768 9590 1820 9596
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1412 9178 1440 9318
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1412 8498 1440 9114
rect 1688 9042 1716 9574
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 2148 9178 2176 9318
rect 3252 9178 3280 9318
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 1596 8634 1624 8910
rect 2424 8634 2452 8910
rect 2608 8634 2636 8978
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 7274 1440 8434
rect 2424 7970 2452 8570
rect 2424 7954 2544 7970
rect 2424 7948 2556 7954
rect 2424 7942 2504 7948
rect 2504 7890 2556 7896
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1964 7342 1992 7822
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1400 7268 1452 7274
rect 1400 7210 1452 7216
rect 1964 6866 1992 7278
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5030 1440 5714
rect 2240 5370 2268 6802
rect 3528 6662 3556 10474
rect 3620 10198 3648 11154
rect 3712 10198 3740 11630
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4264 11354 4292 11494
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4250 10908 4558 10917
rect 4250 10906 4256 10908
rect 4312 10906 4336 10908
rect 4392 10906 4416 10908
rect 4472 10906 4496 10908
rect 4552 10906 4558 10908
rect 4312 10854 4314 10906
rect 4494 10854 4496 10906
rect 4250 10852 4256 10854
rect 4312 10852 4336 10854
rect 4392 10852 4416 10854
rect 4472 10852 4496 10854
rect 4552 10852 4558 10854
rect 4250 10843 4558 10852
rect 4632 10690 4660 12158
rect 4540 10662 4660 10690
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3620 9518 3648 10134
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3804 9722 3832 10066
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9722 4108 9998
rect 4172 9994 4200 10406
rect 4264 10198 4292 10542
rect 4540 10470 4568 10662
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 4250 9820 4558 9829
rect 4250 9818 4256 9820
rect 4312 9818 4336 9820
rect 4392 9818 4416 9820
rect 4472 9818 4496 9820
rect 4552 9818 4558 9820
rect 4312 9766 4314 9818
rect 4494 9766 4496 9818
rect 4250 9764 4256 9766
rect 4312 9764 4336 9766
rect 4392 9764 4416 9766
rect 4472 9764 4496 9766
rect 4552 9764 4558 9766
rect 4250 9755 4558 9764
rect 4724 9722 4752 10066
rect 5000 9994 5028 12582
rect 5368 12434 5396 14554
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 13326 5488 13806
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5828 12434 5856 15302
rect 5998 14920 6054 14929
rect 5998 14855 6054 14864
rect 6092 14884 6144 14890
rect 6012 14822 6040 14855
rect 6092 14826 6144 14832
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5920 14074 5948 14418
rect 6104 14278 6132 14826
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6104 14006 6132 14214
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6104 12782 6132 13942
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 5368 12406 5488 12434
rect 5828 12406 6040 12434
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5276 11218 5304 11834
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5276 10810 5304 11154
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5460 10742 5488 12406
rect 6012 11694 6040 12406
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5644 10810 5672 11630
rect 6104 11354 6132 11766
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6196 11286 6224 17224
rect 6472 17218 6500 17274
rect 6472 17190 6592 17218
rect 6564 16794 6592 17190
rect 7392 17134 7420 18226
rect 7760 17746 7788 18226
rect 7944 18222 7972 18566
rect 8496 18222 8524 18566
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7944 17746 7972 18022
rect 8102 17980 8410 17989
rect 8102 17978 8108 17980
rect 8164 17978 8188 17980
rect 8244 17978 8268 17980
rect 8324 17978 8348 17980
rect 8404 17978 8410 17980
rect 8164 17926 8166 17978
rect 8346 17926 8348 17978
rect 8102 17924 8108 17926
rect 8164 17924 8188 17926
rect 8244 17924 8268 17926
rect 8324 17924 8348 17926
rect 8404 17924 8410 17926
rect 8102 17915 8410 17924
rect 8588 17814 8616 18294
rect 8956 18222 8984 18566
rect 9508 18426 9536 18770
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17134 7972 17478
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6460 16720 6512 16726
rect 6460 16662 6512 16668
rect 6472 16046 6500 16662
rect 7944 16640 7972 17070
rect 8036 16794 8064 17614
rect 9232 17066 9260 18022
rect 9784 17134 9812 18226
rect 9876 18222 9904 18566
rect 10152 18426 10180 18770
rect 10520 18442 10548 18770
rect 10520 18426 10640 18442
rect 10140 18420 10192 18426
rect 10520 18420 10652 18426
rect 10520 18414 10600 18420
rect 10140 18362 10192 18368
rect 10600 18362 10652 18368
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 10152 18136 10180 18362
rect 10324 18148 10376 18154
rect 10152 18108 10324 18136
rect 10324 18090 10376 18096
rect 10796 17134 10824 18770
rect 11440 18358 11468 18770
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 11955 18524 12263 18533
rect 11955 18522 11961 18524
rect 12017 18522 12041 18524
rect 12097 18522 12121 18524
rect 12177 18522 12201 18524
rect 12257 18522 12263 18524
rect 12017 18470 12019 18522
rect 12199 18470 12201 18522
rect 11955 18468 11961 18470
rect 12017 18468 12041 18470
rect 12097 18468 12121 18470
rect 12177 18468 12201 18470
rect 12257 18468 12263 18470
rect 11955 18459 12263 18468
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8102 16892 8410 16901
rect 8102 16890 8108 16892
rect 8164 16890 8188 16892
rect 8244 16890 8268 16892
rect 8324 16890 8348 16892
rect 8404 16890 8410 16892
rect 8164 16838 8166 16890
rect 8346 16838 8348 16890
rect 8102 16836 8108 16838
rect 8164 16836 8188 16838
rect 8244 16836 8268 16838
rect 8324 16836 8348 16838
rect 8404 16836 8410 16838
rect 8102 16827 8410 16836
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8116 16652 8168 16658
rect 7944 16612 8116 16640
rect 8116 16594 8168 16600
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6288 13938 6316 14350
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6380 12434 6408 15846
rect 6472 15570 6500 15982
rect 6564 15638 6592 16390
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6472 15026 6500 15506
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 6460 15020 6512 15026
rect 6460 14962 6512 14968
rect 6472 14482 6500 14962
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6932 13870 6960 14010
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7300 12986 7328 13194
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 6826 12880 6882 12889
rect 6826 12815 6882 12824
rect 6840 12442 6868 12815
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 7116 12442 7144 12650
rect 6828 12436 6880 12442
rect 6380 12406 6592 12434
rect 6564 12374 6592 12406
rect 6828 12378 6880 12384
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6458 12200 6514 12209
rect 6458 12135 6514 12144
rect 6274 11656 6330 11665
rect 6274 11591 6330 11600
rect 6288 11558 6316 11591
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6472 11354 6500 12135
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 5000 9518 5028 9930
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 3620 9178 3648 9454
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3804 8974 3832 9454
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3712 7954 3740 8230
rect 3804 8022 3832 8910
rect 4172 8838 4200 9318
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 8294 4200 8774
rect 4250 8732 4558 8741
rect 4250 8730 4256 8732
rect 4312 8730 4336 8732
rect 4392 8730 4416 8732
rect 4472 8730 4496 8732
rect 4552 8730 4558 8732
rect 4312 8678 4314 8730
rect 4494 8678 4496 8730
rect 4250 8676 4256 8678
rect 4312 8676 4336 8678
rect 4392 8676 4416 8678
rect 4472 8676 4496 8678
rect 4552 8676 4558 8678
rect 4250 8667 4558 8676
rect 5736 8634 5764 11154
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6288 9178 6316 9318
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6656 9110 6684 11562
rect 6840 11558 6868 12242
rect 6932 11830 6960 12310
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11218 6868 11494
rect 7024 11354 7052 12174
rect 7208 12170 7236 12650
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 7116 10538 7144 12038
rect 7208 11014 7236 12106
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7208 10606 7236 10950
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7116 9518 7144 10474
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 9110 6776 9318
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8634 7052 8774
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7392 8537 7420 15302
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7484 12986 7512 13670
rect 7576 13394 7604 13874
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7668 13326 7696 13806
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7484 12374 7512 12582
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7484 10198 7512 12310
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7484 9518 7512 10134
rect 7576 10010 7604 13126
rect 7668 12782 7696 13262
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7760 12434 7788 16390
rect 8404 16114 8432 16662
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8404 15892 8432 16050
rect 8496 16046 8524 16934
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8404 15864 8524 15892
rect 8102 15804 8410 15813
rect 8102 15802 8108 15804
rect 8164 15802 8188 15804
rect 8244 15802 8268 15804
rect 8324 15802 8348 15804
rect 8404 15802 8410 15804
rect 8164 15750 8166 15802
rect 8346 15750 8348 15802
rect 8102 15748 8108 15750
rect 8164 15748 8188 15750
rect 8244 15748 8268 15750
rect 8324 15748 8348 15750
rect 8404 15748 8410 15750
rect 8102 15739 8410 15748
rect 8208 15088 8260 15094
rect 8206 15056 8208 15065
rect 8260 15056 8262 15065
rect 8206 14991 8262 15000
rect 8102 14716 8410 14725
rect 8102 14714 8108 14716
rect 8164 14714 8188 14716
rect 8244 14714 8268 14716
rect 8324 14714 8348 14716
rect 8404 14714 8410 14716
rect 8164 14662 8166 14714
rect 8346 14662 8348 14714
rect 8102 14660 8108 14662
rect 8164 14660 8188 14662
rect 8244 14660 8268 14662
rect 8324 14660 8348 14662
rect 8404 14660 8410 14662
rect 8102 14651 8410 14660
rect 8496 14532 8524 15864
rect 8404 14504 8524 14532
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7852 13870 7880 14010
rect 8404 13938 8432 14504
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 8036 13530 8064 13874
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 8102 13628 8410 13637
rect 8102 13626 8108 13628
rect 8164 13626 8188 13628
rect 8244 13626 8268 13628
rect 8324 13626 8348 13628
rect 8404 13626 8410 13628
rect 8164 13574 8166 13626
rect 8346 13574 8348 13626
rect 8102 13572 8108 13574
rect 8164 13572 8188 13574
rect 8244 13572 8268 13574
rect 8324 13572 8348 13574
rect 8404 13572 8410 13574
rect 8102 13563 8410 13572
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8496 13394 8524 13738
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9324 13190 9352 13262
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12986 9352 13126
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7760 12406 7880 12434
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7760 11898 7788 12310
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7656 11824 7708 11830
rect 7708 11772 7788 11778
rect 7656 11766 7788 11772
rect 7668 11750 7788 11766
rect 7760 11626 7788 11750
rect 7852 11694 7880 12406
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7760 10742 7788 11562
rect 7944 10826 7972 12786
rect 9220 12776 9272 12782
rect 9140 12736 9220 12764
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8036 12442 8064 12582
rect 8102 12540 8410 12549
rect 8102 12538 8108 12540
rect 8164 12538 8188 12540
rect 8244 12538 8268 12540
rect 8324 12538 8348 12540
rect 8404 12538 8410 12540
rect 8164 12486 8166 12538
rect 8346 12486 8348 12538
rect 8102 12484 8108 12486
rect 8164 12484 8188 12486
rect 8244 12484 8268 12486
rect 8324 12484 8348 12486
rect 8404 12484 8410 12486
rect 8102 12475 8410 12484
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 9140 12306 9168 12736
rect 9220 12718 9272 12724
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11694 8064 12038
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8114 11656 8170 11665
rect 8114 11591 8170 11600
rect 8128 11558 8156 11591
rect 9140 11558 9168 12242
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8102 11452 8410 11461
rect 8102 11450 8108 11452
rect 8164 11450 8188 11452
rect 8244 11450 8268 11452
rect 8324 11450 8348 11452
rect 8404 11450 8410 11452
rect 8164 11398 8166 11450
rect 8346 11398 8348 11450
rect 8102 11396 8108 11398
rect 8164 11396 8188 11398
rect 8244 11396 8268 11398
rect 8324 11396 8348 11398
rect 8404 11396 8410 11398
rect 8102 11387 8410 11396
rect 8300 11280 8352 11286
rect 8496 11234 8524 11494
rect 8352 11228 8524 11234
rect 8300 11222 8524 11228
rect 8116 11212 8168 11218
rect 8312 11206 8524 11222
rect 8116 11154 8168 11160
rect 7852 10798 7972 10826
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7760 10130 7788 10542
rect 7852 10198 7880 10798
rect 7930 10704 7986 10713
rect 7930 10639 7986 10648
rect 7944 10470 7972 10639
rect 8128 10520 8156 11154
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8588 10606 8616 11086
rect 9140 10606 9168 11494
rect 9416 11014 9444 16390
rect 10152 16114 10180 16594
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10244 16114 10272 16390
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10152 15706 10180 16050
rect 10244 15706 10272 16050
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10704 15570 10732 15982
rect 10796 15638 10824 17070
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11440 16454 11468 16594
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11072 16250 11100 16390
rect 11440 16250 11468 16390
rect 11624 16250 11652 18022
rect 12268 17882 12296 18158
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 11955 17436 12263 17445
rect 11955 17434 11961 17436
rect 12017 17434 12041 17436
rect 12097 17434 12121 17436
rect 12177 17434 12201 17436
rect 12257 17434 12263 17436
rect 12017 17382 12019 17434
rect 12199 17382 12201 17434
rect 11955 17380 11961 17382
rect 12017 17380 12041 17382
rect 12097 17380 12121 17382
rect 12177 17380 12201 17382
rect 12257 17380 12263 17382
rect 11955 17371 12263 17380
rect 12360 17338 12388 17682
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 10876 16176 10928 16182
rect 10876 16118 10928 16124
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 9508 15162 9536 15506
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9692 14822 9720 15506
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14618 9720 14758
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9784 13326 9812 14418
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 13530 9904 14350
rect 9968 14260 9996 14894
rect 10152 14890 10180 15506
rect 10704 15434 10732 15506
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10796 14958 10824 15574
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10520 14618 10548 14826
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10140 14272 10192 14278
rect 9968 14232 10140 14260
rect 10140 14214 10192 14220
rect 10152 13802 10180 14214
rect 10796 13802 10824 14894
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9692 12442 9720 12718
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9784 12306 9812 13262
rect 9876 12714 9904 13466
rect 10060 12986 10088 13670
rect 10152 13530 10180 13738
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 10060 12628 10088 12922
rect 10888 12753 10916 16118
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11072 14482 11100 14894
rect 11256 14482 11284 15506
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11716 14362 11744 16934
rect 11900 16794 11928 17070
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11796 16652 11848 16658
rect 12176 16640 12204 17070
rect 12452 16794 12480 17070
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12348 16652 12400 16658
rect 12176 16612 12348 16640
rect 11796 16594 11848 16600
rect 12348 16594 12400 16600
rect 11808 16522 11836 16594
rect 11796 16516 11848 16522
rect 11796 16458 11848 16464
rect 11808 15910 11836 16458
rect 11955 16348 12263 16357
rect 11955 16346 11961 16348
rect 12017 16346 12041 16348
rect 12097 16346 12121 16348
rect 12177 16346 12201 16348
rect 12257 16346 12263 16348
rect 12017 16294 12019 16346
rect 12199 16294 12201 16346
rect 11955 16292 11961 16294
rect 12017 16292 12041 16294
rect 12097 16292 12121 16294
rect 12177 16292 12201 16294
rect 12257 16292 12263 16294
rect 11955 16283 12263 16292
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11808 15706 11836 15846
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11900 15638 11928 15982
rect 12360 15978 12388 16594
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 11955 15260 12263 15269
rect 11955 15258 11961 15260
rect 12017 15258 12041 15260
rect 12097 15258 12121 15260
rect 12177 15258 12201 15260
rect 12257 15258 12263 15260
rect 12017 15206 12019 15258
rect 12199 15206 12201 15258
rect 11955 15204 11961 15206
rect 12017 15204 12041 15206
rect 12097 15204 12121 15206
rect 12177 15204 12201 15206
rect 12257 15204 12263 15206
rect 11955 15195 12263 15204
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11716 14334 11836 14362
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 13870 11744 14214
rect 11704 13864 11756 13870
rect 11624 13812 11704 13818
rect 11624 13806 11756 13812
rect 11624 13790 11744 13806
rect 11244 13728 11296 13734
rect 11242 13696 11244 13705
rect 11520 13728 11572 13734
rect 11296 13696 11298 13705
rect 11520 13670 11572 13676
rect 11242 13631 11298 13640
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10874 12744 10930 12753
rect 10874 12679 10930 12688
rect 9968 12600 10088 12628
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9600 11898 9628 12242
rect 9876 11914 9904 12242
rect 9784 11898 9904 11914
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9772 11892 9904 11898
rect 9824 11886 9904 11892
rect 9772 11834 9824 11840
rect 9968 11694 9996 12600
rect 10046 12472 10102 12481
rect 10046 12407 10102 12416
rect 10060 12374 10088 12407
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 10980 12238 11008 12786
rect 11532 12442 11560 13670
rect 11624 13530 11652 13790
rect 11808 13569 11836 14334
rect 11900 14226 11928 14894
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 11880 14198 11928 14226
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 11880 14090 11908 14198
rect 11955 14172 12263 14181
rect 11955 14170 11961 14172
rect 12017 14170 12041 14172
rect 12097 14170 12121 14172
rect 12177 14170 12201 14172
rect 12257 14170 12263 14172
rect 12017 14118 12019 14170
rect 12199 14118 12201 14170
rect 11955 14116 11961 14118
rect 12017 14116 12041 14118
rect 12097 14116 12121 14118
rect 12177 14116 12201 14118
rect 12257 14116 12263 14118
rect 11955 14107 12263 14116
rect 11880 14062 11928 14090
rect 11900 14056 11928 14062
rect 11900 14028 12112 14056
rect 11794 13560 11850 13569
rect 11612 13524 11664 13530
rect 11794 13495 11850 13504
rect 11612 13466 11664 13472
rect 12084 13326 12112 14028
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12176 13394 12204 13738
rect 12360 13530 12388 14214
rect 12452 13938 12480 14350
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12164 13388 12216 13394
rect 12216 13348 12388 13376
rect 12164 13330 12216 13336
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9508 11082 9536 11630
rect 9784 11150 9812 11630
rect 10244 11626 10272 12174
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 9772 11144 9824 11150
rect 9678 11112 9734 11121
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9588 11076 9640 11082
rect 9772 11086 9824 11092
rect 10140 11144 10192 11150
rect 10192 11092 10272 11098
rect 10140 11086 10272 11092
rect 10152 11070 10272 11086
rect 9678 11047 9734 11056
rect 9588 11018 9640 11024
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9508 10810 9536 11018
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 8036 10492 8156 10520
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7840 10192 7892 10198
rect 7840 10134 7892 10140
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7576 9982 7788 10010
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 9518 7604 9862
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 9042 7696 9318
rect 7760 9081 7788 9982
rect 7852 9518 7880 10134
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7852 9110 7880 9318
rect 7840 9104 7892 9110
rect 7746 9072 7802 9081
rect 7656 9036 7708 9042
rect 7840 9046 7892 9052
rect 7746 9007 7802 9016
rect 7656 8978 7708 8984
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7378 8528 7434 8537
rect 7378 8463 7434 8472
rect 7484 8430 7512 8910
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 8498 7880 8774
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 5736 8022 5764 8298
rect 6380 8090 6408 8366
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5736 7750 5764 7822
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 4250 7644 4558 7653
rect 4250 7642 4256 7644
rect 4312 7642 4336 7644
rect 4392 7642 4416 7644
rect 4472 7642 4496 7644
rect 4552 7642 4558 7644
rect 4312 7590 4314 7642
rect 4494 7590 4496 7642
rect 4250 7588 4256 7590
rect 4312 7588 4336 7590
rect 4392 7588 4416 7590
rect 4472 7588 4496 7590
rect 4552 7588 4558 7590
rect 4250 7579 4558 7588
rect 5644 7274 5672 7686
rect 6104 7342 6132 7890
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 7002 5580 7142
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5644 6934 5672 7210
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5642 2452 6054
rect 2608 5914 2636 6190
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2412 5636 2464 5642
rect 2412 5578 2464 5584
rect 2424 5370 2452 5578
rect 2608 5370 2636 5850
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1412 4826 1440 4966
rect 1688 4826 1716 5102
rect 1964 4826 1992 5102
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4282 1532 4422
rect 2240 4298 2268 5306
rect 2700 4758 2728 5782
rect 2976 5778 3004 6258
rect 3620 6254 3648 6598
rect 4250 6556 4558 6565
rect 4250 6554 4256 6556
rect 4312 6554 4336 6556
rect 4392 6554 4416 6556
rect 4472 6554 4496 6556
rect 4552 6554 4558 6556
rect 4312 6502 4314 6554
rect 4494 6502 4496 6554
rect 4250 6500 4256 6502
rect 4312 6500 4336 6502
rect 4392 6500 4416 6502
rect 4472 6500 4496 6502
rect 4552 6500 4558 6502
rect 4250 6491 4558 6500
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 4436 6248 4488 6254
rect 5080 6248 5132 6254
rect 4436 6190 4488 6196
rect 4618 6216 4674 6225
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 3068 5574 3096 6190
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 3160 5778 3188 6054
rect 4172 5846 4200 6054
rect 4448 5914 4476 6190
rect 5080 6190 5132 6196
rect 4618 6151 4674 6160
rect 4896 6180 4948 6186
rect 4632 5914 4660 6151
rect 4896 6122 4948 6128
rect 4908 5914 4936 6122
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 4826 3096 5510
rect 3160 5166 3188 5714
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3528 5098 3556 5714
rect 4172 5166 4200 5782
rect 4250 5468 4558 5477
rect 4250 5466 4256 5468
rect 4312 5466 4336 5468
rect 4392 5466 4416 5468
rect 4472 5466 4496 5468
rect 4552 5466 4558 5468
rect 4312 5414 4314 5466
rect 4494 5414 4496 5466
rect 4250 5412 4256 5414
rect 4312 5412 4336 5414
rect 4392 5412 4416 5414
rect 4472 5412 4496 5414
rect 4552 5412 4558 5414
rect 4250 5403 4558 5412
rect 4908 5302 4936 5850
rect 5092 5778 5120 6190
rect 5736 5778 5764 7278
rect 6012 6458 6040 7278
rect 6196 6866 6224 7414
rect 6288 7342 6316 7686
rect 6276 7336 6328 7342
rect 6380 7324 6408 8026
rect 7392 8022 7420 8230
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6564 7426 6592 7822
rect 6564 7410 6776 7426
rect 6552 7404 6788 7410
rect 6604 7398 6736 7404
rect 6552 7346 6604 7352
rect 6736 7346 6788 7352
rect 6460 7336 6512 7342
rect 6380 7296 6460 7324
rect 6276 7278 6328 7284
rect 6460 7278 6512 7284
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6934 6592 7142
rect 7208 6934 7236 7210
rect 7300 6934 7328 7890
rect 7852 7886 7880 8230
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 8036 7478 8064 10492
rect 8102 10364 8410 10373
rect 8102 10362 8108 10364
rect 8164 10362 8188 10364
rect 8244 10362 8268 10364
rect 8324 10362 8348 10364
rect 8404 10362 8410 10364
rect 8164 10310 8166 10362
rect 8346 10310 8348 10362
rect 8102 10308 8108 10310
rect 8164 10308 8188 10310
rect 8244 10308 8268 10310
rect 8324 10308 8348 10310
rect 8404 10308 8410 10310
rect 8102 10299 8410 10308
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8102 9276 8410 9285
rect 8102 9274 8108 9276
rect 8164 9274 8188 9276
rect 8244 9274 8268 9276
rect 8324 9274 8348 9276
rect 8404 9274 8410 9276
rect 8164 9222 8166 9274
rect 8346 9222 8348 9274
rect 8102 9220 8108 9222
rect 8164 9220 8188 9222
rect 8244 9220 8268 9222
rect 8324 9220 8348 9222
rect 8404 9220 8410 9222
rect 8102 9211 8410 9220
rect 8496 9160 8524 9318
rect 8404 9132 8524 9160
rect 8404 8838 8432 9132
rect 8588 8838 8616 10542
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8680 10062 8708 10474
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8772 9722 8800 10406
rect 9508 10180 9536 10746
rect 9600 10606 9628 11018
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9588 10192 9640 10198
rect 9508 10152 9588 10180
rect 9588 10134 9640 10140
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8404 8430 8432 8774
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8102 8188 8410 8197
rect 8102 8186 8108 8188
rect 8164 8186 8188 8188
rect 8244 8186 8268 8188
rect 8324 8186 8348 8188
rect 8404 8186 8410 8188
rect 8164 8134 8166 8186
rect 8346 8134 8348 8186
rect 8102 8132 8108 8134
rect 8164 8132 8188 8134
rect 8244 8132 8268 8134
rect 8324 8132 8348 8134
rect 8404 8132 8410 8134
rect 8102 8123 8410 8132
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8864 7886 8892 8026
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 8036 6934 8064 7210
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8102 7100 8410 7109
rect 8102 7098 8108 7100
rect 8164 7098 8188 7100
rect 8244 7098 8268 7100
rect 8324 7098 8348 7100
rect 8404 7098 8410 7100
rect 8164 7046 8166 7098
rect 8346 7046 8348 7098
rect 8102 7044 8108 7046
rect 8164 7044 8188 7046
rect 8244 7044 8268 7046
rect 8324 7044 8348 7046
rect 8404 7044 8410 7046
rect 8102 7035 8410 7044
rect 8680 7002 8708 7142
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7288 6928 7340 6934
rect 8024 6928 8076 6934
rect 7288 6870 7340 6876
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6000 6452 6052 6458
rect 6196 6440 6224 6802
rect 6276 6452 6328 6458
rect 6196 6412 6276 6440
rect 6000 6394 6052 6400
rect 6276 6394 6328 6400
rect 6564 6254 6592 6870
rect 7484 6866 7788 6882
rect 8024 6870 8076 6876
rect 8680 6866 8708 6938
rect 7472 6860 7800 6866
rect 7524 6854 7748 6860
rect 7472 6802 7524 6808
rect 7748 6802 7800 6808
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5000 5370 5028 5714
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 5092 5302 5120 5714
rect 5460 5370 5488 5714
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 3516 5092 3568 5098
rect 3516 5034 3568 5040
rect 5092 5030 5120 5238
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 6932 4758 6960 6734
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 6458 8524 6598
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8772 6322 8800 7346
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8864 6254 8892 6666
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8956 6254 8984 6598
rect 9692 6338 9720 11047
rect 10244 11014 10272 11070
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10060 10441 10088 10950
rect 10152 10674 10180 10950
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10244 10470 10272 10950
rect 10796 10606 10824 11154
rect 10784 10600 10836 10606
rect 11256 10577 11284 11494
rect 11336 11280 11388 11286
rect 11440 11268 11468 11562
rect 11532 11558 11560 12378
rect 11624 12170 11652 13126
rect 11808 12986 11836 13126
rect 11955 13084 12263 13093
rect 11955 13082 11961 13084
rect 12017 13082 12041 13084
rect 12097 13082 12121 13084
rect 12177 13082 12201 13084
rect 12257 13082 12263 13084
rect 12017 13030 12019 13082
rect 12199 13030 12201 13082
rect 11955 13028 11961 13030
rect 12017 13028 12041 13030
rect 12097 13028 12121 13030
rect 12177 13028 12201 13030
rect 12257 13028 12263 13030
rect 11955 13019 12263 13028
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 11888 12436 11940 12442
rect 11992 12434 12020 12582
rect 11992 12406 12112 12434
rect 11888 12378 11940 12384
rect 11900 12306 11928 12378
rect 12084 12374 12112 12406
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11388 11240 11468 11268
rect 11336 11222 11388 11228
rect 10784 10542 10836 10548
rect 11242 10568 11298 10577
rect 11242 10503 11298 10512
rect 10232 10464 10284 10470
rect 10046 10432 10102 10441
rect 10232 10406 10284 10412
rect 10046 10367 10102 10376
rect 10244 8362 10272 10406
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10980 8430 11008 9454
rect 11348 9382 11376 11222
rect 11532 11218 11560 11494
rect 11624 11286 11652 12106
rect 11900 12050 11928 12242
rect 12176 12084 12204 12582
rect 12268 12442 12296 12582
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12360 12152 12388 13348
rect 12452 12782 12480 13874
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12360 12124 12480 12152
rect 12176 12056 12388 12084
rect 11880 12022 11928 12050
rect 11880 11914 11908 12022
rect 11955 11996 12263 12005
rect 11955 11994 11961 11996
rect 12017 11994 12041 11996
rect 12097 11994 12121 11996
rect 12177 11994 12201 11996
rect 12257 11994 12263 11996
rect 12017 11942 12019 11994
rect 12199 11942 12201 11994
rect 11955 11940 11961 11942
rect 12017 11940 12041 11942
rect 12097 11940 12121 11942
rect 12177 11940 12201 11942
rect 12257 11940 12263 11942
rect 11955 11931 12263 11940
rect 11880 11886 11928 11914
rect 11900 11694 11928 11886
rect 11980 11824 12032 11830
rect 12032 11784 12112 11812
rect 11980 11766 12032 11772
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11808 11506 11836 11630
rect 11992 11529 12020 11630
rect 11978 11520 12034 11529
rect 11808 11478 11978 11506
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11624 9518 11652 11222
rect 11808 10130 11836 11478
rect 11978 11455 12034 11464
rect 12084 11014 12112 11784
rect 11888 11008 11940 11014
rect 11880 10956 11888 10962
rect 11880 10950 11940 10956
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 11880 10934 11928 10950
rect 11880 10826 11908 10934
rect 11955 10908 12263 10917
rect 11955 10906 11961 10908
rect 12017 10906 12041 10908
rect 12097 10906 12121 10908
rect 12177 10906 12201 10908
rect 12257 10906 12263 10908
rect 12017 10854 12019 10906
rect 12199 10854 12201 10906
rect 11955 10852 11961 10854
rect 12017 10852 12041 10854
rect 12097 10852 12121 10854
rect 12177 10852 12201 10854
rect 12257 10852 12263 10854
rect 11955 10843 12263 10852
rect 11880 10798 11928 10826
rect 11900 10606 11928 10798
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11796 10124 11848 10130
rect 11900 10112 11928 10542
rect 11980 10124 12032 10130
rect 11900 10084 11980 10112
rect 11796 10066 11848 10072
rect 11980 10066 12032 10072
rect 11955 9820 12263 9829
rect 11955 9818 11961 9820
rect 12017 9818 12041 9820
rect 12097 9818 12121 9820
rect 12177 9818 12201 9820
rect 12257 9818 12263 9820
rect 12017 9766 12019 9818
rect 12199 9766 12201 9818
rect 11955 9764 11961 9766
rect 12017 9764 12041 9766
rect 12097 9764 12121 9766
rect 12177 9764 12201 9766
rect 12257 9764 12263 9766
rect 11955 9755 12263 9764
rect 12360 9674 12388 12056
rect 12452 9897 12480 12124
rect 12544 10538 12572 18566
rect 13648 18340 13676 18702
rect 14200 18426 14228 18770
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14004 18352 14056 18358
rect 13648 18312 14004 18340
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 13004 17882 13032 18158
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13372 17882 13400 18022
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 12820 17746 12940 17762
rect 13648 17746 13676 18312
rect 14004 18294 14056 18300
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13740 17882 13768 18158
rect 15028 18057 15056 18566
rect 16224 18222 16252 18770
rect 16960 18222 16988 18770
rect 17420 18714 17448 19600
rect 17868 18760 17920 18766
rect 17420 18686 17632 18714
rect 17868 18702 17920 18708
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 15014 18048 15070 18057
rect 15014 17983 15070 17992
rect 15807 17980 16115 17989
rect 15807 17978 15813 17980
rect 15869 17978 15893 17980
rect 15949 17978 15973 17980
rect 16029 17978 16053 17980
rect 16109 17978 16115 17980
rect 15869 17926 15871 17978
rect 16051 17926 16053 17978
rect 15807 17924 15813 17926
rect 15869 17924 15893 17926
rect 15949 17924 15973 17926
rect 16029 17924 16053 17926
rect 16109 17924 16115 17926
rect 15807 17915 16115 17924
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 16224 17746 16252 18158
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 12820 17740 12952 17746
rect 12820 17734 12900 17740
rect 12820 17270 12848 17734
rect 12900 17682 12952 17688
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 13004 17626 13032 17682
rect 12912 17598 13032 17626
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12912 16998 12940 17598
rect 13648 17202 13676 17682
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16794 12940 16934
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 13648 16726 13676 17138
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12636 16046 12664 16526
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12636 15706 12664 15982
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12820 13258 12848 13670
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12636 10538 12664 12378
rect 12912 12322 12940 15302
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13096 14482 13124 14962
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13280 14074 13308 14214
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13372 13870 13400 14350
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 13004 12434 13032 13398
rect 13096 13258 13124 13670
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 13188 12986 13216 13670
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13096 12434 13124 12582
rect 13004 12406 13124 12434
rect 13096 12374 13124 12406
rect 12992 12368 13044 12374
rect 12912 12316 12992 12322
rect 12912 12310 13044 12316
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 12912 12294 13032 12310
rect 13096 12220 13124 12310
rect 12820 12192 13124 12220
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12438 9888 12494 9897
rect 12438 9823 12494 9832
rect 12268 9646 12388 9674
rect 12268 9586 12296 9646
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10336 6662 10364 7890
rect 10980 7886 11008 8366
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10980 7274 11008 7822
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 7274 11284 7686
rect 11532 7546 11560 8774
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9600 6310 9720 6338
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 8102 6012 8410 6021
rect 8102 6010 8108 6012
rect 8164 6010 8188 6012
rect 8244 6010 8268 6012
rect 8324 6010 8348 6012
rect 8404 6010 8410 6012
rect 8164 5958 8166 6010
rect 8346 5958 8348 6010
rect 8102 5956 8108 5958
rect 8164 5956 8188 5958
rect 8244 5956 8268 5958
rect 8324 5956 8348 5958
rect 8404 5956 8410 5958
rect 8102 5947 8410 5956
rect 8956 5914 8984 6054
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 5166 7328 5510
rect 7760 5302 7788 5714
rect 8220 5302 8248 5714
rect 9048 5574 9076 6054
rect 9600 5914 9628 6310
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9692 5778 9720 6122
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9218 5400 9274 5409
rect 9218 5335 9220 5344
rect 9272 5335 9274 5344
rect 9220 5306 9272 5312
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7760 5030 7788 5238
rect 9324 5166 9352 5510
rect 9508 5302 9536 5578
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 6920 4752 6972 4758
rect 7208 4729 7236 4762
rect 7392 4758 7420 4966
rect 8102 4924 8410 4933
rect 8102 4922 8108 4924
rect 8164 4922 8188 4924
rect 8244 4922 8268 4924
rect 8324 4922 8348 4924
rect 8404 4922 8410 4924
rect 8164 4870 8166 4922
rect 8346 4870 8348 4922
rect 8102 4868 8108 4870
rect 8164 4868 8188 4870
rect 8244 4868 8268 4870
rect 8324 4868 8348 4870
rect 8404 4868 8410 4870
rect 8102 4859 8410 4868
rect 7380 4752 7432 4758
rect 6920 4694 6972 4700
rect 7194 4720 7250 4729
rect 7380 4694 7432 4700
rect 7194 4655 7250 4664
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 3516 4616 3568 4622
rect 7288 4616 7340 4622
rect 3516 4558 3568 4564
rect 4894 4584 4950 4593
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 1492 4276 1544 4282
rect 1492 4218 1544 4224
rect 1872 4270 2268 4298
rect 3436 4282 3464 4422
rect 1872 4078 1900 4270
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 1964 4078 1992 4150
rect 2240 4078 2268 4270
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 1872 2990 1900 3674
rect 2056 3602 2084 3878
rect 2332 3602 2360 4082
rect 3528 4078 3556 4558
rect 7288 4558 7340 4564
rect 4894 4519 4896 4528
rect 4948 4519 4950 4528
rect 4896 4490 4948 4496
rect 4250 4380 4558 4389
rect 4250 4378 4256 4380
rect 4312 4378 4336 4380
rect 4392 4378 4416 4380
rect 4472 4378 4496 4380
rect 4552 4378 4558 4380
rect 4312 4326 4314 4378
rect 4494 4326 4496 4378
rect 4250 4324 4256 4326
rect 4312 4324 4336 4326
rect 4392 4324 4416 4326
rect 4472 4324 4496 4326
rect 4552 4324 4558 4326
rect 4250 4315 4558 4324
rect 7300 4078 7328 4558
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2516 3738 2544 3946
rect 3528 3738 3556 4014
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 2148 2990 2176 3470
rect 2516 2990 2544 3674
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3068 3398 3096 3538
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3068 3194 3096 3334
rect 4250 3292 4558 3301
rect 4250 3290 4256 3292
rect 4312 3290 4336 3292
rect 4392 3290 4416 3292
rect 4472 3290 4496 3292
rect 4552 3290 4558 3292
rect 4312 3238 4314 3290
rect 4494 3238 4496 3290
rect 4250 3236 4256 3238
rect 4312 3236 4336 3238
rect 4392 3236 4416 3238
rect 4472 3236 4496 3238
rect 4552 3236 4558 3238
rect 4250 3227 4558 3236
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2412 2848 2464 2854
rect 2412 2790 2464 2796
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2424 2650 2452 2790
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2700 2582 2728 2790
rect 3068 2774 3096 3130
rect 5460 3074 5488 3946
rect 7300 3670 7328 4014
rect 9140 3942 9168 4626
rect 9324 4078 9352 5102
rect 9508 4758 9536 5238
rect 9784 5166 9812 6394
rect 10336 6254 10364 6598
rect 10520 6458 10548 6802
rect 10980 6798 11008 7210
rect 11624 7206 11652 8978
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10980 6322 11008 6734
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5914 10364 6054
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9968 5370 9996 5714
rect 10336 5370 10364 5850
rect 10428 5778 10456 6190
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10414 5400 10470 5409
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10324 5364 10376 5370
rect 10414 5335 10416 5344
rect 10324 5306 10376 5312
rect 10468 5335 10470 5344
rect 10416 5306 10468 5312
rect 10612 5234 10640 6258
rect 11624 6254 11652 7142
rect 10692 6248 10744 6254
rect 11612 6248 11664 6254
rect 10692 6190 10744 6196
rect 11532 6208 11612 6236
rect 10704 5710 10732 6190
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9416 4078 9444 4422
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 8102 3836 8410 3845
rect 8102 3834 8108 3836
rect 8164 3834 8188 3836
rect 8244 3834 8268 3836
rect 8324 3834 8348 3836
rect 8404 3834 8410 3836
rect 8164 3782 8166 3834
rect 8346 3782 8348 3834
rect 8102 3780 8108 3782
rect 8164 3780 8188 3782
rect 8244 3780 8268 3782
rect 8324 3780 8348 3782
rect 8404 3780 8410 3782
rect 8102 3771 8410 3780
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 5460 3046 5580 3074
rect 5262 2952 5318 2961
rect 3976 2916 4028 2922
rect 5448 2916 5500 2922
rect 5262 2887 5318 2896
rect 3976 2858 4028 2864
rect 2792 2746 3096 2774
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 2700 2106 2728 2518
rect 2792 2514 2820 2746
rect 3988 2650 4016 2858
rect 5276 2854 5304 2887
rect 5368 2876 5448 2904
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 5368 2582 5396 2876
rect 5448 2858 5500 2864
rect 5552 2802 5580 3046
rect 5460 2774 5580 2802
rect 5356 2576 5408 2582
rect 5356 2518 5408 2524
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2688 2100 2740 2106
rect 2688 2042 2740 2048
rect 2792 1902 2820 2450
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3344 2106 3372 2314
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 4250 2204 4558 2213
rect 4250 2202 4256 2204
rect 4312 2202 4336 2204
rect 4392 2202 4416 2204
rect 4472 2202 4496 2204
rect 4552 2202 4558 2204
rect 4312 2150 4314 2202
rect 4494 2150 4496 2202
rect 4250 2148 4256 2150
rect 4312 2148 4336 2150
rect 4392 2148 4416 2150
rect 4472 2148 4496 2150
rect 4552 2148 4558 2150
rect 4250 2139 4558 2148
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 4632 1902 4660 2246
rect 4724 2038 4752 2246
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 5184 1902 5212 2246
rect 5460 1902 5488 2774
rect 6840 2038 6868 3538
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7116 2774 7144 2858
rect 7024 2746 7144 2774
rect 7024 2582 7052 2746
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 7024 2038 7052 2518
rect 7208 2106 7236 3130
rect 7944 3058 7972 3470
rect 8128 3194 8156 3538
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7944 2514 7972 2994
rect 9416 2990 9444 4014
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 8102 2748 8410 2757
rect 8102 2746 8108 2748
rect 8164 2746 8188 2748
rect 8244 2746 8268 2748
rect 8324 2746 8348 2748
rect 8404 2746 8410 2748
rect 8164 2694 8166 2746
rect 8346 2694 8348 2746
rect 8102 2692 8108 2694
rect 8164 2692 8188 2694
rect 8244 2692 8268 2694
rect 8324 2692 8348 2694
rect 8404 2692 8410 2694
rect 8102 2683 8410 2692
rect 9416 2514 9444 2926
rect 10428 2922 10456 4966
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10704 4146 10732 4694
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 11256 3126 11284 4966
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11348 4078 11376 4762
rect 11428 4480 11480 4486
rect 11532 4468 11560 6208
rect 11612 6190 11664 6196
rect 11610 5944 11666 5953
rect 11610 5879 11666 5888
rect 11624 5846 11652 5879
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11612 4548 11664 4554
rect 11716 4536 11744 9454
rect 11888 9444 11940 9450
rect 12072 9444 12124 9450
rect 11940 9404 12072 9432
rect 11888 9386 11940 9392
rect 12072 9386 12124 9392
rect 11955 8732 12263 8741
rect 11955 8730 11961 8732
rect 12017 8730 12041 8732
rect 12097 8730 12121 8732
rect 12177 8730 12201 8732
rect 12257 8730 12263 8732
rect 12017 8678 12019 8730
rect 12199 8678 12201 8730
rect 11955 8676 11961 8678
rect 12017 8676 12041 8678
rect 12097 8676 12121 8678
rect 12177 8676 12201 8678
rect 12257 8676 12263 8678
rect 11955 8667 12263 8676
rect 11888 8560 11940 8566
rect 11808 8520 11888 8548
rect 11808 5352 11836 8520
rect 11888 8502 11940 8508
rect 12360 8430 12388 9454
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 11955 7644 12263 7653
rect 11955 7642 11961 7644
rect 12017 7642 12041 7644
rect 12097 7642 12121 7644
rect 12177 7642 12201 7644
rect 12257 7642 12263 7644
rect 12017 7590 12019 7642
rect 12199 7590 12201 7642
rect 11955 7588 11961 7590
rect 12017 7588 12041 7590
rect 12097 7588 12121 7590
rect 12177 7588 12201 7590
rect 12257 7588 12263 7590
rect 11955 7579 12263 7588
rect 12452 7342 12480 9823
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12544 8430 12572 9658
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 9178 12756 9454
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12728 8673 12756 8774
rect 12714 8664 12770 8673
rect 12714 8599 12770 8608
rect 12532 8424 12584 8430
rect 12716 8424 12768 8430
rect 12532 8366 12584 8372
rect 12714 8392 12716 8401
rect 12768 8392 12770 8401
rect 12544 7954 12572 8366
rect 12714 8327 12770 8336
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12820 7834 12848 12192
rect 13188 12102 13216 12922
rect 13464 12646 13492 15846
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13648 13802 13676 14758
rect 13740 13802 13768 15098
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14200 14618 14228 14758
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13648 13161 13676 13398
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13634 13152 13690 13161
rect 13634 13087 13690 13096
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12912 11218 12940 11562
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 13188 10810 13216 12038
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 8634 12940 10406
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13280 9761 13308 9930
rect 13266 9752 13322 9761
rect 13266 9687 13322 9696
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13004 8634 13032 8978
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 8090 13032 8230
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12728 7806 12848 7834
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12452 6914 12480 7278
rect 12360 6886 12480 6914
rect 12532 6928 12584 6934
rect 12254 6760 12310 6769
rect 12254 6695 12256 6704
rect 12308 6695 12310 6704
rect 12256 6666 12308 6672
rect 11955 6556 12263 6565
rect 11955 6554 11961 6556
rect 12017 6554 12041 6556
rect 12097 6554 12121 6556
rect 12177 6554 12201 6556
rect 12257 6554 12263 6556
rect 12017 6502 12019 6554
rect 12199 6502 12201 6554
rect 11955 6500 11961 6502
rect 12017 6500 12041 6502
rect 12097 6500 12121 6502
rect 12177 6500 12201 6502
rect 12257 6500 12263 6502
rect 11955 6491 12263 6500
rect 12360 5914 12388 6886
rect 12532 6870 12584 6876
rect 12544 6225 12572 6870
rect 12636 6780 12664 7686
rect 12728 7206 12756 7806
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12820 7041 12848 7686
rect 12912 7546 12940 7686
rect 13004 7546 13032 7686
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12806 7032 12862 7041
rect 12806 6967 12862 6976
rect 13096 6798 13124 8978
rect 12716 6792 12768 6798
rect 12636 6752 12716 6780
rect 12716 6734 12768 6740
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 6458 12756 6598
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 13082 6352 13138 6361
rect 13082 6287 13138 6296
rect 12530 6216 12586 6225
rect 12530 6151 12586 6160
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12728 5914 12756 6122
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12268 5556 12296 5714
rect 12440 5568 12492 5574
rect 12268 5528 12388 5556
rect 11955 5468 12263 5477
rect 11955 5466 11961 5468
rect 12017 5466 12041 5468
rect 12097 5466 12121 5468
rect 12177 5466 12201 5468
rect 12257 5466 12263 5468
rect 12017 5414 12019 5466
rect 12199 5414 12201 5466
rect 11955 5412 11961 5414
rect 12017 5412 12041 5414
rect 12097 5412 12121 5414
rect 12177 5412 12201 5414
rect 12257 5412 12263 5414
rect 11955 5403 12263 5412
rect 12360 5370 12388 5528
rect 12440 5510 12492 5516
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12348 5364 12400 5370
rect 11808 5324 12112 5352
rect 12084 4826 12112 5324
rect 12348 5306 12400 5312
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12176 4758 12204 5034
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11664 4508 11744 4536
rect 11612 4490 11664 4496
rect 11480 4440 11560 4468
rect 11428 4422 11480 4428
rect 11532 4282 11560 4440
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11808 4010 11836 4626
rect 11980 4480 12032 4486
rect 11900 4440 11980 4468
rect 11900 4434 11928 4440
rect 11880 4406 11928 4434
rect 11980 4422 12032 4428
rect 11880 4298 11908 4406
rect 11955 4380 12263 4389
rect 11955 4378 11961 4380
rect 12017 4378 12041 4380
rect 12097 4378 12121 4380
rect 12177 4378 12201 4380
rect 12257 4378 12263 4380
rect 12017 4326 12019 4378
rect 12199 4326 12201 4378
rect 11955 4324 11961 4326
rect 12017 4324 12041 4326
rect 12097 4324 12121 4326
rect 12177 4324 12201 4326
rect 12257 4324 12263 4326
rect 11955 4315 12263 4324
rect 11880 4282 11928 4298
rect 11880 4276 11940 4282
rect 11880 4270 11888 4276
rect 11888 4218 11940 4224
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 11532 3194 11560 3946
rect 11978 3768 12034 3777
rect 11978 3703 12034 3712
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 10416 2916 10468 2922
rect 10416 2858 10468 2864
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 6828 2032 6880 2038
rect 6828 1974 6880 1980
rect 7012 2032 7064 2038
rect 7012 1974 7064 1980
rect 6840 1902 6868 1974
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 4620 1896 4672 1902
rect 4620 1838 4672 1844
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 5448 1896 5500 1902
rect 5448 1838 5500 1844
rect 6828 1896 6880 1902
rect 6828 1838 6880 1844
rect 7208 1562 7236 2042
rect 7300 2038 7328 2246
rect 8220 2106 8248 2450
rect 9692 2106 9720 2450
rect 7840 2100 7892 2106
rect 7840 2042 7892 2048
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 7288 2032 7340 2038
rect 7288 1974 7340 1980
rect 7300 1562 7328 1974
rect 7852 1562 7880 2042
rect 9876 1902 9904 2858
rect 8116 1896 8168 1902
rect 8116 1838 8168 1844
rect 9496 1896 9548 1902
rect 9496 1838 9548 1844
rect 9864 1896 9916 1902
rect 9864 1838 9916 1844
rect 8128 1748 8156 1838
rect 8036 1720 8156 1748
rect 9404 1760 9456 1766
rect 7196 1556 7248 1562
rect 7196 1498 7248 1504
rect 7288 1556 7340 1562
rect 7288 1498 7340 1504
rect 7840 1556 7892 1562
rect 7840 1498 7892 1504
rect 4250 1116 4558 1125
rect 4250 1114 4256 1116
rect 4312 1114 4336 1116
rect 4392 1114 4416 1116
rect 4472 1114 4496 1116
rect 4552 1114 4558 1116
rect 4312 1062 4314 1114
rect 4494 1062 4496 1114
rect 4250 1060 4256 1062
rect 4312 1060 4336 1062
rect 4392 1060 4416 1062
rect 4472 1060 4496 1062
rect 4552 1060 4558 1062
rect 4250 1051 4558 1060
rect 7852 814 7880 1498
rect 8036 1358 8064 1720
rect 9404 1702 9456 1708
rect 8102 1660 8410 1669
rect 8102 1658 8108 1660
rect 8164 1658 8188 1660
rect 8244 1658 8268 1660
rect 8324 1658 8348 1660
rect 8404 1658 8410 1660
rect 8164 1606 8166 1658
rect 8346 1606 8348 1658
rect 8102 1604 8108 1606
rect 8164 1604 8188 1606
rect 8244 1604 8268 1606
rect 8324 1604 8348 1606
rect 8404 1604 8410 1606
rect 8102 1595 8410 1604
rect 9416 1494 9444 1702
rect 9508 1562 9536 1838
rect 9680 1760 9732 1766
rect 9680 1702 9732 1708
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 8484 1488 8536 1494
rect 8484 1430 8536 1436
rect 9404 1488 9456 1494
rect 9404 1430 9456 1436
rect 8024 1352 8076 1358
rect 8024 1294 8076 1300
rect 8036 1018 8064 1294
rect 8496 1018 8524 1430
rect 9416 1018 9444 1430
rect 9692 1426 9720 1702
rect 9680 1420 9732 1426
rect 9680 1362 9732 1368
rect 9692 1018 9720 1362
rect 8024 1012 8076 1018
rect 8024 954 8076 960
rect 8484 1012 8536 1018
rect 8484 954 8536 960
rect 9404 1012 9456 1018
rect 9404 954 9456 960
rect 9680 1012 9732 1018
rect 9680 954 9732 960
rect 9876 882 9904 1838
rect 10600 1828 10652 1834
rect 10600 1770 10652 1776
rect 10612 1426 10640 1770
rect 11072 1494 11100 2858
rect 11624 2650 11652 3606
rect 11992 3398 12020 3703
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11955 3292 12263 3301
rect 11955 3290 11961 3292
rect 12017 3290 12041 3292
rect 12097 3290 12121 3292
rect 12177 3290 12201 3292
rect 12257 3290 12263 3292
rect 12017 3238 12019 3290
rect 12199 3238 12201 3290
rect 11955 3236 11961 3238
rect 12017 3236 12041 3238
rect 12097 3236 12121 3238
rect 12177 3236 12201 3238
rect 12257 3236 12263 3238
rect 11955 3227 12263 3236
rect 12452 2990 12480 5510
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12544 3641 12572 3946
rect 12530 3632 12586 3641
rect 12636 3602 12664 3946
rect 12530 3567 12586 3576
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12728 3194 12756 3538
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12820 3194 12848 3334
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12912 2922 12940 5510
rect 13096 5302 13124 6287
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11532 2106 11560 2450
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 11164 1494 11192 2042
rect 11612 1896 11664 1902
rect 11612 1838 11664 1844
rect 11624 1562 11652 1838
rect 11612 1556 11664 1562
rect 11612 1498 11664 1504
rect 11060 1488 11112 1494
rect 11060 1430 11112 1436
rect 11152 1488 11204 1494
rect 11152 1430 11204 1436
rect 10600 1420 10652 1426
rect 10600 1362 10652 1368
rect 9864 876 9916 882
rect 9864 818 9916 824
rect 10612 814 10640 1362
rect 11072 1018 11100 1430
rect 11612 1216 11664 1222
rect 11716 1170 11744 2450
rect 11955 2204 12263 2213
rect 11955 2202 11961 2204
rect 12017 2202 12041 2204
rect 12097 2202 12121 2204
rect 12177 2202 12201 2204
rect 12257 2202 12263 2204
rect 12017 2150 12019 2202
rect 12199 2150 12201 2202
rect 11955 2148 11961 2150
rect 12017 2148 12041 2150
rect 12097 2148 12121 2150
rect 12177 2148 12201 2150
rect 12257 2148 12263 2150
rect 11955 2139 12263 2148
rect 12348 1760 12400 1766
rect 12348 1702 12400 1708
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 11664 1164 11744 1170
rect 11612 1158 11744 1164
rect 11624 1142 11744 1158
rect 11060 1012 11112 1018
rect 11060 954 11112 960
rect 11716 950 11744 1142
rect 11955 1116 12263 1125
rect 11955 1114 11961 1116
rect 12017 1114 12041 1116
rect 12097 1114 12121 1116
rect 12177 1114 12201 1116
rect 12257 1114 12263 1116
rect 12017 1062 12019 1114
rect 12199 1062 12201 1114
rect 11955 1060 11961 1062
rect 12017 1060 12041 1062
rect 12097 1060 12121 1062
rect 12177 1060 12201 1062
rect 12257 1060 12263 1062
rect 11955 1051 12263 1060
rect 11704 944 11756 950
rect 11704 886 11756 892
rect 12360 814 12388 1702
rect 12636 1426 12664 1702
rect 12820 1562 12848 2858
rect 13004 2106 13032 5034
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13096 2650 13124 4558
rect 13188 3194 13216 9522
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13280 8634 13308 8978
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13372 8566 13400 12038
rect 13556 11608 13584 12718
rect 13740 12434 13768 13330
rect 13464 11580 13584 11608
rect 13648 12406 13768 12434
rect 13464 9518 13492 11580
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13556 9926 13584 11086
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13450 8936 13506 8945
rect 13450 8871 13452 8880
rect 13504 8871 13506 8880
rect 13544 8900 13596 8906
rect 13452 8842 13504 8848
rect 13544 8842 13596 8848
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13372 8022 13400 8366
rect 13450 8120 13506 8129
rect 13450 8055 13506 8064
rect 13464 8022 13492 8055
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13452 8016 13504 8022
rect 13452 7958 13504 7964
rect 13280 6934 13308 7958
rect 13464 7342 13492 7958
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13464 7002 13492 7278
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13280 6718 13492 6746
rect 13280 5574 13308 6718
rect 13464 6662 13492 6718
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13372 6458 13400 6598
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13372 5386 13400 6190
rect 13280 5358 13400 5386
rect 13280 4826 13308 5358
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13280 4457 13308 4762
rect 13464 4690 13492 5102
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13266 4448 13322 4457
rect 13266 4383 13322 4392
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13280 2922 13308 3538
rect 13372 3210 13400 4558
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 13464 3534 13492 3606
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13556 3398 13584 8842
rect 13648 6118 13676 12406
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13740 10130 13768 12310
rect 13832 12238 13860 14010
rect 14016 13870 14044 14486
rect 14476 14482 14504 14758
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14004 13728 14056 13734
rect 13910 13696 13966 13705
rect 14004 13670 14056 13676
rect 13910 13631 13966 13640
rect 13924 12866 13952 13631
rect 14016 12986 14044 13670
rect 14108 13376 14136 13874
rect 14200 13512 14228 14214
rect 14292 13938 14320 14214
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14200 13484 14412 13512
rect 14384 13394 14412 13484
rect 14280 13388 14332 13394
rect 14108 13348 14228 13376
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13924 12838 14044 12866
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13924 12617 13952 12718
rect 13910 12608 13966 12617
rect 13910 12543 13966 12552
rect 13910 12472 13966 12481
rect 13910 12407 13966 12416
rect 14016 12434 14044 12838
rect 14108 12764 14136 13194
rect 14200 12986 14228 13348
rect 14280 13330 14332 13336
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14292 12889 14320 13330
rect 14568 13308 14596 16390
rect 14456 13280 14596 13308
rect 14456 13274 14484 13280
rect 14384 13246 14484 13274
rect 14278 12880 14334 12889
rect 14278 12815 14334 12824
rect 14188 12776 14240 12782
rect 14108 12736 14188 12764
rect 14188 12718 14240 12724
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13818 11792 13874 11801
rect 13818 11727 13874 11736
rect 13832 11694 13860 11727
rect 13924 11694 13952 12407
rect 14016 12406 14136 12434
rect 14108 11762 14136 12406
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13924 10826 13952 11630
rect 13832 10798 13952 10826
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9722 13768 9862
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13832 9602 13860 10798
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13924 10198 13952 10678
rect 14016 10305 14044 11630
rect 14200 11529 14228 12718
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 14186 11520 14242 11529
rect 14186 11455 14242 11464
rect 14200 11218 14228 11455
rect 14292 11354 14320 11562
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14384 10538 14412 13246
rect 14660 13172 14688 17478
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14844 13938 14872 16186
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15488 15706 15516 15914
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 14936 14958 14964 15370
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 15016 14544 15068 14550
rect 15014 14512 15016 14521
rect 15068 14512 15070 14521
rect 15014 14447 15070 14456
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14568 13144 14688 13172
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14476 10810 14504 10950
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14568 10538 14596 13144
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 14660 11694 14688 12854
rect 14752 12714 14780 13874
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14844 13394 14872 13670
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14844 12730 14872 13126
rect 14936 12918 14964 13874
rect 15120 13802 15148 15302
rect 15396 15162 15424 15302
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15200 14476 15252 14482
rect 15304 14464 15332 15030
rect 15488 15026 15516 15302
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15580 14890 15608 15370
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15252 14436 15332 14464
rect 15200 14418 15252 14424
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15212 13802 15240 13942
rect 15304 13938 15332 14214
rect 15488 14074 15516 14282
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15200 13796 15252 13802
rect 15384 13796 15436 13802
rect 15200 13738 15252 13744
rect 15304 13756 15384 13784
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 14740 12708 14792 12714
rect 14844 12702 15056 12730
rect 14740 12650 14792 12656
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14752 11626 14780 12650
rect 15028 12434 15056 12702
rect 15028 12406 15148 12434
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14740 11620 14792 11626
rect 14740 11562 14792 11568
rect 14752 10810 14780 11562
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14738 10704 14794 10713
rect 14738 10639 14794 10648
rect 14752 10538 14780 10639
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 14556 10532 14608 10538
rect 14556 10474 14608 10480
rect 14740 10532 14792 10538
rect 14740 10474 14792 10480
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14186 10432 14242 10441
rect 14002 10296 14058 10305
rect 14002 10231 14058 10240
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13740 9574 13860 9602
rect 13740 7970 13768 9574
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13832 8090 13860 8366
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13740 7942 13860 7970
rect 13832 7750 13860 7942
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13726 6896 13782 6905
rect 13832 6866 13860 7686
rect 13924 7546 13952 9658
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 13726 6831 13782 6840
rect 13820 6860 13872 6866
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13634 5128 13690 5137
rect 13634 5063 13690 5072
rect 13648 4826 13676 5063
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13648 4282 13676 4626
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13740 3466 13768 6831
rect 13820 6802 13872 6808
rect 13924 6338 13952 6938
rect 14016 6866 14044 10231
rect 14108 9926 14136 10406
rect 14186 10367 14242 10376
rect 14200 10130 14228 10367
rect 14278 10160 14334 10169
rect 14188 10124 14240 10130
rect 14844 10146 14872 11834
rect 14936 10810 14964 12174
rect 15014 11792 15070 11801
rect 15014 11727 15070 11736
rect 15028 11558 15056 11727
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14924 10464 14976 10470
rect 14976 10424 15056 10452
rect 14924 10406 14976 10412
rect 14278 10095 14280 10104
rect 14188 10066 14240 10072
rect 14332 10095 14334 10104
rect 14384 10118 14872 10146
rect 14280 10066 14332 10072
rect 14278 10024 14334 10033
rect 14278 9959 14334 9968
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14292 9489 14320 9959
rect 14278 9480 14334 9489
rect 14278 9415 14334 9424
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14200 8566 14228 9114
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14096 7812 14148 7818
rect 14096 7754 14148 7760
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14002 6488 14058 6497
rect 14002 6423 14004 6432
rect 14056 6423 14058 6432
rect 14004 6394 14056 6400
rect 13924 6310 14044 6338
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13832 4826 13860 6190
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13832 3466 13860 3878
rect 13924 3738 13952 6190
rect 14016 4486 14044 6310
rect 14108 5846 14136 7754
rect 14200 6746 14228 8366
rect 14292 7993 14320 8774
rect 14278 7984 14334 7993
rect 14278 7919 14334 7928
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7342 14320 7822
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14292 6934 14320 7278
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 14200 6718 14320 6746
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 14108 5370 14136 5782
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14200 4826 14228 6598
rect 14292 5914 14320 6718
rect 14384 6458 14412 10118
rect 14740 10056 14792 10062
rect 14476 10016 14740 10044
rect 14476 6458 14504 10016
rect 14740 9998 14792 10004
rect 14556 9920 14608 9926
rect 14648 9920 14700 9926
rect 14556 9862 14608 9868
rect 14646 9888 14648 9897
rect 14740 9920 14792 9926
rect 14700 9888 14702 9897
rect 14568 9178 14596 9862
rect 14740 9862 14792 9868
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14646 9823 14702 9832
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14568 9042 14596 9114
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14554 8664 14610 8673
rect 14554 8599 14556 8608
rect 14608 8599 14610 8608
rect 14556 8570 14608 8576
rect 14568 8430 14596 8570
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 8129 14596 8230
rect 14554 8120 14610 8129
rect 14554 8055 14610 8064
rect 14568 7410 14596 8055
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14660 7002 14688 9658
rect 14752 9500 14780 9862
rect 14844 9722 14872 9862
rect 14922 9752 14978 9761
rect 14832 9716 14884 9722
rect 14922 9687 14924 9696
rect 14832 9658 14884 9664
rect 14976 9687 14978 9696
rect 14924 9658 14976 9664
rect 14922 9616 14978 9625
rect 14922 9551 14978 9560
rect 14832 9512 14884 9518
rect 14752 9472 14832 9500
rect 14832 9454 14884 9460
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14752 8294 14780 9318
rect 14844 8820 14872 9318
rect 14936 9178 14964 9551
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14924 8832 14976 8838
rect 14844 8792 14924 8820
rect 14924 8774 14976 8780
rect 15028 8634 15056 10424
rect 15120 9722 15148 12406
rect 15212 12306 15240 13126
rect 15304 12306 15332 13756
rect 15384 13738 15436 13744
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15396 12442 15424 13398
rect 15488 13190 15516 14010
rect 15568 13796 15620 13802
rect 15672 13784 15700 17478
rect 15807 16892 16115 16901
rect 15807 16890 15813 16892
rect 15869 16890 15893 16892
rect 15949 16890 15973 16892
rect 16029 16890 16053 16892
rect 16109 16890 16115 16892
rect 15869 16838 15871 16890
rect 16051 16838 16053 16890
rect 15807 16836 15813 16838
rect 15869 16836 15893 16838
rect 15949 16836 15973 16838
rect 16029 16836 16053 16838
rect 16109 16836 16115 16838
rect 15807 16827 16115 16836
rect 16026 16008 16082 16017
rect 16026 15943 16082 15952
rect 16040 15910 16068 15943
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 15807 15804 16115 15813
rect 15807 15802 15813 15804
rect 15869 15802 15893 15804
rect 15949 15802 15973 15804
rect 16029 15802 16053 15804
rect 16109 15802 16115 15804
rect 15869 15750 15871 15802
rect 16051 15750 16053 15802
rect 15807 15748 15813 15750
rect 15869 15748 15893 15750
rect 15949 15748 15973 15750
rect 16029 15748 16053 15750
rect 16109 15748 16115 15750
rect 15807 15739 16115 15748
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15856 14958 15884 15438
rect 16224 15026 16252 17682
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15807 14716 16115 14725
rect 15807 14714 15813 14716
rect 15869 14714 15893 14716
rect 15949 14714 15973 14716
rect 16029 14714 16053 14716
rect 16109 14714 16115 14716
rect 15869 14662 15871 14714
rect 16051 14662 16053 14714
rect 15807 14660 15813 14662
rect 15869 14660 15893 14662
rect 15949 14660 15973 14662
rect 16029 14660 16053 14662
rect 16109 14660 16115 14662
rect 15807 14651 16115 14660
rect 16224 14482 16252 14962
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16120 13864 16172 13870
rect 16172 13824 16252 13852
rect 16120 13806 16172 13812
rect 15936 13796 15988 13802
rect 15672 13756 15936 13784
rect 15568 13738 15620 13744
rect 15936 13738 15988 13744
rect 15580 13297 15608 13738
rect 15807 13628 16115 13637
rect 15807 13626 15813 13628
rect 15869 13626 15893 13628
rect 15949 13626 15973 13628
rect 16029 13626 16053 13628
rect 16109 13626 16115 13628
rect 15869 13574 15871 13626
rect 16051 13574 16053 13626
rect 15807 13572 15813 13574
rect 15869 13572 15893 13574
rect 15949 13572 15973 13574
rect 16029 13572 16053 13574
rect 16109 13572 16115 13574
rect 15807 13563 16115 13572
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15566 13288 15622 13297
rect 15566 13223 15622 13232
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15658 13152 15714 13161
rect 15658 13087 15714 13096
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15488 12481 15516 12718
rect 15474 12472 15530 12481
rect 15384 12436 15436 12442
rect 15474 12407 15476 12416
rect 15384 12378 15436 12384
rect 15528 12407 15530 12416
rect 15672 12434 15700 13087
rect 15764 12782 15792 13330
rect 16224 12918 16252 13824
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15807 12540 16115 12549
rect 15807 12538 15813 12540
rect 15869 12538 15893 12540
rect 15949 12538 15973 12540
rect 16029 12538 16053 12540
rect 16109 12538 16115 12540
rect 15869 12486 15871 12538
rect 16051 12486 16053 12538
rect 15807 12484 15813 12486
rect 15869 12484 15893 12486
rect 15949 12484 15973 12486
rect 16029 12484 16053 12486
rect 16109 12484 16115 12486
rect 15807 12475 16115 12484
rect 15672 12406 15792 12434
rect 15476 12378 15528 12384
rect 15764 12306 15792 12406
rect 16026 12336 16082 12345
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15752 12300 15804 12306
rect 16026 12271 16082 12280
rect 15752 12242 15804 12248
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15212 12073 15240 12106
rect 15198 12064 15254 12073
rect 15198 11999 15254 12008
rect 15580 11626 15608 12242
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15108 9580 15160 9586
rect 15212 9568 15240 10406
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15304 9761 15332 9998
rect 15396 9926 15424 10406
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15290 9752 15346 9761
rect 15290 9687 15346 9696
rect 15212 9540 15332 9568
rect 15108 9522 15160 9528
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14752 8266 14872 8294
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14844 7834 14872 8266
rect 15120 8090 15148 9522
rect 15198 9480 15254 9489
rect 15198 9415 15200 9424
rect 15252 9415 15254 9424
rect 15200 9386 15252 9392
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15212 8090 15240 8842
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15304 8022 15332 9540
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15396 9178 15424 9454
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15488 8974 15516 10474
rect 15580 10130 15608 11562
rect 15672 11393 15700 12242
rect 15934 12200 15990 12209
rect 16040 12170 16068 12271
rect 15934 12135 15936 12144
rect 15988 12135 15990 12144
rect 16028 12164 16080 12170
rect 15936 12106 15988 12112
rect 16028 12106 16080 12112
rect 16026 11792 16082 11801
rect 16082 11750 16252 11778
rect 16026 11727 16082 11736
rect 16224 11529 16252 11750
rect 16210 11520 16266 11529
rect 15807 11452 16115 11461
rect 16210 11455 16266 11464
rect 15807 11450 15813 11452
rect 15869 11450 15893 11452
rect 15949 11450 15973 11452
rect 16029 11450 16053 11452
rect 16109 11450 16115 11452
rect 15869 11398 15871 11450
rect 16051 11398 16053 11450
rect 15807 11396 15813 11398
rect 15869 11396 15893 11398
rect 15949 11396 15973 11398
rect 16029 11396 16053 11398
rect 16109 11396 16115 11398
rect 15658 11384 15714 11393
rect 15807 11387 16115 11396
rect 15658 11319 15714 11328
rect 16028 11348 16080 11354
rect 16316 11336 16344 18022
rect 16488 17808 16540 17814
rect 16592 17796 16620 18022
rect 16540 17768 16620 17796
rect 16488 17750 16540 17756
rect 16960 17746 16988 18022
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16856 17264 16908 17270
rect 16856 17206 16908 17212
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16500 13784 16528 15846
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16776 14958 16804 15302
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16764 13864 16816 13870
rect 16762 13832 16764 13841
rect 16816 13832 16818 13841
rect 16672 13796 16724 13802
rect 16500 13756 16672 13784
rect 16762 13767 16818 13776
rect 16672 13738 16724 13744
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16408 13190 16436 13670
rect 16868 13530 16896 17206
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16486 13152 16542 13161
rect 16486 13087 16542 13096
rect 16500 12986 16528 13087
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16486 12472 16542 12481
rect 16486 12407 16542 12416
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16028 11290 16080 11296
rect 16132 11308 16344 11336
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15750 10840 15806 10849
rect 15660 10804 15712 10810
rect 15750 10775 15806 10784
rect 15660 10746 15712 10752
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15672 9674 15700 10746
rect 15764 10577 15792 10775
rect 15856 10606 15884 11018
rect 16040 11014 16068 11290
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15844 10600 15896 10606
rect 15750 10568 15806 10577
rect 15936 10600 15988 10606
rect 15844 10542 15896 10548
rect 15934 10568 15936 10577
rect 15988 10568 15990 10577
rect 15750 10503 15806 10512
rect 15934 10503 15990 10512
rect 16040 10452 16068 10746
rect 16132 10674 16160 11308
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16316 10588 16344 10950
rect 16408 10810 16436 12242
rect 16500 12238 16528 12407
rect 16592 12306 16620 13466
rect 16776 13433 16804 13466
rect 16762 13424 16818 13433
rect 16960 13410 16988 13670
rect 16868 13394 16988 13410
rect 16762 13359 16818 13368
rect 16856 13388 16988 13394
rect 16908 13382 16988 13388
rect 16856 13330 16908 13336
rect 17052 13308 17080 18566
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17144 13394 17172 13670
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 16960 13280 17080 13308
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16868 13025 16896 13126
rect 16854 13016 16910 13025
rect 16672 12980 16724 12986
rect 16854 12951 16910 12960
rect 16672 12922 16724 12928
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16396 10600 16448 10606
rect 16316 10560 16396 10588
rect 16396 10542 16448 10548
rect 16304 10464 16356 10470
rect 16040 10441 16252 10452
rect 16040 10432 16266 10441
rect 16040 10424 16210 10432
rect 16304 10406 16356 10412
rect 15807 10364 16115 10373
rect 16210 10367 16266 10376
rect 15807 10362 15813 10364
rect 15869 10362 15893 10364
rect 15949 10362 15973 10364
rect 16029 10362 16053 10364
rect 16109 10362 16115 10364
rect 15869 10310 15871 10362
rect 16051 10310 16053 10362
rect 15807 10308 15813 10310
rect 15869 10308 15893 10310
rect 15949 10308 15973 10310
rect 16029 10308 16053 10310
rect 16109 10308 16115 10310
rect 15807 10299 16115 10308
rect 16224 10248 16252 10367
rect 16316 10305 16344 10406
rect 16132 10220 16252 10248
rect 16302 10296 16358 10305
rect 16302 10231 16358 10240
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15764 9897 15792 10066
rect 15750 9888 15806 9897
rect 15750 9823 15806 9832
rect 15580 9646 15700 9674
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15384 8424 15436 8430
rect 15476 8424 15528 8430
rect 15384 8366 15436 8372
rect 15474 8392 15476 8401
rect 15528 8392 15530 8401
rect 15292 8016 15344 8022
rect 15292 7958 15344 7964
rect 14922 7848 14978 7857
rect 14752 7546 14780 7822
rect 14844 7806 14922 7834
rect 14922 7783 14978 7792
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14752 6866 14780 7142
rect 15106 7032 15162 7041
rect 15028 6990 15106 7018
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14462 6216 14518 6225
rect 14372 6180 14424 6186
rect 14462 6151 14518 6160
rect 14372 6122 14424 6128
rect 14384 5953 14412 6122
rect 14370 5944 14426 5953
rect 14280 5908 14332 5914
rect 14370 5879 14426 5888
rect 14280 5850 14332 5856
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14292 4690 14320 5850
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14016 4282 14044 4422
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14292 3777 14320 3946
rect 14278 3768 14334 3777
rect 13912 3732 13964 3738
rect 14278 3703 14334 3712
rect 13912 3674 13964 3680
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 3210 13676 3334
rect 13372 3194 13676 3210
rect 13360 3188 13676 3194
rect 13412 3182 13676 3188
rect 13360 3130 13412 3136
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 13556 2774 13584 2926
rect 13556 2746 13676 2774
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 13648 2582 13676 2746
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 12992 2100 13044 2106
rect 12992 2042 13044 2048
rect 13188 1562 13216 2450
rect 12808 1556 12860 1562
rect 12808 1498 12860 1504
rect 13176 1556 13228 1562
rect 13176 1498 13228 1504
rect 12624 1420 12676 1426
rect 12624 1362 12676 1368
rect 13176 1420 13228 1426
rect 13176 1362 13228 1368
rect 12636 1018 12664 1362
rect 12624 1012 12676 1018
rect 12624 954 12676 960
rect 13188 814 13216 1362
rect 13740 1358 13768 2450
rect 14200 2310 14228 3606
rect 14384 3210 14412 4150
rect 14476 3534 14504 6151
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14568 3466 14596 6666
rect 14844 6458 14872 6734
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 14936 5778 14964 6190
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14936 5080 14964 5714
rect 15028 5522 15056 6990
rect 15106 6967 15162 6976
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15120 5914 15148 6598
rect 15212 6254 15240 7414
rect 15304 7002 15332 7958
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15304 6458 15332 6802
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15028 5494 15148 5522
rect 15016 5092 15068 5098
rect 14936 5052 15016 5080
rect 15016 5034 15068 5040
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14752 4758 14780 4966
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14660 4185 14688 4558
rect 14646 4176 14702 4185
rect 14646 4111 14702 4120
rect 14660 4010 14688 4111
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 14752 3720 14780 4694
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 14844 4282 14872 4558
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14844 4078 14872 4218
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14832 3732 14884 3738
rect 14752 3692 14832 3720
rect 14832 3674 14884 3680
rect 14648 3664 14700 3670
rect 14648 3606 14700 3612
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14384 3194 14504 3210
rect 14384 3188 14516 3194
rect 14384 3182 14464 3188
rect 14464 3130 14516 3136
rect 14372 2916 14424 2922
rect 14372 2858 14424 2864
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14384 1850 14412 2858
rect 14660 2650 14688 3606
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14936 3194 14964 3538
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 14384 1822 14780 1850
rect 13728 1352 13780 1358
rect 13728 1294 13780 1300
rect 13740 814 13768 1294
rect 14384 1290 14412 1822
rect 14464 1760 14516 1766
rect 14464 1702 14516 1708
rect 14556 1760 14608 1766
rect 14556 1702 14608 1708
rect 14476 1494 14504 1702
rect 14568 1562 14596 1702
rect 14752 1562 14780 1822
rect 14556 1556 14608 1562
rect 14556 1498 14608 1504
rect 14740 1556 14792 1562
rect 14740 1498 14792 1504
rect 14464 1488 14516 1494
rect 14464 1430 14516 1436
rect 14372 1284 14424 1290
rect 14372 1226 14424 1232
rect 14188 1216 14240 1222
rect 14188 1158 14240 1164
rect 14200 1018 14228 1158
rect 14476 1018 14504 1430
rect 14648 1216 14700 1222
rect 14648 1158 14700 1164
rect 14740 1216 14792 1222
rect 14740 1158 14792 1164
rect 14188 1012 14240 1018
rect 14188 954 14240 960
rect 14464 1012 14516 1018
rect 14464 954 14516 960
rect 14660 814 14688 1158
rect 14752 950 14780 1158
rect 15028 1018 15056 5034
rect 15120 3738 15148 5494
rect 15396 5370 15424 8366
rect 15474 8327 15530 8336
rect 15580 7954 15608 9646
rect 16132 9625 16160 10220
rect 16118 9616 16174 9625
rect 16118 9551 16174 9560
rect 16408 9518 16436 10542
rect 15660 9512 15712 9518
rect 16396 9512 16448 9518
rect 15660 9454 15712 9460
rect 15750 9480 15806 9489
rect 15672 8974 15700 9454
rect 16396 9454 16448 9460
rect 15750 9415 15752 9424
rect 15804 9415 15806 9424
rect 16120 9444 16172 9450
rect 15752 9386 15804 9392
rect 16500 9432 16528 11766
rect 16592 11762 16620 12038
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16578 11520 16634 11529
rect 16578 11455 16634 11464
rect 16592 11200 16620 11455
rect 16684 11354 16712 12922
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12306 16896 12582
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16776 11898 16804 12242
rect 16960 12220 16988 13280
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17052 12374 17080 12718
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 17040 12232 17092 12238
rect 16960 12192 17040 12220
rect 17040 12174 17092 12180
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16868 11801 16896 12038
rect 16960 11830 16988 12038
rect 16948 11824 17000 11830
rect 16854 11792 16910 11801
rect 16948 11766 17000 11772
rect 17236 11762 17264 13126
rect 16854 11727 16910 11736
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16762 11520 16818 11529
rect 16762 11455 16818 11464
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16672 11212 16724 11218
rect 16592 11172 16672 11200
rect 16672 11154 16724 11160
rect 16776 10962 16804 11455
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16868 11121 16896 11154
rect 16854 11112 16910 11121
rect 16854 11047 16910 11056
rect 16776 10934 16896 10962
rect 16578 10840 16634 10849
rect 16762 10840 16818 10849
rect 16684 10810 16762 10826
rect 16578 10775 16634 10784
rect 16672 10804 16762 10810
rect 16592 10520 16620 10775
rect 16724 10798 16762 10804
rect 16762 10775 16818 10784
rect 16672 10746 16724 10752
rect 16868 10674 16896 10934
rect 16856 10668 16908 10674
rect 16776 10628 16856 10656
rect 16672 10532 16724 10538
rect 16592 10492 16672 10520
rect 16672 10474 16724 10480
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 9722 16620 9862
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16670 9616 16726 9625
rect 16670 9551 16726 9560
rect 16172 9404 16252 9432
rect 16500 9404 16620 9432
rect 16120 9386 16172 9392
rect 15807 9276 16115 9285
rect 15807 9274 15813 9276
rect 15869 9274 15893 9276
rect 15949 9274 15973 9276
rect 16029 9274 16053 9276
rect 16109 9274 16115 9276
rect 15869 9222 15871 9274
rect 16051 9222 16053 9274
rect 15807 9220 15813 9222
rect 15869 9220 15893 9222
rect 15949 9220 15973 9222
rect 16029 9220 16053 9222
rect 16109 9220 16115 9222
rect 15807 9211 16115 9220
rect 16120 9172 16172 9178
rect 16040 9132 16120 9160
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15856 8430 15884 8570
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 16040 8294 16068 9132
rect 16120 9114 16172 9120
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16132 8566 16160 8978
rect 16120 8560 16172 8566
rect 16120 8502 16172 8508
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15580 7546 15608 7890
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15672 6934 15700 8230
rect 15807 8188 16115 8197
rect 15807 8186 15813 8188
rect 15869 8186 15893 8188
rect 15949 8186 15973 8188
rect 16029 8186 16053 8188
rect 16109 8186 16115 8188
rect 15869 8134 15871 8186
rect 16051 8134 16053 8186
rect 15807 8132 15813 8134
rect 15869 8132 15893 8134
rect 15949 8132 15973 8134
rect 16029 8132 16053 8134
rect 16109 8132 16115 8134
rect 15807 8123 16115 8132
rect 16224 7546 16252 9404
rect 16394 9208 16450 9217
rect 16592 9194 16620 9404
rect 16394 9143 16450 9152
rect 16500 9166 16620 9194
rect 16684 9178 16712 9551
rect 16672 9172 16724 9178
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16316 7478 16344 8842
rect 16408 8634 16436 9143
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16408 8090 16436 8298
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16408 7478 16436 7890
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16500 7426 16528 9166
rect 16672 9114 16724 9120
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16592 8673 16620 8842
rect 16670 8800 16726 8809
rect 16670 8735 16726 8744
rect 16578 8664 16634 8673
rect 16578 8599 16634 8608
rect 16684 8548 16712 8735
rect 16776 8634 16804 10628
rect 16856 10610 16908 10616
rect 16960 10248 16988 11630
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17038 11248 17094 11257
rect 17038 11183 17040 11192
rect 17092 11183 17094 11192
rect 17040 11154 17092 11160
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 17052 10810 17080 11018
rect 17236 10985 17264 11290
rect 17222 10976 17278 10985
rect 17222 10911 17278 10920
rect 17328 10810 17356 13670
rect 17420 12850 17448 16934
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17512 12918 17540 14010
rect 17604 13734 17632 18686
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17788 16697 17816 17478
rect 17880 17202 17908 18702
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17774 16688 17830 16697
rect 17880 16658 17908 17138
rect 17774 16623 17830 16632
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17880 16114 17908 16594
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17682 15056 17738 15065
rect 17682 14991 17738 15000
rect 17696 14958 17724 14991
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17880 14657 17908 14894
rect 17866 14648 17922 14657
rect 17866 14583 17922 14592
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17788 13462 17816 13806
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17774 13152 17830 13161
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 11626 17448 12582
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17406 11384 17462 11393
rect 17512 11354 17540 12854
rect 17406 11319 17462 11328
rect 17500 11348 17552 11354
rect 17420 11218 17448 11319
rect 17500 11290 17552 11296
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17500 11144 17552 11150
rect 17604 11132 17632 13126
rect 17774 13087 17830 13096
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17696 12442 17724 12922
rect 17788 12918 17816 13087
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 17880 12782 17908 14350
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17972 12866 18000 14214
rect 18064 13802 18092 19600
rect 18708 19530 18736 19600
rect 18800 19530 18828 19638
rect 18708 19502 18828 19530
rect 18696 18148 18748 18154
rect 18696 18090 18748 18096
rect 18708 17814 18736 18090
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18696 17808 18748 17814
rect 18696 17750 18748 17756
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18156 16046 18184 16390
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18340 15570 18368 15846
rect 18524 15638 18552 15846
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18800 15162 18828 18022
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18696 14952 18748 14958
rect 18694 14920 18696 14929
rect 18748 14920 18750 14929
rect 18694 14855 18750 14864
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 18248 14618 18276 14758
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18878 14512 18934 14521
rect 18878 14447 18934 14456
rect 18892 14278 18920 14447
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 18328 13456 18380 13462
rect 18328 13398 18380 13404
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18064 13190 18092 13330
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 17972 12838 18092 12866
rect 17776 12776 17828 12782
rect 17774 12744 17776 12753
rect 17868 12776 17920 12782
rect 17828 12744 17830 12753
rect 17868 12718 17920 12724
rect 17774 12679 17830 12688
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17696 11529 17724 12242
rect 17682 11520 17738 11529
rect 17682 11455 17738 11464
rect 17788 11354 17816 12310
rect 17880 12170 17908 12718
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17880 11354 17908 11494
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17552 11104 17632 11132
rect 17500 11086 17552 11092
rect 17406 10976 17462 10985
rect 17406 10911 17462 10920
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 16868 10220 16988 10248
rect 16868 9722 16896 10220
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16960 9518 16988 10066
rect 17052 9722 17080 10406
rect 17144 9722 17172 10678
rect 17420 10674 17448 10911
rect 17696 10810 17724 11290
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17236 10169 17264 10406
rect 17222 10160 17278 10169
rect 17222 10095 17278 10104
rect 17328 9874 17356 10406
rect 17788 10169 17816 10406
rect 17774 10160 17830 10169
rect 17236 9846 17356 9874
rect 17696 10118 17774 10146
rect 17236 9722 17264 9846
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 17604 9625 17632 9658
rect 17590 9616 17646 9625
rect 17590 9551 17646 9560
rect 17696 9568 17724 10118
rect 17774 10095 17830 10104
rect 17880 9602 17908 11154
rect 17972 10130 18000 11562
rect 18064 11370 18092 12838
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18156 12442 18184 12718
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18248 12374 18276 13126
rect 18236 12368 18288 12374
rect 18142 12336 18198 12345
rect 18236 12310 18288 12316
rect 18142 12271 18198 12280
rect 18156 12238 18184 12271
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18248 11694 18276 12038
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18064 11342 18184 11370
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 18064 9674 18092 11222
rect 18156 10538 18184 11342
rect 18236 11212 18288 11218
rect 18236 11154 18288 11160
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 18142 10296 18198 10305
rect 18142 10231 18198 10240
rect 18156 9908 18184 10231
rect 18248 10062 18276 11154
rect 18340 11014 18368 13398
rect 18524 12442 18552 13942
rect 18696 13796 18748 13802
rect 18696 13738 18748 13744
rect 18708 13705 18736 13738
rect 18892 13734 18920 14214
rect 18788 13728 18840 13734
rect 18694 13696 18750 13705
rect 18788 13670 18840 13676
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18694 13631 18750 13640
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18616 12850 18644 13330
rect 18800 12866 18828 13670
rect 18892 13462 18920 13670
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18708 12838 18828 12866
rect 18602 12472 18658 12481
rect 18512 12436 18564 12442
rect 18602 12407 18658 12416
rect 18512 12378 18564 12384
rect 18616 12170 18644 12407
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18418 11928 18474 11937
rect 18418 11863 18474 11872
rect 18432 11694 18460 11863
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18340 10713 18368 10950
rect 18326 10704 18382 10713
rect 18326 10639 18382 10648
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18156 9880 18276 9908
rect 18064 9646 18184 9674
rect 18248 9654 18276 9880
rect 17880 9574 17954 9602
rect 17696 9540 17816 9568
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 17132 9512 17184 9518
rect 17788 9512 17816 9540
rect 17776 9506 17828 9512
rect 17184 9472 17264 9500
rect 17132 9454 17184 9460
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16592 8520 16712 8548
rect 16592 7857 16620 8520
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16684 8090 16712 8366
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 8090 16804 8230
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16578 7848 16634 7857
rect 16578 7783 16634 7792
rect 16500 7398 16620 7426
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 15807 7100 16115 7109
rect 15807 7098 15813 7100
rect 15869 7098 15893 7100
rect 15949 7098 15973 7100
rect 16029 7098 16053 7100
rect 16109 7098 16115 7100
rect 15869 7046 15871 7098
rect 16051 7046 16053 7098
rect 15807 7044 15813 7046
rect 15869 7044 15893 7046
rect 15949 7044 15973 7046
rect 16029 7044 16053 7046
rect 16109 7044 16115 7046
rect 15807 7035 16115 7044
rect 16500 7002 16528 7278
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 15948 6390 15976 6802
rect 16132 6390 16160 6802
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 15936 6384 15988 6390
rect 15936 6326 15988 6332
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15580 5778 15608 6190
rect 15807 6012 16115 6021
rect 15807 6010 15813 6012
rect 15869 6010 15893 6012
rect 15949 6010 15973 6012
rect 16029 6010 16053 6012
rect 16109 6010 16115 6012
rect 15869 5958 15871 6010
rect 16051 5958 16053 6010
rect 15807 5956 15813 5958
rect 15869 5956 15893 5958
rect 15949 5956 15973 5958
rect 16029 5956 16053 5958
rect 16109 5956 16115 5958
rect 15807 5947 16115 5956
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15580 5302 15608 5714
rect 16316 5534 16344 6598
rect 16592 6474 16620 7398
rect 16684 7342 16712 8026
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16776 6798 16804 6938
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16592 6446 16712 6474
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16224 5506 16344 5534
rect 15934 5400 15990 5409
rect 15934 5335 15936 5344
rect 15988 5335 15990 5344
rect 15936 5306 15988 5312
rect 15568 5296 15620 5302
rect 15290 5264 15346 5273
rect 15568 5238 15620 5244
rect 15290 5199 15346 5208
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15212 4282 15240 4558
rect 15304 4282 15332 5199
rect 16224 5166 16252 5506
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 15384 5160 15436 5166
rect 15660 5160 15712 5166
rect 15436 5120 15608 5148
rect 15384 5102 15436 5108
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15212 3398 15240 4218
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 15396 2394 15424 4694
rect 15488 4486 15516 4966
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15580 4321 15608 5120
rect 15660 5102 15712 5108
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 15672 4758 15700 5102
rect 15807 4924 16115 4933
rect 15807 4922 15813 4924
rect 15869 4922 15893 4924
rect 15949 4922 15973 4924
rect 16029 4922 16053 4924
rect 16109 4922 16115 4924
rect 15869 4870 15871 4922
rect 16051 4870 16053 4922
rect 15807 4868 15813 4870
rect 15869 4868 15893 4870
rect 15949 4868 15973 4870
rect 16029 4868 16053 4870
rect 16109 4868 16115 4870
rect 15807 4859 16115 4868
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 15566 4312 15622 4321
rect 15672 4282 15700 4694
rect 15844 4480 15896 4486
rect 15842 4448 15844 4457
rect 15896 4448 15898 4457
rect 15842 4383 15898 4392
rect 15566 4247 15622 4256
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15566 4176 15622 4185
rect 15566 4111 15622 4120
rect 15580 4078 15608 4111
rect 15856 4078 15884 4383
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15807 3836 16115 3845
rect 15807 3834 15813 3836
rect 15869 3834 15893 3836
rect 15949 3834 15973 3836
rect 16029 3834 16053 3836
rect 16109 3834 16115 3836
rect 15869 3782 15871 3834
rect 16051 3782 16053 3834
rect 15807 3780 15813 3782
rect 15869 3780 15893 3782
rect 15949 3780 15973 3782
rect 16029 3780 16053 3782
rect 16109 3780 16115 3782
rect 15807 3771 16115 3780
rect 16224 3670 16252 5102
rect 16316 4826 16344 5306
rect 16500 5302 16528 5714
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15488 2582 15516 2926
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 15807 2748 16115 2757
rect 15807 2746 15813 2748
rect 15869 2746 15893 2748
rect 15949 2746 15973 2748
rect 16029 2746 16053 2748
rect 16109 2746 16115 2748
rect 15869 2694 15871 2746
rect 16051 2694 16053 2746
rect 15807 2692 15813 2694
rect 15869 2692 15893 2694
rect 15949 2692 15973 2694
rect 16029 2692 16053 2694
rect 16109 2692 16115 2694
rect 15807 2683 16115 2692
rect 15476 2576 15528 2582
rect 16224 2530 16252 2858
rect 16316 2650 16344 3606
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 15476 2518 15528 2524
rect 16132 2502 16252 2530
rect 15396 2366 15608 2394
rect 15580 2310 15608 2366
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 16132 2106 16160 2502
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16120 2100 16172 2106
rect 16120 2042 16172 2048
rect 15200 1896 15252 1902
rect 15200 1838 15252 1844
rect 15476 1896 15528 1902
rect 15476 1838 15528 1844
rect 15660 1896 15712 1902
rect 15660 1838 15712 1844
rect 15212 1494 15240 1838
rect 15488 1562 15516 1838
rect 15672 1562 15700 1838
rect 15807 1660 16115 1669
rect 15807 1658 15813 1660
rect 15869 1658 15893 1660
rect 15949 1658 15973 1660
rect 16029 1658 16053 1660
rect 16109 1658 16115 1660
rect 15869 1606 15871 1658
rect 16051 1606 16053 1658
rect 15807 1604 15813 1606
rect 15869 1604 15893 1606
rect 15949 1604 15973 1606
rect 16029 1604 16053 1606
rect 16109 1604 16115 1606
rect 15807 1595 16115 1604
rect 15476 1556 15528 1562
rect 15476 1498 15528 1504
rect 15660 1556 15712 1562
rect 15660 1498 15712 1504
rect 15200 1488 15252 1494
rect 15200 1430 15252 1436
rect 15016 1012 15068 1018
rect 15016 954 15068 960
rect 14740 944 14792 950
rect 14740 886 14792 892
rect 16224 814 16252 2382
rect 16304 1896 16356 1902
rect 16304 1838 16356 1844
rect 16316 1562 16344 1838
rect 16408 1562 16436 5034
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16500 3738 16528 4422
rect 16592 4282 16620 4966
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16578 4040 16634 4049
rect 16578 3975 16634 3984
rect 16592 3942 16620 3975
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16684 3738 16712 6446
rect 16776 4758 16804 6598
rect 16868 6390 16896 9318
rect 17038 9072 17094 9081
rect 16948 9036 17000 9042
rect 17038 9007 17094 9016
rect 16948 8978 17000 8984
rect 16960 8430 16988 8978
rect 17052 8974 17080 9007
rect 17040 8968 17092 8974
rect 17092 8928 17172 8956
rect 17040 8910 17092 8916
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 17052 8294 17080 8774
rect 17144 8634 17172 8928
rect 17236 8820 17264 9472
rect 17776 9448 17828 9454
rect 17316 9376 17368 9382
rect 17926 9364 17954 9574
rect 17368 9336 17540 9364
rect 17316 9318 17368 9324
rect 17408 8832 17460 8838
rect 17236 8792 17408 8820
rect 17408 8774 17460 8780
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17316 8424 17368 8430
rect 17314 8392 17316 8401
rect 17408 8424 17460 8430
rect 17368 8392 17370 8401
rect 17408 8366 17460 8372
rect 17314 8327 17370 8336
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 16946 8120 17002 8129
rect 16946 8055 17002 8064
rect 17040 8084 17092 8090
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16868 5778 16896 6122
rect 16960 5778 16988 8055
rect 17040 8026 17092 8032
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16868 5098 16896 5714
rect 17052 5534 17080 8026
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 17236 7342 17264 7754
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17236 7002 17264 7278
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17328 6934 17356 7278
rect 17132 6928 17184 6934
rect 17132 6870 17184 6876
rect 17316 6928 17368 6934
rect 17316 6870 17368 6876
rect 17144 5794 17172 6870
rect 17144 5778 17356 5794
rect 17144 5772 17368 5778
rect 17144 5766 17316 5772
rect 17316 5714 17368 5720
rect 17052 5506 17356 5534
rect 16856 5092 16908 5098
rect 16856 5034 16908 5040
rect 16948 5024 17000 5030
rect 16868 4972 16948 4978
rect 16868 4966 17000 4972
rect 16868 4950 16988 4966
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16764 4276 16816 4282
rect 16764 4218 16816 4224
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16776 3398 16804 4218
rect 16868 4010 16896 4950
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16960 4321 16988 4422
rect 16946 4312 17002 4321
rect 17002 4270 17080 4298
rect 16946 4247 17002 4256
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 16960 3194 16988 3946
rect 17052 3942 17080 4270
rect 17328 4010 17356 5506
rect 17420 4282 17448 8366
rect 17512 8242 17540 9336
rect 17880 9336 17954 9364
rect 18050 9344 18106 9353
rect 17592 9104 17644 9110
rect 17590 9072 17592 9081
rect 17644 9072 17646 9081
rect 17590 9007 17646 9016
rect 17880 8922 17908 9336
rect 18050 9279 18106 9288
rect 18064 9042 18092 9279
rect 18156 9042 18184 9646
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18248 9092 18276 9590
rect 18340 9450 18368 10066
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18328 9104 18380 9110
rect 18248 9064 18328 9092
rect 18328 9046 18380 9052
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 17788 8894 17908 8922
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17682 8800 17738 8809
rect 17604 8498 17632 8774
rect 17682 8735 17738 8744
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17512 8214 17632 8242
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17512 6186 17540 6802
rect 17604 6769 17632 8214
rect 17696 8090 17724 8735
rect 17788 8634 17816 8894
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17880 8090 17908 8774
rect 17972 8430 18000 8910
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 18248 7993 18276 8570
rect 18234 7984 18290 7993
rect 18144 7948 18196 7954
rect 18234 7919 18290 7928
rect 18144 7890 18196 7896
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17696 7342 17724 7822
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17590 6760 17646 6769
rect 17590 6695 17646 6704
rect 17696 6662 17724 7278
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17500 6180 17552 6186
rect 17500 6122 17552 6128
rect 17512 5710 17540 6122
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17512 5166 17540 5510
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17052 3754 17080 3878
rect 17052 3738 17264 3754
rect 17052 3732 17276 3738
rect 17052 3726 17224 3732
rect 17224 3674 17276 3680
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17222 3632 17278 3641
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 16868 1970 16896 2450
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 16856 1760 16908 1766
rect 16856 1702 16908 1708
rect 16868 1562 16896 1702
rect 16304 1556 16356 1562
rect 16304 1498 16356 1504
rect 16396 1556 16448 1562
rect 16396 1498 16448 1504
rect 16856 1556 16908 1562
rect 16856 1498 16908 1504
rect 16304 1420 16356 1426
rect 16304 1362 16356 1368
rect 7840 808 7892 814
rect 7840 750 7892 756
rect 10600 808 10652 814
rect 10600 750 10652 756
rect 12348 808 12400 814
rect 12348 750 12400 756
rect 13176 808 13228 814
rect 13176 750 13228 756
rect 13728 808 13780 814
rect 13728 750 13780 756
rect 14648 808 14700 814
rect 14648 750 14700 756
rect 16212 808 16264 814
rect 16212 750 16264 756
rect 15660 740 15712 746
rect 15660 682 15712 688
rect 8102 572 8410 581
rect 8102 570 8108 572
rect 8164 570 8188 572
rect 8244 570 8268 572
rect 8324 570 8348 572
rect 8404 570 8410 572
rect 8164 518 8166 570
rect 8346 518 8348 570
rect 8102 516 8108 518
rect 8164 516 8188 518
rect 8244 516 8268 518
rect 8324 516 8348 518
rect 8404 516 8410 518
rect 8102 507 8410 516
rect 15672 490 15700 682
rect 15807 572 16115 581
rect 15807 570 15813 572
rect 15869 570 15893 572
rect 15949 570 15973 572
rect 16029 570 16053 572
rect 16109 570 16115 572
rect 15869 518 15871 570
rect 16051 518 16053 570
rect 15807 516 15813 518
rect 15869 516 15893 518
rect 15949 516 15973 518
rect 16029 516 16053 518
rect 16109 516 16115 518
rect 15807 507 16115 516
rect 15488 462 15700 490
rect 15488 400 15516 462
rect 16316 406 16344 1362
rect 17144 1018 17172 3606
rect 17328 3618 17356 3946
rect 17512 3738 17540 4014
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17278 3590 17356 3618
rect 17222 3567 17278 3576
rect 17592 1828 17644 1834
rect 17592 1770 17644 1776
rect 17604 1562 17632 1770
rect 17592 1556 17644 1562
rect 17592 1498 17644 1504
rect 17500 1420 17552 1426
rect 17420 1380 17500 1408
rect 17132 1012 17184 1018
rect 17132 954 17184 960
rect 16764 740 16816 746
rect 16764 682 16816 688
rect 16120 400 16172 406
rect 16304 400 16356 406
rect 16776 400 16804 682
rect 17420 400 17448 1380
rect 17500 1362 17552 1368
rect 17604 1290 17632 1498
rect 17592 1284 17644 1290
rect 17592 1226 17644 1232
rect 17696 796 17724 6598
rect 17788 6186 17816 6802
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17880 6322 17908 6598
rect 17972 6497 18000 6598
rect 17958 6488 18014 6497
rect 17958 6423 18014 6432
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17866 6216 17922 6225
rect 17776 6180 17828 6186
rect 17866 6151 17922 6160
rect 17776 6122 17828 6128
rect 17788 1562 17816 6122
rect 17880 5574 17908 6151
rect 18156 6118 18184 7890
rect 18340 7478 18368 8910
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 18340 7002 18368 7414
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 18432 5234 18460 11494
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 9654 18552 10406
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 18512 9104 18564 9110
rect 18510 9072 18512 9081
rect 18564 9072 18566 9081
rect 18510 9007 18566 9016
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18524 8401 18552 8774
rect 18510 8392 18566 8401
rect 18510 8327 18566 8336
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18524 6866 18552 7890
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18524 5642 18552 6190
rect 18512 5636 18564 5642
rect 18512 5578 18564 5584
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18064 4593 18092 4626
rect 18050 4584 18106 4593
rect 18050 4519 18106 4528
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18340 4282 18368 4422
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17972 2650 18000 3946
rect 18064 3398 18092 4218
rect 18432 3466 18460 4422
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18248 2106 18276 2450
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 17972 1986 18000 2042
rect 17972 1958 18092 1986
rect 17960 1896 18012 1902
rect 17960 1838 18012 1844
rect 17972 1562 18000 1838
rect 18064 1562 18092 1958
rect 18524 1562 18552 5578
rect 18616 4826 18644 11698
rect 18708 11150 18736 12838
rect 18984 12730 19012 19638
rect 19338 19600 19394 20000
rect 19982 19600 20038 20000
rect 20088 19638 20300 19666
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19260 17814 19288 18022
rect 19248 17808 19300 17814
rect 19248 17750 19300 17756
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 19260 16998 19288 17478
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19260 16726 19288 16934
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19076 15706 19104 15846
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 19076 15094 19104 15302
rect 19064 15088 19116 15094
rect 19064 15030 19116 15036
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19076 14414 19104 14894
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19168 13462 19196 16390
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19260 15706 19288 15846
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19352 15586 19380 19600
rect 19996 19530 20024 19600
rect 20088 19530 20116 19638
rect 19996 19502 20116 19530
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19660 18524 19968 18533
rect 19660 18522 19666 18524
rect 19722 18522 19746 18524
rect 19802 18522 19826 18524
rect 19882 18522 19906 18524
rect 19962 18522 19968 18524
rect 19722 18470 19724 18522
rect 19904 18470 19906 18522
rect 19660 18468 19666 18470
rect 19722 18468 19746 18470
rect 19802 18468 19826 18470
rect 19882 18468 19906 18470
rect 19962 18468 19968 18470
rect 19660 18459 19968 18468
rect 19996 18290 20024 18566
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19536 17338 19564 17478
rect 19660 17436 19968 17445
rect 19660 17434 19666 17436
rect 19722 17434 19746 17436
rect 19802 17434 19826 17436
rect 19882 17434 19906 17436
rect 19962 17434 19968 17436
rect 19722 17382 19724 17434
rect 19904 17382 19906 17434
rect 19660 17380 19666 17382
rect 19722 17380 19746 17382
rect 19802 17380 19826 17382
rect 19882 17380 19906 17382
rect 19962 17380 19968 17382
rect 19660 17371 19968 17380
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19536 17202 19564 17274
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19996 17134 20024 17478
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 19444 16046 19472 16458
rect 19660 16348 19968 16357
rect 19660 16346 19666 16348
rect 19722 16346 19746 16348
rect 19802 16346 19826 16348
rect 19882 16346 19906 16348
rect 19962 16346 19968 16348
rect 19722 16294 19724 16346
rect 19904 16294 19906 16346
rect 19660 16292 19666 16294
rect 19722 16292 19746 16294
rect 19802 16292 19826 16294
rect 19882 16292 19906 16294
rect 19962 16292 19968 16294
rect 19660 16283 19968 16292
rect 19996 16182 20024 16458
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19996 15706 20024 15846
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19352 15558 19564 15586
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19352 14958 19380 15438
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19352 14550 19380 14894
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19430 14376 19486 14385
rect 19430 14311 19432 14320
rect 19484 14311 19486 14320
rect 19432 14282 19484 14288
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19156 13456 19208 13462
rect 19156 13398 19208 13404
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19076 12986 19104 13126
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19168 12850 19196 13194
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19260 12782 19288 13670
rect 19352 13394 19380 13670
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19338 13288 19394 13297
rect 19338 13223 19394 13232
rect 19248 12776 19300 12782
rect 18788 12708 18840 12714
rect 18984 12702 19196 12730
rect 19248 12718 19300 12724
rect 18840 12668 18920 12696
rect 18788 12650 18840 12656
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18800 12073 18828 12378
rect 18786 12064 18842 12073
rect 18786 11999 18842 12008
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18800 10810 18828 11999
rect 18892 11801 18920 12668
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18878 11792 18934 11801
rect 18878 11727 18934 11736
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18892 10849 18920 11630
rect 18984 11150 19012 12582
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 19076 11898 19104 12310
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19062 11792 19118 11801
rect 19168 11762 19196 12702
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19260 12374 19288 12582
rect 19352 12442 19380 13223
rect 19444 13190 19472 13330
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19062 11727 19118 11736
rect 19156 11756 19208 11762
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18972 11008 19024 11014
rect 18972 10950 19024 10956
rect 18878 10840 18934 10849
rect 18788 10804 18840 10810
rect 18878 10775 18934 10784
rect 18788 10746 18840 10752
rect 18694 9616 18750 9625
rect 18694 9551 18750 9560
rect 18708 9110 18736 9551
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18708 7750 18736 8910
rect 18800 7954 18828 10746
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18800 6322 18828 7686
rect 18892 6798 18920 9930
rect 18984 8294 19012 10950
rect 19076 8838 19104 11727
rect 19156 11698 19208 11704
rect 19352 11665 19380 12242
rect 19338 11656 19394 11665
rect 19338 11591 19394 11600
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19168 11286 19196 11494
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 19168 8650 19196 11086
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19260 9897 19288 10610
rect 19246 9888 19302 9897
rect 19246 9823 19302 9832
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19076 8622 19196 8650
rect 19076 8430 19104 8622
rect 19154 8528 19210 8537
rect 19154 8463 19210 8472
rect 19168 8430 19196 8463
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 19260 8090 19288 8366
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 18984 7857 19012 7958
rect 19248 7880 19300 7886
rect 18970 7848 19026 7857
rect 19248 7822 19300 7828
rect 18970 7783 19026 7792
rect 19260 7206 19288 7822
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 19064 6724 19116 6730
rect 19064 6666 19116 6672
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18800 5574 18828 6258
rect 18880 6248 18932 6254
rect 18878 6216 18880 6225
rect 18932 6216 18934 6225
rect 18878 6151 18934 6160
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18788 5568 18840 5574
rect 18788 5510 18840 5516
rect 18800 5370 18828 5510
rect 18788 5364 18840 5370
rect 18788 5306 18840 5312
rect 18892 5098 18920 5714
rect 19076 5574 19104 6666
rect 19260 5846 19288 7142
rect 19352 6322 19380 9454
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 19338 5672 19394 5681
rect 19338 5607 19394 5616
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 18880 5092 18932 5098
rect 18880 5034 18932 5040
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18708 4690 18736 4966
rect 19168 4826 19196 5102
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 18984 4729 19012 4762
rect 18970 4720 19026 4729
rect 18696 4684 18748 4690
rect 19352 4690 19380 5607
rect 19444 4826 19472 12718
rect 19536 12442 19564 15558
rect 19660 15260 19968 15269
rect 19660 15258 19666 15260
rect 19722 15258 19746 15260
rect 19802 15258 19826 15260
rect 19882 15258 19906 15260
rect 19962 15258 19968 15260
rect 19722 15206 19724 15258
rect 19904 15206 19906 15258
rect 19660 15204 19666 15206
rect 19722 15204 19746 15206
rect 19802 15204 19826 15206
rect 19882 15204 19906 15206
rect 19962 15204 19968 15206
rect 19660 15195 19968 15204
rect 19800 15088 19852 15094
rect 19800 15030 19852 15036
rect 19812 14482 19840 15030
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19660 14172 19968 14181
rect 19660 14170 19666 14172
rect 19722 14170 19746 14172
rect 19802 14170 19826 14172
rect 19882 14170 19906 14172
rect 19962 14170 19968 14172
rect 19722 14118 19724 14170
rect 19904 14118 19906 14170
rect 19660 14116 19666 14118
rect 19722 14116 19746 14118
rect 19802 14116 19826 14118
rect 19882 14116 19906 14118
rect 19962 14116 19968 14118
rect 19660 14107 19968 14116
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 19996 13977 20024 14010
rect 19982 13968 20038 13977
rect 19982 13903 20038 13912
rect 19800 13796 19852 13802
rect 19852 13756 20024 13784
rect 19800 13738 19852 13744
rect 19660 13084 19968 13093
rect 19660 13082 19666 13084
rect 19722 13082 19746 13084
rect 19802 13082 19826 13084
rect 19882 13082 19906 13084
rect 19962 13082 19968 13084
rect 19722 13030 19724 13082
rect 19904 13030 19906 13082
rect 19660 13028 19666 13030
rect 19722 13028 19746 13030
rect 19802 13028 19826 13030
rect 19882 13028 19906 13030
rect 19962 13028 19968 13030
rect 19660 13019 19968 13028
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19890 12336 19946 12345
rect 19616 12300 19668 12306
rect 19536 12260 19616 12288
rect 19536 9654 19564 12260
rect 19890 12271 19946 12280
rect 19616 12242 19668 12248
rect 19904 12170 19932 12271
rect 19892 12164 19944 12170
rect 19892 12106 19944 12112
rect 19660 11996 19968 12005
rect 19660 11994 19666 11996
rect 19722 11994 19746 11996
rect 19802 11994 19826 11996
rect 19882 11994 19906 11996
rect 19962 11994 19968 11996
rect 19722 11942 19724 11994
rect 19904 11942 19906 11994
rect 19660 11940 19666 11942
rect 19722 11940 19746 11942
rect 19802 11940 19826 11942
rect 19882 11940 19906 11942
rect 19962 11940 19968 11942
rect 19660 11931 19968 11940
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19628 11558 19656 11834
rect 19798 11792 19854 11801
rect 19798 11727 19854 11736
rect 19708 11688 19760 11694
rect 19706 11656 19708 11665
rect 19760 11656 19762 11665
rect 19812 11626 19840 11727
rect 19706 11591 19762 11600
rect 19800 11620 19852 11626
rect 19800 11562 19852 11568
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19660 10908 19968 10917
rect 19660 10906 19666 10908
rect 19722 10906 19746 10908
rect 19802 10906 19826 10908
rect 19882 10906 19906 10908
rect 19962 10906 19968 10908
rect 19722 10854 19724 10906
rect 19904 10854 19906 10906
rect 19660 10852 19666 10854
rect 19722 10852 19746 10854
rect 19802 10852 19826 10854
rect 19882 10852 19906 10854
rect 19962 10852 19968 10854
rect 19660 10843 19968 10852
rect 19890 10704 19946 10713
rect 19890 10639 19946 10648
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19800 10600 19852 10606
rect 19800 10542 19852 10548
rect 19720 10441 19748 10542
rect 19706 10432 19762 10441
rect 19706 10367 19762 10376
rect 19812 10169 19840 10542
rect 19798 10160 19854 10169
rect 19798 10095 19854 10104
rect 19904 9908 19932 10639
rect 19996 10130 20024 13756
rect 20088 13326 20116 14010
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20180 13394 20208 13670
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20272 13274 20300 19638
rect 20626 19600 20682 20000
rect 27710 19600 27766 20000
rect 28354 19600 28410 20000
rect 20444 17264 20496 17270
rect 20444 17206 20496 17212
rect 20456 16726 20484 17206
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20548 16046 20576 16186
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20456 14521 20484 14554
rect 20442 14512 20498 14521
rect 20442 14447 20498 14456
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20352 13796 20404 13802
rect 20352 13738 20404 13744
rect 20364 13433 20392 13738
rect 20350 13424 20406 13433
rect 20350 13359 20406 13368
rect 20088 12782 20116 13262
rect 20272 13246 20392 13274
rect 20166 12880 20222 12889
rect 20166 12815 20222 12824
rect 20180 12782 20208 12815
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20088 12434 20116 12718
rect 20260 12708 20312 12714
rect 20260 12650 20312 12656
rect 20088 12406 20208 12434
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 20088 11801 20116 12106
rect 20074 11792 20130 11801
rect 20074 11727 20130 11736
rect 20074 11384 20130 11393
rect 20074 11319 20076 11328
rect 20128 11319 20130 11328
rect 20076 11290 20128 11296
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 20088 10606 20116 10950
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19904 9880 20024 9908
rect 19660 9820 19968 9829
rect 19660 9818 19666 9820
rect 19722 9818 19746 9820
rect 19802 9818 19826 9820
rect 19882 9818 19906 9820
rect 19962 9818 19968 9820
rect 19722 9766 19724 9818
rect 19904 9766 19906 9818
rect 19660 9764 19666 9766
rect 19722 9764 19746 9766
rect 19802 9764 19826 9766
rect 19882 9764 19906 9766
rect 19962 9764 19968 9766
rect 19660 9755 19968 9764
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19536 8498 19564 9386
rect 19720 9178 19748 9590
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19996 9110 20024 9880
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 19984 9104 20036 9110
rect 19890 9072 19946 9081
rect 19984 9046 20036 9052
rect 19890 9007 19946 9016
rect 19904 8838 19932 9007
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19660 8732 19968 8741
rect 19660 8730 19666 8732
rect 19722 8730 19746 8732
rect 19802 8730 19826 8732
rect 19882 8730 19906 8732
rect 19962 8730 19968 8732
rect 19722 8678 19724 8730
rect 19904 8678 19906 8730
rect 19660 8676 19666 8678
rect 19722 8676 19746 8678
rect 19802 8676 19826 8678
rect 19882 8676 19906 8678
rect 19962 8676 19968 8678
rect 19660 8667 19968 8676
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19892 8492 19944 8498
rect 19892 8434 19944 8440
rect 19536 6118 19564 8434
rect 19628 8090 19656 8434
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19812 8090 19840 8366
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19708 8016 19760 8022
rect 19706 7984 19708 7993
rect 19760 7984 19762 7993
rect 19706 7919 19762 7928
rect 19904 7732 19932 8434
rect 19996 7886 20024 8570
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19904 7704 20024 7732
rect 19660 7644 19968 7653
rect 19660 7642 19666 7644
rect 19722 7642 19746 7644
rect 19802 7642 19826 7644
rect 19882 7642 19906 7644
rect 19962 7642 19968 7644
rect 19722 7590 19724 7642
rect 19904 7590 19906 7642
rect 19660 7588 19666 7590
rect 19722 7588 19746 7590
rect 19802 7588 19826 7590
rect 19882 7588 19906 7590
rect 19962 7588 19968 7590
rect 19660 7579 19968 7588
rect 19708 6928 19760 6934
rect 19706 6896 19708 6905
rect 19760 6896 19762 6905
rect 19706 6831 19762 6840
rect 19660 6556 19968 6565
rect 19660 6554 19666 6556
rect 19722 6554 19746 6556
rect 19802 6554 19826 6556
rect 19882 6554 19906 6556
rect 19962 6554 19968 6556
rect 19722 6502 19724 6554
rect 19904 6502 19906 6554
rect 19660 6500 19666 6502
rect 19722 6500 19746 6502
rect 19802 6500 19826 6502
rect 19882 6500 19906 6502
rect 19962 6500 19968 6502
rect 19660 6491 19968 6500
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19536 5370 19564 6054
rect 19890 5944 19946 5953
rect 19812 5902 19890 5930
rect 19812 5846 19840 5902
rect 19996 5914 20024 7704
rect 19890 5879 19946 5888
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 19800 5840 19852 5846
rect 19892 5840 19944 5846
rect 19800 5782 19852 5788
rect 19890 5808 19892 5817
rect 19944 5808 19946 5817
rect 19890 5743 19946 5752
rect 19614 5672 19670 5681
rect 19614 5607 19616 5616
rect 19668 5607 19670 5616
rect 19616 5578 19668 5584
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19660 5468 19968 5477
rect 19660 5466 19666 5468
rect 19722 5466 19746 5468
rect 19802 5466 19826 5468
rect 19882 5466 19906 5468
rect 19962 5466 19968 5468
rect 19722 5414 19724 5466
rect 19904 5414 19906 5466
rect 19660 5412 19666 5414
rect 19722 5412 19746 5414
rect 19802 5412 19826 5414
rect 19882 5412 19906 5414
rect 19962 5412 19968 5414
rect 19660 5403 19968 5412
rect 19996 5370 20024 5510
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19536 5234 19564 5306
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 18970 4655 19026 4664
rect 19340 4684 19392 4690
rect 18696 4626 18748 4632
rect 19340 4626 19392 4632
rect 19062 4584 19118 4593
rect 19996 4554 20024 5102
rect 19062 4519 19118 4528
rect 19984 4548 20036 4554
rect 18878 4448 18934 4457
rect 18878 4383 18934 4392
rect 18892 3738 18920 4383
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 19076 3670 19104 4519
rect 19984 4490 20036 4496
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19352 3738 19380 4422
rect 19660 4380 19968 4389
rect 19660 4378 19666 4380
rect 19722 4378 19746 4380
rect 19802 4378 19826 4380
rect 19882 4378 19906 4380
rect 19962 4378 19968 4380
rect 19722 4326 19724 4378
rect 19904 4326 19906 4378
rect 19660 4324 19666 4326
rect 19722 4324 19746 4326
rect 19802 4324 19826 4326
rect 19882 4324 19906 4326
rect 19962 4324 19968 4326
rect 19660 4315 19968 4324
rect 20088 4146 20116 9454
rect 20180 8498 20208 12406
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20180 6730 20208 7686
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 20180 4826 20208 6190
rect 20272 5370 20300 12650
rect 20364 12073 20392 13246
rect 20456 13190 20484 13806
rect 20548 13394 20576 14962
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20548 13002 20576 13194
rect 20456 12974 20576 13002
rect 20350 12064 20406 12073
rect 20350 11999 20406 12008
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20364 10810 20392 11630
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20456 10198 20484 12974
rect 20640 12850 20668 19600
rect 23512 19068 23820 19077
rect 23512 19066 23518 19068
rect 23574 19066 23598 19068
rect 23654 19066 23678 19068
rect 23734 19066 23758 19068
rect 23814 19066 23820 19068
rect 23574 19014 23576 19066
rect 23756 19014 23758 19066
rect 23512 19012 23518 19014
rect 23574 19012 23598 19014
rect 23654 19012 23678 19014
rect 23734 19012 23758 19014
rect 23814 19012 23820 19014
rect 23512 19003 23820 19012
rect 27724 18834 27752 19600
rect 28368 18834 28396 19600
rect 31666 19136 31722 19145
rect 31217 19068 31525 19077
rect 31666 19071 31722 19080
rect 31217 19066 31223 19068
rect 31279 19066 31303 19068
rect 31359 19066 31383 19068
rect 31439 19066 31463 19068
rect 31519 19066 31525 19068
rect 31279 19014 31281 19066
rect 31461 19014 31463 19066
rect 31217 19012 31223 19014
rect 31279 19012 31303 19014
rect 31359 19012 31383 19014
rect 31439 19012 31463 19014
rect 31519 19012 31525 19014
rect 31217 19003 31525 19012
rect 31680 18834 31708 19071
rect 20812 18828 20864 18834
rect 20812 18770 20864 18776
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 27712 18828 27764 18834
rect 27712 18770 27764 18776
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 31668 18828 31720 18834
rect 31668 18770 31720 18776
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20732 16776 20760 18566
rect 20824 18426 20852 18770
rect 21008 18426 21036 18770
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 22296 18154 22324 18566
rect 22756 18426 22784 18566
rect 23032 18426 23060 18566
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 23216 18222 23244 18770
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 24032 18624 24084 18630
rect 24032 18566 24084 18572
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 22284 18148 22336 18154
rect 22284 18090 22336 18096
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22388 17814 22416 18022
rect 22848 17814 22876 18158
rect 23512 17980 23820 17989
rect 23512 17978 23518 17980
rect 23574 17978 23598 17980
rect 23654 17978 23678 17980
rect 23734 17978 23758 17980
rect 23814 17978 23820 17980
rect 23574 17926 23576 17978
rect 23756 17926 23758 17978
rect 23512 17924 23518 17926
rect 23574 17924 23598 17926
rect 23654 17924 23678 17926
rect 23734 17924 23758 17926
rect 23814 17924 23820 17926
rect 23512 17915 23820 17924
rect 22376 17808 22428 17814
rect 22376 17750 22428 17756
rect 22836 17808 22888 17814
rect 22836 17750 22888 17756
rect 21916 17740 21968 17746
rect 21916 17682 21968 17688
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 21100 16794 21128 16934
rect 21088 16788 21140 16794
rect 20732 16748 20852 16776
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20732 16182 20760 16594
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20536 12368 20588 12374
rect 20536 12310 20588 12316
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20548 9722 20576 12310
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20534 9616 20590 9625
rect 20456 9574 20534 9602
rect 20456 9518 20484 9574
rect 20534 9551 20590 9560
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20272 4758 20300 5102
rect 20260 4752 20312 4758
rect 20260 4694 20312 4700
rect 20364 4690 20392 9386
rect 20456 9217 20484 9454
rect 20442 9208 20498 9217
rect 20548 9178 20576 9454
rect 20442 9143 20498 9152
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20640 9042 20668 12582
rect 20732 9500 20760 15302
rect 20824 13802 20852 16748
rect 21088 16730 21140 16736
rect 20996 15972 21048 15978
rect 20996 15914 21048 15920
rect 21008 15706 21036 15914
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20916 15042 20944 15302
rect 21008 15162 21036 15302
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20916 15014 21036 15042
rect 21008 14958 21036 15014
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 20902 14376 20958 14385
rect 20902 14311 20958 14320
rect 20916 13870 20944 14311
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21008 13870 21036 14010
rect 21100 13870 21128 14214
rect 21192 14074 21220 14826
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21178 13968 21234 13977
rect 21178 13903 21234 13912
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 20812 13796 20864 13802
rect 20812 13738 20864 13744
rect 21192 13734 21220 13903
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20916 12238 20944 12718
rect 21192 12458 21220 13330
rect 21008 12430 21220 12458
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20824 11665 20852 11834
rect 20916 11694 20944 12174
rect 20904 11688 20956 11694
rect 20810 11656 20866 11665
rect 20904 11630 20956 11636
rect 20810 11591 20866 11600
rect 20810 11384 20866 11393
rect 20810 11319 20866 11328
rect 20824 11082 20852 11319
rect 21008 11218 21036 12430
rect 21284 11370 21312 17478
rect 21928 17338 21956 17682
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 21916 17332 21968 17338
rect 21916 17274 21968 17280
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21560 16658 21588 16934
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21468 16046 21496 16390
rect 21928 16046 21956 17274
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 22020 16114 22048 16390
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 21928 15570 21956 15982
rect 22020 15638 22048 16050
rect 22388 16046 22416 16594
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 22008 15632 22060 15638
rect 22008 15574 22060 15580
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21376 14226 21404 14758
rect 21928 14618 21956 15506
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21640 14476 21692 14482
rect 21640 14418 21692 14424
rect 21376 14198 21496 14226
rect 21362 13968 21418 13977
rect 21362 13903 21418 13912
rect 21376 13870 21404 13903
rect 21468 13870 21496 14198
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21456 13864 21508 13870
rect 21548 13864 21600 13870
rect 21456 13806 21508 13812
rect 21546 13832 21548 13841
rect 21600 13832 21602 13841
rect 21364 13320 21416 13326
rect 21362 13288 21364 13297
rect 21416 13288 21418 13297
rect 21362 13223 21418 13232
rect 21468 12374 21496 13806
rect 21546 13767 21602 13776
rect 21560 13394 21588 13767
rect 21652 13462 21680 14418
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 21744 13870 21772 14010
rect 21732 13864 21784 13870
rect 21732 13806 21784 13812
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21744 13326 21772 13806
rect 22008 13796 22060 13802
rect 22112 13784 22140 14758
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22296 14074 22324 14214
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 22060 13756 22140 13784
rect 22008 13738 22060 13744
rect 22388 13734 22416 13942
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21652 12442 21680 13126
rect 21836 12986 21864 13330
rect 22204 13297 22232 13330
rect 22190 13288 22246 13297
rect 22190 13223 22246 13232
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 21640 12436 21692 12442
rect 21560 12396 21640 12424
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21192 11342 21312 11370
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 21008 10130 21036 11154
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 20812 9648 20864 9654
rect 21192 9636 21220 11342
rect 21272 11280 21324 11286
rect 21272 11222 21324 11228
rect 21284 10674 21312 11222
rect 21468 11014 21496 11630
rect 21456 11008 21508 11014
rect 21456 10950 21508 10956
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21284 10266 21312 10610
rect 21560 10538 21588 12396
rect 21640 12378 21692 12384
rect 21638 12064 21694 12073
rect 21638 11999 21694 12008
rect 21652 11762 21680 11999
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21548 10532 21600 10538
rect 21548 10474 21600 10480
rect 21732 10532 21784 10538
rect 21732 10474 21784 10480
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21284 9722 21312 10202
rect 21546 10160 21602 10169
rect 21744 10130 21772 10474
rect 21546 10095 21602 10104
rect 21640 10124 21692 10130
rect 21560 9994 21588 10095
rect 21640 10066 21692 10072
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21362 9752 21418 9761
rect 21272 9716 21324 9722
rect 21652 9722 21680 10066
rect 21362 9687 21418 9696
rect 21640 9716 21692 9722
rect 21272 9658 21324 9664
rect 20864 9608 21220 9636
rect 20812 9590 20864 9596
rect 20904 9512 20956 9518
rect 20732 9472 20904 9500
rect 20904 9454 20956 9460
rect 21088 9444 21140 9450
rect 21008 9404 21088 9432
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20456 8809 20484 8910
rect 20442 8800 20498 8809
rect 20442 8735 20498 8744
rect 20442 8256 20498 8265
rect 20442 8191 20498 8200
rect 20626 8256 20682 8265
rect 20626 8191 20682 8200
rect 20456 5658 20484 8191
rect 20536 8084 20588 8090
rect 20640 8072 20668 8191
rect 20588 8044 20668 8072
rect 20536 8026 20588 8032
rect 20548 7002 20576 8026
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20824 6254 20852 7142
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20456 5630 20668 5658
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20456 5370 20484 5510
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20640 5234 20668 5630
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20732 5273 20760 5306
rect 20718 5264 20774 5273
rect 20628 5228 20680 5234
rect 20718 5199 20774 5208
rect 20628 5170 20680 5176
rect 20824 5030 20852 5306
rect 21008 5302 21036 9404
rect 21088 9386 21140 9392
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 20996 5296 21048 5302
rect 20996 5238 21048 5244
rect 21008 5166 21036 5238
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 21100 4690 21128 8570
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21284 7478 21312 7754
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 21192 6730 21220 7278
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 21376 6610 21404 9687
rect 21640 9658 21692 9664
rect 21732 8628 21784 8634
rect 21836 8616 21864 12922
rect 22008 11824 22060 11830
rect 22006 11792 22008 11801
rect 22060 11792 22062 11801
rect 22296 11778 22324 13670
rect 22480 12434 22508 13806
rect 22572 13802 22600 14418
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22664 14074 22692 14214
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22560 13796 22612 13802
rect 22560 13738 22612 13744
rect 22560 12776 22612 12782
rect 22560 12718 22612 12724
rect 22388 12406 22508 12434
rect 22388 12102 22416 12406
rect 22572 12186 22600 12718
rect 22756 12714 22784 15030
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22940 14385 22968 14418
rect 22926 14376 22982 14385
rect 22926 14311 22982 14320
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22848 14074 22876 14214
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22834 13560 22890 13569
rect 22834 13495 22836 13504
rect 22888 13495 22890 13504
rect 22836 13466 22888 13472
rect 22744 12708 22796 12714
rect 22744 12650 22796 12656
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22848 12306 22876 12582
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 22572 12170 22692 12186
rect 22572 12164 22704 12170
rect 22572 12158 22652 12164
rect 22652 12106 22704 12112
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22296 11750 22692 11778
rect 22006 11727 22062 11736
rect 22560 11688 22612 11694
rect 22560 11630 22612 11636
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 22020 10266 22048 11154
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22112 10266 22140 10746
rect 22204 10674 22232 11222
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22192 10464 22244 10470
rect 22296 10452 22324 11494
rect 22572 11218 22600 11630
rect 22560 11212 22612 11218
rect 22560 11154 22612 11160
rect 22244 10424 22324 10452
rect 22192 10406 22244 10412
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21784 8588 21864 8616
rect 21732 8570 21784 8576
rect 21652 8214 21864 8242
rect 21652 8090 21680 8214
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 21652 7750 21680 8026
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21744 7546 21772 8026
rect 21836 8022 21864 8214
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21836 7546 21864 7958
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21732 7540 21784 7546
rect 21732 7482 21784 7488
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21468 7342 21496 7482
rect 21928 7410 21956 10134
rect 22204 10130 22232 10406
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 22560 10124 22612 10130
rect 22560 10066 22612 10072
rect 22192 9512 22244 9518
rect 22296 9466 22324 10066
rect 22572 9722 22600 10066
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22374 9616 22430 9625
rect 22430 9574 22508 9602
rect 22374 9551 22430 9560
rect 22480 9518 22508 9574
rect 22468 9512 22520 9518
rect 22244 9460 22416 9466
rect 22192 9454 22416 9460
rect 22468 9454 22520 9460
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22100 9444 22152 9450
rect 22204 9438 22416 9454
rect 22100 9386 22152 9392
rect 22112 9178 22140 9386
rect 22388 9382 22416 9438
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22376 9376 22428 9382
rect 22376 9318 22428 9324
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22008 8900 22060 8906
rect 22008 8842 22060 8848
rect 22020 8634 22048 8842
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 22112 8362 22140 8978
rect 22296 8838 22324 9318
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22112 8090 22140 8298
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 22204 7546 22232 7890
rect 22284 7744 22336 7750
rect 22388 7732 22416 9318
rect 22572 9042 22600 9454
rect 22560 9036 22612 9042
rect 22560 8978 22612 8984
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22480 8430 22508 8910
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22572 8090 22600 8978
rect 22664 8566 22692 11750
rect 22756 11393 22784 12242
rect 22940 12220 22968 14311
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 23032 12646 23060 13806
rect 23020 12640 23072 12646
rect 23020 12582 23072 12588
rect 23032 12374 23060 12582
rect 23124 12374 23152 16934
rect 23216 14550 23244 17478
rect 23512 16892 23820 16901
rect 23512 16890 23518 16892
rect 23574 16890 23598 16892
rect 23654 16890 23678 16892
rect 23734 16890 23758 16892
rect 23814 16890 23820 16892
rect 23574 16838 23576 16890
rect 23756 16838 23758 16890
rect 23512 16836 23518 16838
rect 23574 16836 23598 16838
rect 23654 16836 23678 16838
rect 23734 16836 23758 16838
rect 23814 16836 23820 16838
rect 23512 16827 23820 16836
rect 23664 16652 23716 16658
rect 23860 16640 23888 17478
rect 23716 16612 23888 16640
rect 23664 16594 23716 16600
rect 23676 16046 23704 16594
rect 23940 16176 23992 16182
rect 23940 16118 23992 16124
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 23848 15904 23900 15910
rect 23848 15846 23900 15852
rect 23512 15804 23820 15813
rect 23512 15802 23518 15804
rect 23574 15802 23598 15804
rect 23654 15802 23678 15804
rect 23734 15802 23758 15804
rect 23814 15802 23820 15804
rect 23574 15750 23576 15802
rect 23756 15750 23758 15802
rect 23512 15748 23518 15750
rect 23574 15748 23598 15750
rect 23654 15748 23678 15750
rect 23734 15748 23758 15750
rect 23814 15748 23820 15750
rect 23512 15739 23820 15748
rect 23860 15706 23888 15846
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 23952 15450 23980 16118
rect 23860 15422 23980 15450
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23204 14544 23256 14550
rect 23204 14486 23256 14492
rect 23308 14362 23336 14962
rect 23512 14716 23820 14725
rect 23512 14714 23518 14716
rect 23574 14714 23598 14716
rect 23654 14714 23678 14716
rect 23734 14714 23758 14716
rect 23814 14714 23820 14716
rect 23574 14662 23576 14714
rect 23756 14662 23758 14714
rect 23512 14660 23518 14662
rect 23574 14660 23598 14662
rect 23654 14660 23678 14662
rect 23734 14660 23758 14662
rect 23814 14660 23820 14662
rect 23512 14651 23820 14660
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23216 14334 23336 14362
rect 23480 14408 23532 14414
rect 23676 14385 23704 14486
rect 23480 14350 23532 14356
rect 23662 14376 23718 14385
rect 23216 13734 23244 14334
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23308 14074 23336 14214
rect 23492 14074 23520 14350
rect 23662 14311 23718 14320
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23492 13841 23520 14010
rect 23570 13968 23626 13977
rect 23570 13903 23626 13912
rect 23584 13870 23612 13903
rect 23572 13864 23624 13870
rect 23478 13832 23534 13841
rect 23572 13806 23624 13812
rect 23860 13802 23888 15422
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23952 14958 23980 15302
rect 23940 14952 23992 14958
rect 23940 14894 23992 14900
rect 23938 14512 23994 14521
rect 24044 14482 24072 18566
rect 24308 18216 24360 18222
rect 24308 18158 24360 18164
rect 24952 18216 25004 18222
rect 24952 18158 25004 18164
rect 24320 17882 24348 18158
rect 24964 17882 24992 18158
rect 24308 17876 24360 17882
rect 24308 17818 24360 17824
rect 24952 17876 25004 17882
rect 24952 17818 25004 17824
rect 24308 17740 24360 17746
rect 24308 17682 24360 17688
rect 24320 17066 24348 17682
rect 25240 17678 25268 18702
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 27365 18524 27673 18533
rect 27365 18522 27371 18524
rect 27427 18522 27451 18524
rect 27507 18522 27531 18524
rect 27587 18522 27611 18524
rect 27667 18522 27673 18524
rect 27427 18470 27429 18522
rect 27609 18470 27611 18522
rect 27365 18468 27371 18470
rect 27427 18468 27451 18470
rect 27507 18468 27531 18470
rect 27587 18468 27611 18470
rect 27667 18468 27673 18470
rect 27365 18459 27673 18468
rect 31036 18465 31064 18566
rect 31022 18456 31078 18465
rect 31022 18391 31078 18400
rect 31217 17980 31525 17989
rect 31217 17978 31223 17980
rect 31279 17978 31303 17980
rect 31359 17978 31383 17980
rect 31439 17978 31463 17980
rect 31519 17978 31525 17980
rect 31279 17926 31281 17978
rect 31461 17926 31463 17978
rect 31217 17924 31223 17926
rect 31279 17924 31303 17926
rect 31359 17924 31383 17926
rect 31439 17924 31463 17926
rect 31519 17924 31525 17926
rect 31217 17915 31525 17924
rect 25320 17740 25372 17746
rect 25320 17682 25372 17688
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 25332 17338 25360 17682
rect 25320 17332 25372 17338
rect 25320 17274 25372 17280
rect 25332 17202 25360 17274
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 25412 17128 25464 17134
rect 25412 17070 25464 17076
rect 24308 17060 24360 17066
rect 24308 17002 24360 17008
rect 24320 16658 24348 17002
rect 25424 16658 25452 17070
rect 25608 16998 25636 17682
rect 25688 17128 25740 17134
rect 25688 17070 25740 17076
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25700 16794 25728 17070
rect 26160 17066 26188 17682
rect 27365 17436 27673 17445
rect 27365 17434 27371 17436
rect 27427 17434 27451 17436
rect 27507 17434 27531 17436
rect 27587 17434 27611 17436
rect 27667 17434 27673 17436
rect 27427 17382 27429 17434
rect 27609 17382 27611 17434
rect 27365 17380 27371 17382
rect 27427 17380 27451 17382
rect 27507 17380 27531 17382
rect 27587 17380 27611 17382
rect 27667 17380 27673 17382
rect 27365 17371 27673 17380
rect 27068 17128 27120 17134
rect 27068 17070 27120 17076
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 25688 16788 25740 16794
rect 25688 16730 25740 16736
rect 24308 16652 24360 16658
rect 24308 16594 24360 16600
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 24952 16448 25004 16454
rect 24952 16390 25004 16396
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24308 15564 24360 15570
rect 24308 15506 24360 15512
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 24216 15496 24268 15502
rect 24216 15438 24268 15444
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 23938 14447 23940 14456
rect 23992 14447 23994 14456
rect 24032 14476 24084 14482
rect 23940 14418 23992 14424
rect 24032 14418 24084 14424
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 23478 13767 23534 13776
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 23204 13728 23256 13734
rect 23204 13670 23256 13676
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23020 12368 23072 12374
rect 23020 12310 23072 12316
rect 23112 12368 23164 12374
rect 23112 12310 23164 12316
rect 23216 12306 23244 13670
rect 23294 13560 23350 13569
rect 23400 13530 23428 13670
rect 23512 13628 23820 13637
rect 23512 13626 23518 13628
rect 23574 13626 23598 13628
rect 23654 13626 23678 13628
rect 23734 13626 23758 13628
rect 23814 13626 23820 13628
rect 23574 13574 23576 13626
rect 23756 13574 23758 13626
rect 23512 13572 23518 13574
rect 23574 13572 23598 13574
rect 23654 13572 23678 13574
rect 23734 13572 23758 13574
rect 23814 13572 23820 13574
rect 23512 13563 23820 13572
rect 23294 13495 23350 13504
rect 23388 13524 23440 13530
rect 23308 13258 23336 13495
rect 23388 13466 23440 13472
rect 23480 13320 23532 13326
rect 23478 13288 23480 13297
rect 23532 13288 23534 13297
rect 23296 13252 23348 13258
rect 23478 13223 23534 13232
rect 23296 13194 23348 13200
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23400 12782 23428 12922
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23204 12300 23256 12306
rect 23204 12242 23256 12248
rect 22940 12192 23152 12220
rect 22836 12164 22888 12170
rect 22836 12106 22888 12112
rect 22848 11830 22876 12106
rect 22836 11824 22888 11830
rect 22836 11766 22888 11772
rect 22836 11552 22888 11558
rect 22836 11494 22888 11500
rect 22742 11384 22798 11393
rect 22742 11319 22798 11328
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 22756 10266 22784 11154
rect 22848 10606 22876 11494
rect 23018 11384 23074 11393
rect 23018 11319 23074 11328
rect 23032 10690 23060 11319
rect 22940 10662 23060 10690
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22848 10266 22876 10542
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22652 8560 22704 8566
rect 22940 8514 22968 10662
rect 23018 10568 23074 10577
rect 23018 10503 23074 10512
rect 22652 8502 22704 8508
rect 22756 8486 22968 8514
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22336 7704 22416 7732
rect 22284 7686 22336 7692
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22296 7426 22324 7686
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 22204 7398 22324 7426
rect 21456 7336 21508 7342
rect 21456 7278 21508 7284
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21468 6798 21496 7278
rect 21560 7206 21588 7278
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21560 7002 21588 7142
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21836 6848 21864 7278
rect 21652 6820 21864 6848
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21652 6662 21680 6820
rect 21284 6582 21404 6610
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 20352 4684 20404 4690
rect 20352 4626 20404 4632
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20180 4282 20208 4558
rect 20272 4282 20300 4558
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19628 3738 19656 4082
rect 20640 3738 20668 4422
rect 20732 4282 20760 4422
rect 20720 4276 20772 4282
rect 20720 4218 20772 4224
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 19156 3664 19208 3670
rect 19156 3606 19208 3612
rect 19984 3664 20036 3670
rect 19984 3606 20036 3612
rect 19064 3528 19116 3534
rect 19062 3496 19064 3505
rect 19116 3496 19118 3505
rect 19062 3431 19118 3440
rect 19076 3398 19104 3431
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 18984 3074 19012 3334
rect 19064 3188 19116 3194
rect 19168 3176 19196 3606
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19116 3148 19196 3176
rect 19064 3130 19116 3136
rect 19260 3074 19288 3334
rect 18984 3046 19288 3074
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 18696 1964 18748 1970
rect 18696 1906 18748 1912
rect 17776 1556 17828 1562
rect 17776 1498 17828 1504
rect 17960 1556 18012 1562
rect 17960 1498 18012 1504
rect 18052 1556 18104 1562
rect 18052 1498 18104 1504
rect 18512 1556 18564 1562
rect 18512 1498 18564 1504
rect 18236 1420 18288 1426
rect 18064 1380 18236 1408
rect 17868 808 17920 814
rect 17696 768 17868 796
rect 17868 750 17920 756
rect 18064 400 18092 1380
rect 18236 1362 18288 1368
rect 18708 882 18736 1906
rect 19064 1896 19116 1902
rect 19064 1838 19116 1844
rect 18788 1760 18840 1766
rect 18788 1702 18840 1708
rect 18800 1562 18828 1702
rect 19076 1562 19104 1838
rect 19444 1834 19472 2858
rect 19536 2650 19564 3470
rect 19660 3292 19968 3301
rect 19660 3290 19666 3292
rect 19722 3290 19746 3292
rect 19802 3290 19826 3292
rect 19882 3290 19906 3292
rect 19962 3290 19968 3292
rect 19722 3238 19724 3290
rect 19904 3238 19906 3290
rect 19660 3236 19666 3238
rect 19722 3236 19746 3238
rect 19802 3236 19826 3238
rect 19882 3236 19906 3238
rect 19962 3236 19968 3238
rect 19660 3227 19968 3236
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 19660 2204 19968 2213
rect 19660 2202 19666 2204
rect 19722 2202 19746 2204
rect 19802 2202 19826 2204
rect 19882 2202 19906 2204
rect 19962 2202 19968 2204
rect 19722 2150 19724 2202
rect 19904 2150 19906 2202
rect 19660 2148 19666 2150
rect 19722 2148 19746 2150
rect 19802 2148 19826 2150
rect 19882 2148 19906 2150
rect 19962 2148 19968 2150
rect 19660 2139 19968 2148
rect 19432 1828 19484 1834
rect 19432 1770 19484 1776
rect 19444 1562 19472 1770
rect 19524 1760 19576 1766
rect 19524 1702 19576 1708
rect 18788 1556 18840 1562
rect 18788 1498 18840 1504
rect 19064 1556 19116 1562
rect 19064 1498 19116 1504
rect 19432 1556 19484 1562
rect 19432 1498 19484 1504
rect 19536 1426 19564 1702
rect 19524 1420 19576 1426
rect 19524 1362 19576 1368
rect 18696 876 18748 882
rect 18696 818 18748 824
rect 19536 814 19564 1362
rect 19660 1116 19968 1125
rect 19660 1114 19666 1116
rect 19722 1114 19746 1116
rect 19802 1114 19826 1116
rect 19882 1114 19906 1116
rect 19962 1114 19968 1116
rect 19722 1062 19724 1114
rect 19904 1062 19906 1114
rect 19660 1060 19666 1062
rect 19722 1060 19746 1062
rect 19802 1060 19826 1062
rect 19882 1060 19906 1062
rect 19962 1060 19968 1062
rect 19660 1051 19968 1060
rect 19996 1018 20024 3606
rect 20718 3496 20774 3505
rect 20718 3431 20774 3440
rect 20732 3398 20760 3431
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20824 3194 20852 4422
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 21192 2990 21220 6122
rect 21284 3738 21312 6582
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21376 5778 21404 6190
rect 21468 5846 21496 6394
rect 21456 5840 21508 5846
rect 21456 5782 21508 5788
rect 21652 5828 21680 6598
rect 21928 6254 21956 7346
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22112 6458 22140 6734
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21732 5840 21784 5846
rect 21652 5800 21732 5828
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 21548 5772 21600 5778
rect 21652 5760 21680 5800
rect 21732 5782 21784 5788
rect 21600 5732 21680 5760
rect 21548 5714 21600 5720
rect 21376 4690 21404 5714
rect 21640 5160 21692 5166
rect 21640 5102 21692 5108
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 21652 4593 21680 5102
rect 22204 4758 22232 7398
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22296 6458 22324 6802
rect 22388 6730 22416 7278
rect 22376 6724 22428 6730
rect 22376 6666 22428 6672
rect 22664 6662 22692 7890
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 22664 6390 22692 6598
rect 22652 6384 22704 6390
rect 22652 6326 22704 6332
rect 22664 6118 22692 6326
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22388 5846 22416 6054
rect 22376 5840 22428 5846
rect 22376 5782 22428 5788
rect 22652 5568 22704 5574
rect 22652 5510 22704 5516
rect 22664 5234 22692 5510
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22756 5137 22784 8486
rect 22928 8424 22980 8430
rect 22928 8366 22980 8372
rect 22940 7886 22968 8366
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22940 7274 22968 7822
rect 22928 7268 22980 7274
rect 22928 7210 22980 7216
rect 22940 6662 22968 7210
rect 22836 6656 22888 6662
rect 22834 6624 22836 6633
rect 22928 6656 22980 6662
rect 22888 6624 22890 6633
rect 22928 6598 22980 6604
rect 22834 6559 22890 6568
rect 22926 5944 22982 5953
rect 22926 5879 22982 5888
rect 22940 5642 22968 5879
rect 23032 5794 23060 10503
rect 23124 8430 23152 12192
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 23202 11520 23258 11529
rect 23202 11455 23258 11464
rect 23216 11354 23244 11455
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23308 10441 23336 11766
rect 23294 10432 23350 10441
rect 23294 10367 23350 10376
rect 23400 10062 23428 12582
rect 23512 12540 23820 12549
rect 23512 12538 23518 12540
rect 23574 12538 23598 12540
rect 23654 12538 23678 12540
rect 23734 12538 23758 12540
rect 23814 12538 23820 12540
rect 23574 12486 23576 12538
rect 23756 12486 23758 12538
rect 23512 12484 23518 12486
rect 23574 12484 23598 12486
rect 23654 12484 23678 12486
rect 23734 12484 23758 12486
rect 23814 12484 23820 12486
rect 23512 12475 23820 12484
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23492 11694 23520 12378
rect 23572 12164 23624 12170
rect 23572 12106 23624 12112
rect 23584 11762 23612 12106
rect 23860 11762 23888 12718
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23952 11694 23980 14214
rect 24044 12306 24072 14214
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 24032 11824 24084 11830
rect 24030 11792 24032 11801
rect 24084 11792 24086 11801
rect 24030 11727 24086 11736
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 24032 11620 24084 11626
rect 24032 11562 24084 11568
rect 24044 11506 24072 11562
rect 23952 11478 24072 11506
rect 23512 11452 23820 11461
rect 23512 11450 23518 11452
rect 23574 11450 23598 11452
rect 23654 11450 23678 11452
rect 23734 11450 23758 11452
rect 23814 11450 23820 11452
rect 23574 11398 23576 11450
rect 23756 11398 23758 11450
rect 23512 11396 23518 11398
rect 23574 11396 23598 11398
rect 23654 11396 23678 11398
rect 23734 11396 23758 11398
rect 23814 11396 23820 11398
rect 23512 11387 23820 11396
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23512 10364 23820 10373
rect 23512 10362 23518 10364
rect 23574 10362 23598 10364
rect 23654 10362 23678 10364
rect 23734 10362 23758 10364
rect 23814 10362 23820 10364
rect 23574 10310 23576 10362
rect 23756 10310 23758 10362
rect 23512 10308 23518 10310
rect 23574 10308 23598 10310
rect 23654 10308 23678 10310
rect 23734 10308 23758 10310
rect 23814 10308 23820 10310
rect 23512 10299 23820 10308
rect 23860 10266 23888 10406
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23388 10056 23440 10062
rect 23202 10024 23258 10033
rect 23388 9998 23440 10004
rect 23202 9959 23204 9968
rect 23256 9959 23258 9968
rect 23204 9930 23256 9936
rect 23848 9920 23900 9926
rect 23848 9862 23900 9868
rect 23512 9276 23820 9285
rect 23512 9274 23518 9276
rect 23574 9274 23598 9276
rect 23654 9274 23678 9276
rect 23734 9274 23758 9276
rect 23814 9274 23820 9276
rect 23574 9222 23576 9274
rect 23756 9222 23758 9274
rect 23512 9220 23518 9222
rect 23574 9220 23598 9222
rect 23654 9220 23678 9222
rect 23734 9220 23758 9222
rect 23814 9220 23820 9222
rect 23512 9211 23820 9220
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23492 8634 23520 8978
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 23676 8634 23704 8842
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23112 8424 23164 8430
rect 23112 8366 23164 8372
rect 23124 8265 23152 8366
rect 23110 8256 23166 8265
rect 23110 8191 23166 8200
rect 23512 8188 23820 8197
rect 23512 8186 23518 8188
rect 23574 8186 23598 8188
rect 23654 8186 23678 8188
rect 23734 8186 23758 8188
rect 23814 8186 23820 8188
rect 23574 8134 23576 8186
rect 23756 8134 23758 8186
rect 23512 8132 23518 8134
rect 23574 8132 23598 8134
rect 23654 8132 23678 8134
rect 23734 8132 23758 8134
rect 23814 8132 23820 8134
rect 23512 8123 23820 8132
rect 23204 7200 23256 7206
rect 23204 7142 23256 7148
rect 23216 5846 23244 7142
rect 23512 7100 23820 7109
rect 23512 7098 23518 7100
rect 23574 7098 23598 7100
rect 23654 7098 23678 7100
rect 23734 7098 23758 7100
rect 23814 7098 23820 7100
rect 23574 7046 23576 7098
rect 23756 7046 23758 7098
rect 23512 7044 23518 7046
rect 23574 7044 23598 7046
rect 23654 7044 23678 7046
rect 23734 7044 23758 7046
rect 23814 7044 23820 7046
rect 23512 7035 23820 7044
rect 23860 6934 23888 9862
rect 23952 9042 23980 11478
rect 24032 9988 24084 9994
rect 24032 9930 24084 9936
rect 23940 9036 23992 9042
rect 23940 8978 23992 8984
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 23952 6322 23980 6802
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 23756 6248 23808 6254
rect 23756 6190 23808 6196
rect 23768 6100 23796 6190
rect 23768 6072 23980 6100
rect 23512 6012 23820 6021
rect 23512 6010 23518 6012
rect 23574 6010 23598 6012
rect 23654 6010 23678 6012
rect 23734 6010 23758 6012
rect 23814 6010 23820 6012
rect 23574 5958 23576 6010
rect 23756 5958 23758 6010
rect 23512 5956 23518 5958
rect 23574 5956 23598 5958
rect 23654 5956 23678 5958
rect 23734 5956 23758 5958
rect 23814 5956 23820 5958
rect 23512 5947 23820 5956
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23204 5840 23256 5846
rect 23032 5766 23152 5794
rect 23204 5782 23256 5788
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 22836 5636 22888 5642
rect 22836 5578 22888 5584
rect 22928 5636 22980 5642
rect 22928 5578 22980 5584
rect 22742 5128 22798 5137
rect 22848 5098 22876 5578
rect 22928 5296 22980 5302
rect 22928 5238 22980 5244
rect 22742 5063 22798 5072
rect 22836 5092 22888 5098
rect 22836 5034 22888 5040
rect 22192 4752 22244 4758
rect 22192 4694 22244 4700
rect 21638 4584 21694 4593
rect 21638 4519 21694 4528
rect 22848 4282 22876 5034
rect 22940 4282 22968 5238
rect 23032 4826 23060 5646
rect 23124 5302 23152 5766
rect 23112 5296 23164 5302
rect 23112 5238 23164 5244
rect 23112 5160 23164 5166
rect 23216 5148 23244 5782
rect 23296 5772 23348 5778
rect 23348 5732 23428 5760
rect 23296 5714 23348 5720
rect 23164 5120 23244 5148
rect 23112 5102 23164 5108
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23124 4826 23152 4966
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 23018 4584 23074 4593
rect 23216 4570 23244 4966
rect 23074 4542 23244 4570
rect 23018 4519 23074 4528
rect 21732 4276 21784 4282
rect 21732 4218 21784 4224
rect 22652 4276 22704 4282
rect 22836 4276 22888 4282
rect 22704 4236 22836 4264
rect 22652 4218 22704 4224
rect 22836 4218 22888 4224
rect 22928 4276 22980 4282
rect 23032 4264 23060 4519
rect 23112 4276 23164 4282
rect 23032 4236 23112 4264
rect 22928 4218 22980 4224
rect 23112 4218 23164 4224
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 21468 3194 21496 3946
rect 21548 3664 21600 3670
rect 21548 3606 21600 3612
rect 21560 3194 21588 3606
rect 21744 3398 21772 4218
rect 23124 4146 23152 4218
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 22376 4004 22428 4010
rect 22376 3946 22428 3952
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21836 3720 21864 3878
rect 21916 3732 21968 3738
rect 21836 3692 21916 3720
rect 21916 3674 21968 3680
rect 22008 3664 22060 3670
rect 22008 3606 22060 3612
rect 21732 3392 21784 3398
rect 21732 3334 21784 3340
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 20088 1970 20116 2926
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20272 2650 20300 2858
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 20180 2106 20208 2450
rect 20168 2100 20220 2106
rect 20168 2042 20220 2048
rect 20076 1964 20128 1970
rect 20076 1906 20128 1912
rect 20076 1556 20128 1562
rect 20076 1498 20128 1504
rect 20088 1290 20116 1498
rect 20180 1358 20208 2042
rect 20272 1562 20300 2586
rect 21928 2582 21956 2926
rect 21916 2576 21968 2582
rect 21916 2518 21968 2524
rect 20444 1828 20496 1834
rect 20444 1770 20496 1776
rect 20260 1556 20312 1562
rect 20260 1498 20312 1504
rect 20456 1426 20484 1770
rect 20444 1420 20496 1426
rect 20444 1362 20496 1368
rect 21824 1420 21876 1426
rect 21824 1362 21876 1368
rect 20168 1352 20220 1358
rect 20168 1294 20220 1300
rect 20076 1284 20128 1290
rect 20076 1226 20128 1232
rect 20456 1018 20484 1362
rect 21732 1352 21784 1358
rect 21732 1294 21784 1300
rect 21272 1216 21324 1222
rect 21272 1158 21324 1164
rect 19984 1012 20036 1018
rect 19984 954 20036 960
rect 20444 1012 20496 1018
rect 20444 954 20496 960
rect 21284 814 21312 1158
rect 21744 814 21772 1294
rect 21836 1018 21864 1362
rect 21824 1012 21876 1018
rect 21824 954 21876 960
rect 21928 882 21956 2518
rect 22020 2106 22048 3606
rect 22388 2106 22416 3946
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22572 2854 22600 3878
rect 22664 3738 22692 4082
rect 22926 4040 22982 4049
rect 22926 3975 22928 3984
rect 22980 3975 22982 3984
rect 23296 4004 23348 4010
rect 22928 3946 22980 3952
rect 23296 3946 23348 3952
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23216 3738 23244 3878
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 23308 3194 23336 3946
rect 23400 3194 23428 5732
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23492 5030 23520 5646
rect 23584 5370 23612 5850
rect 23952 5778 23980 6072
rect 23940 5772 23992 5778
rect 23940 5714 23992 5720
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 23848 5092 23900 5098
rect 23848 5034 23900 5040
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23512 4924 23820 4933
rect 23512 4922 23518 4924
rect 23574 4922 23598 4924
rect 23654 4922 23678 4924
rect 23734 4922 23758 4924
rect 23814 4922 23820 4924
rect 23574 4870 23576 4922
rect 23756 4870 23758 4922
rect 23512 4868 23518 4870
rect 23574 4868 23598 4870
rect 23654 4868 23678 4870
rect 23734 4868 23758 4870
rect 23814 4868 23820 4870
rect 23512 4859 23820 4868
rect 23512 3836 23820 3845
rect 23512 3834 23518 3836
rect 23574 3834 23598 3836
rect 23654 3834 23678 3836
rect 23734 3834 23758 3836
rect 23814 3834 23820 3836
rect 23574 3782 23576 3834
rect 23756 3782 23758 3834
rect 23512 3780 23518 3782
rect 23574 3780 23598 3782
rect 23654 3780 23678 3782
rect 23734 3780 23758 3782
rect 23814 3780 23820 3782
rect 23512 3771 23820 3780
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 23512 2748 23820 2757
rect 23512 2746 23518 2748
rect 23574 2746 23598 2748
rect 23654 2746 23678 2748
rect 23734 2746 23758 2748
rect 23814 2746 23820 2748
rect 23574 2694 23576 2746
rect 23756 2694 23758 2746
rect 23512 2692 23518 2694
rect 23574 2692 23598 2694
rect 23654 2692 23678 2694
rect 23734 2692 23758 2694
rect 23814 2692 23820 2694
rect 23512 2683 23820 2692
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22008 2100 22060 2106
rect 22008 2042 22060 2048
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 22848 1902 22876 2450
rect 22836 1896 22888 1902
rect 22836 1838 22888 1844
rect 22008 1760 22060 1766
rect 22008 1702 22060 1708
rect 22100 1760 22152 1766
rect 22100 1702 22152 1708
rect 22020 1562 22048 1702
rect 22008 1556 22060 1562
rect 22008 1498 22060 1504
rect 22112 1222 22140 1702
rect 22848 1562 22876 1838
rect 23512 1660 23820 1669
rect 23512 1658 23518 1660
rect 23574 1658 23598 1660
rect 23654 1658 23678 1660
rect 23734 1658 23758 1660
rect 23814 1658 23820 1660
rect 23574 1606 23576 1658
rect 23756 1606 23758 1658
rect 23512 1604 23518 1606
rect 23574 1604 23598 1606
rect 23654 1604 23678 1606
rect 23734 1604 23758 1606
rect 23814 1604 23820 1606
rect 23512 1595 23820 1604
rect 23860 1562 23888 5034
rect 24044 4146 24072 9930
rect 24136 9518 24164 15302
rect 24228 14482 24256 15438
rect 24320 14958 24348 15506
rect 24412 15162 24440 15506
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24308 14816 24360 14822
rect 24360 14764 24440 14770
rect 24308 14758 24440 14764
rect 24320 14742 24440 14758
rect 24216 14476 24268 14482
rect 24216 14418 24268 14424
rect 24228 14090 24256 14418
rect 24228 14062 24348 14090
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 24122 9208 24178 9217
rect 24122 9143 24178 9152
rect 24136 9110 24164 9143
rect 24124 9104 24176 9110
rect 24124 9046 24176 9052
rect 24228 8922 24256 13670
rect 24320 12186 24348 14062
rect 24412 13682 24440 14742
rect 24596 14482 24624 14894
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24412 13654 24532 13682
rect 24400 13388 24452 13394
rect 24400 13330 24452 13336
rect 24412 12782 24440 13330
rect 24400 12776 24452 12782
rect 24400 12718 24452 12724
rect 24412 12442 24440 12718
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24398 12200 24454 12209
rect 24320 12158 24398 12186
rect 24398 12135 24454 12144
rect 24504 12050 24532 13654
rect 24596 13326 24624 14418
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 24688 12434 24716 14214
rect 24136 8894 24256 8922
rect 24320 12022 24532 12050
rect 24596 12406 24716 12434
rect 24136 8838 24164 8894
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 24124 8424 24176 8430
rect 24124 8366 24176 8372
rect 24136 4282 24164 8366
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 24228 6254 24256 6394
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24320 5710 24348 12022
rect 24596 11914 24624 12406
rect 24676 12300 24728 12306
rect 24676 12242 24728 12248
rect 24412 11886 24624 11914
rect 24412 11744 24440 11886
rect 24582 11792 24638 11801
rect 24412 11716 24532 11744
rect 24582 11727 24638 11736
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24412 9926 24440 11290
rect 24504 10130 24532 11716
rect 24596 11626 24624 11727
rect 24584 11620 24636 11626
rect 24584 11562 24636 11568
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24400 9920 24452 9926
rect 24400 9862 24452 9868
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 24504 9081 24532 9454
rect 24596 9450 24624 11562
rect 24688 11082 24716 12242
rect 24780 11762 24808 15846
rect 24964 14550 24992 16390
rect 25424 15978 25452 16594
rect 25412 15972 25464 15978
rect 25412 15914 25464 15920
rect 25964 15564 26016 15570
rect 25964 15506 26016 15512
rect 25976 14958 26004 15506
rect 26240 15360 26292 15366
rect 26240 15302 26292 15308
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24872 14074 24900 14214
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 25976 13870 26004 14894
rect 26252 14890 26280 15302
rect 26240 14884 26292 14890
rect 26240 14826 26292 14832
rect 25964 13864 26016 13870
rect 25964 13806 26016 13812
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 25056 13394 25084 13670
rect 25044 13388 25096 13394
rect 24964 13348 25044 13376
rect 24964 12986 24992 13348
rect 25044 13330 25096 13336
rect 25976 13326 26004 13806
rect 25412 13320 25464 13326
rect 25412 13262 25464 13268
rect 25688 13320 25740 13326
rect 25688 13262 25740 13268
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 25056 12986 25084 13126
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25056 12782 25084 12922
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 25424 12646 25452 13262
rect 25700 12850 25728 13262
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 24872 11642 24900 12378
rect 25332 12345 25360 12582
rect 25318 12336 25374 12345
rect 25318 12271 25374 12280
rect 24780 11614 24900 11642
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 25964 11620 26016 11626
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24688 9518 24716 11018
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24584 9444 24636 9450
rect 24584 9386 24636 9392
rect 24490 9072 24546 9081
rect 24400 9036 24452 9042
rect 24490 9007 24546 9016
rect 24400 8978 24452 8984
rect 24412 8430 24440 8978
rect 24780 8945 24808 11614
rect 25964 11562 26016 11568
rect 24860 11552 24912 11558
rect 24860 11494 24912 11500
rect 24872 9178 24900 11494
rect 25504 11212 25556 11218
rect 25504 11154 25556 11160
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25424 10130 25452 10542
rect 25516 10470 25544 11154
rect 25596 11008 25648 11014
rect 25596 10950 25648 10956
rect 25504 10464 25556 10470
rect 25504 10406 25556 10412
rect 25516 10198 25544 10406
rect 25504 10192 25556 10198
rect 25504 10134 25556 10140
rect 25412 10124 25464 10130
rect 25412 10066 25464 10072
rect 25608 10062 25636 10950
rect 25976 10810 26004 11562
rect 26252 11286 26280 11630
rect 26240 11280 26292 11286
rect 26240 11222 26292 11228
rect 25688 10804 25740 10810
rect 25688 10746 25740 10752
rect 25964 10804 26016 10810
rect 25964 10746 26016 10752
rect 25700 10470 25728 10746
rect 25976 10674 26004 10746
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 25688 10464 25740 10470
rect 25688 10406 25740 10412
rect 25700 10266 25728 10406
rect 25688 10260 25740 10266
rect 25688 10202 25740 10208
rect 25596 10056 25648 10062
rect 25596 9998 25648 10004
rect 25686 9616 25742 9625
rect 25686 9551 25688 9560
rect 25740 9551 25742 9560
rect 25688 9522 25740 9528
rect 26344 9489 26372 16934
rect 26424 16584 26476 16590
rect 26424 16526 26476 16532
rect 26436 15978 26464 16526
rect 26884 16448 26936 16454
rect 26884 16390 26936 16396
rect 26896 16250 26924 16390
rect 26884 16244 26936 16250
rect 26884 16186 26936 16192
rect 27080 16114 27108 17070
rect 27436 17060 27488 17066
rect 27436 17002 27488 17008
rect 27160 16788 27212 16794
rect 27160 16730 27212 16736
rect 27172 16590 27200 16730
rect 27448 16658 27476 17002
rect 30012 16992 30064 16998
rect 30012 16934 30064 16940
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 28724 16652 28776 16658
rect 28724 16594 28776 16600
rect 29184 16652 29236 16658
rect 29184 16594 29236 16600
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 27365 16348 27673 16357
rect 27365 16346 27371 16348
rect 27427 16346 27451 16348
rect 27507 16346 27531 16348
rect 27587 16346 27611 16348
rect 27667 16346 27673 16348
rect 27427 16294 27429 16346
rect 27609 16294 27611 16346
rect 27365 16292 27371 16294
rect 27427 16292 27451 16294
rect 27507 16292 27531 16294
rect 27587 16292 27611 16294
rect 27667 16292 27673 16294
rect 27365 16283 27673 16292
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 26424 15972 26476 15978
rect 26424 15914 26476 15920
rect 27080 15570 27108 16050
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27540 15638 27568 15982
rect 27528 15632 27580 15638
rect 27528 15574 27580 15580
rect 27068 15564 27120 15570
rect 27068 15506 27120 15512
rect 27365 15260 27673 15269
rect 27365 15258 27371 15260
rect 27427 15258 27451 15260
rect 27507 15258 27531 15260
rect 27587 15258 27611 15260
rect 27667 15258 27673 15260
rect 27427 15206 27429 15258
rect 27609 15206 27611 15258
rect 27365 15204 27371 15206
rect 27427 15204 27451 15206
rect 27507 15204 27531 15206
rect 27587 15204 27611 15206
rect 27667 15204 27673 15206
rect 27365 15195 27673 15204
rect 26792 14884 26844 14890
rect 26792 14826 26844 14832
rect 26804 14618 26832 14826
rect 26792 14612 26844 14618
rect 26792 14554 26844 14560
rect 26792 14476 26844 14482
rect 26792 14418 26844 14424
rect 27804 14476 27856 14482
rect 27804 14418 27856 14424
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26620 13938 26648 14350
rect 26804 14074 26832 14418
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27365 14172 27673 14181
rect 27365 14170 27371 14172
rect 27427 14170 27451 14172
rect 27507 14170 27531 14172
rect 27587 14170 27611 14172
rect 27667 14170 27673 14172
rect 27427 14118 27429 14170
rect 27609 14118 27611 14170
rect 27365 14116 27371 14118
rect 27427 14116 27451 14118
rect 27507 14116 27531 14118
rect 27587 14116 27611 14118
rect 27667 14116 27673 14118
rect 27365 14107 27673 14116
rect 27724 14074 27752 14350
rect 26792 14068 26844 14074
rect 26792 14010 26844 14016
rect 27712 14068 27764 14074
rect 27712 14010 27764 14016
rect 27816 13938 27844 14418
rect 28080 14340 28132 14346
rect 28080 14282 28132 14288
rect 28092 14006 28120 14282
rect 28080 14000 28132 14006
rect 28080 13942 28132 13948
rect 26608 13932 26660 13938
rect 26608 13874 26660 13880
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 26516 13864 26568 13870
rect 26516 13806 26568 13812
rect 26528 13394 26556 13806
rect 26620 13734 26648 13874
rect 26792 13796 26844 13802
rect 26792 13738 26844 13744
rect 28080 13796 28132 13802
rect 28080 13738 28132 13744
rect 26608 13728 26660 13734
rect 26608 13670 26660 13676
rect 26620 13530 26648 13670
rect 26804 13530 26832 13738
rect 26608 13524 26660 13530
rect 26608 13466 26660 13472
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 26516 13388 26568 13394
rect 26516 13330 26568 13336
rect 26424 12708 26476 12714
rect 26528 12696 26556 13330
rect 27365 13084 27673 13093
rect 27365 13082 27371 13084
rect 27427 13082 27451 13084
rect 27507 13082 27531 13084
rect 27587 13082 27611 13084
rect 27667 13082 27673 13084
rect 27427 13030 27429 13082
rect 27609 13030 27611 13082
rect 27365 13028 27371 13030
rect 27427 13028 27451 13030
rect 27507 13028 27531 13030
rect 27587 13028 27611 13030
rect 27667 13028 27673 13030
rect 27365 13019 27673 13028
rect 26476 12668 26556 12696
rect 26976 12708 27028 12714
rect 26424 12650 26476 12656
rect 26976 12650 27028 12656
rect 26988 12374 27016 12650
rect 26976 12368 27028 12374
rect 26976 12310 27028 12316
rect 26988 11694 27016 12310
rect 27365 11996 27673 12005
rect 27365 11994 27371 11996
rect 27427 11994 27451 11996
rect 27507 11994 27531 11996
rect 27587 11994 27611 11996
rect 27667 11994 27673 11996
rect 27427 11942 27429 11994
rect 27609 11942 27611 11994
rect 27365 11940 27371 11942
rect 27427 11940 27451 11942
rect 27507 11940 27531 11942
rect 27587 11940 27611 11942
rect 27667 11940 27673 11942
rect 27365 11931 27673 11940
rect 26976 11688 27028 11694
rect 26976 11630 27028 11636
rect 27252 11620 27304 11626
rect 27252 11562 27304 11568
rect 27264 11354 27292 11562
rect 27252 11348 27304 11354
rect 27252 11290 27304 11296
rect 27724 11257 27752 13466
rect 28092 13462 28120 13738
rect 28080 13456 28132 13462
rect 28080 13398 28132 13404
rect 28172 12300 28224 12306
rect 28172 12242 28224 12248
rect 28184 11762 28212 12242
rect 28172 11756 28224 11762
rect 28172 11698 28224 11704
rect 27988 11620 28040 11626
rect 27988 11562 28040 11568
rect 27710 11248 27766 11257
rect 27710 11183 27766 11192
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 27252 11144 27304 11150
rect 27252 11086 27304 11092
rect 26436 10810 26464 11086
rect 26792 11008 26844 11014
rect 26792 10950 26844 10956
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26436 10606 26464 10746
rect 26804 10606 26832 10950
rect 27264 10810 27292 11086
rect 28000 11082 28028 11562
rect 28184 11354 28212 11698
rect 28172 11348 28224 11354
rect 28172 11290 28224 11296
rect 28080 11280 28132 11286
rect 28080 11222 28132 11228
rect 27988 11076 28040 11082
rect 27988 11018 28040 11024
rect 27365 10908 27673 10917
rect 27365 10906 27371 10908
rect 27427 10906 27451 10908
rect 27507 10906 27531 10908
rect 27587 10906 27611 10908
rect 27667 10906 27673 10908
rect 27427 10854 27429 10906
rect 27609 10854 27611 10906
rect 27365 10852 27371 10854
rect 27427 10852 27451 10854
rect 27507 10852 27531 10854
rect 27587 10852 27611 10854
rect 27667 10852 27673 10854
rect 27365 10843 27673 10852
rect 28092 10810 28120 11222
rect 28184 10810 28212 11290
rect 27252 10804 27304 10810
rect 27252 10746 27304 10752
rect 28080 10804 28132 10810
rect 28080 10746 28132 10752
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 27264 10674 27292 10746
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 26424 10600 26476 10606
rect 26424 10542 26476 10548
rect 26792 10600 26844 10606
rect 26792 10542 26844 10548
rect 26330 9480 26386 9489
rect 26804 9450 26832 10542
rect 26884 10260 26936 10266
rect 26884 10202 26936 10208
rect 26896 10169 26924 10202
rect 27988 10192 28040 10198
rect 26882 10160 26938 10169
rect 28092 10180 28120 10746
rect 28040 10152 28120 10180
rect 27988 10134 28040 10140
rect 26882 10095 26938 10104
rect 27365 9820 27673 9829
rect 27365 9818 27371 9820
rect 27427 9818 27451 9820
rect 27507 9818 27531 9820
rect 27587 9818 27611 9820
rect 27667 9818 27673 9820
rect 27427 9766 27429 9818
rect 27609 9766 27611 9818
rect 27365 9764 27371 9766
rect 27427 9764 27451 9766
rect 27507 9764 27531 9766
rect 27587 9764 27611 9766
rect 27667 9764 27673 9766
rect 27365 9755 27673 9764
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 26330 9415 26386 9424
rect 26792 9444 26844 9450
rect 26792 9386 26844 9392
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24766 8936 24822 8945
rect 24766 8871 24822 8880
rect 24872 8809 24900 9114
rect 27908 9042 27936 9454
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 27896 9036 27948 9042
rect 27896 8978 27948 8984
rect 25320 8832 25372 8838
rect 24858 8800 24914 8809
rect 25320 8774 25372 8780
rect 24858 8735 24914 8744
rect 25332 8634 25360 8774
rect 26528 8634 26556 8978
rect 27365 8732 27673 8741
rect 27365 8730 27371 8732
rect 27427 8730 27451 8732
rect 27507 8730 27531 8732
rect 27587 8730 27611 8732
rect 27667 8730 27673 8732
rect 27427 8678 27429 8730
rect 27609 8678 27611 8730
rect 27365 8676 27371 8678
rect 27427 8676 27451 8678
rect 27507 8676 27531 8678
rect 27587 8676 27611 8678
rect 27667 8676 27673 8678
rect 27365 8667 27673 8676
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 27908 8498 27936 8978
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 24400 8424 24452 8430
rect 24400 8366 24452 8372
rect 24412 7206 24440 8366
rect 25780 8356 25832 8362
rect 25780 8298 25832 8304
rect 24492 8288 24544 8294
rect 24492 8230 24544 8236
rect 24504 8090 24532 8230
rect 24492 8084 24544 8090
rect 24492 8026 24544 8032
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 24688 7478 24716 7686
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24400 6928 24452 6934
rect 24400 6870 24452 6876
rect 24308 5704 24360 5710
rect 24308 5646 24360 5652
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 22468 1556 22520 1562
rect 22468 1498 22520 1504
rect 22836 1556 22888 1562
rect 22836 1498 22888 1504
rect 23848 1556 23900 1562
rect 23848 1498 23900 1504
rect 22100 1216 22152 1222
rect 22100 1158 22152 1164
rect 22112 1018 22140 1158
rect 22480 1018 22508 1498
rect 22928 1420 22980 1426
rect 22928 1362 22980 1368
rect 23572 1420 23624 1426
rect 23572 1362 23624 1368
rect 22100 1012 22152 1018
rect 22100 954 22152 960
rect 22468 1012 22520 1018
rect 22468 954 22520 960
rect 21916 876 21968 882
rect 21916 818 21968 824
rect 22940 814 22968 1362
rect 23584 1018 23612 1362
rect 23572 1012 23624 1018
rect 23572 954 23624 960
rect 23848 944 23900 950
rect 23952 932 23980 4014
rect 24412 3738 24440 6870
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 24492 6112 24544 6118
rect 24492 6054 24544 6060
rect 24504 5914 24532 6054
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 25148 5846 25176 6190
rect 25320 5908 25372 5914
rect 25320 5850 25372 5856
rect 25136 5840 25188 5846
rect 25136 5782 25188 5788
rect 25332 5710 25360 5850
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 25320 5704 25372 5710
rect 25320 5646 25372 5652
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24872 5098 24900 5306
rect 24964 5166 24992 5646
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 25056 5370 25084 5510
rect 25044 5364 25096 5370
rect 25044 5306 25096 5312
rect 25424 5234 25452 7822
rect 25792 6254 25820 8298
rect 27908 8090 27936 8434
rect 27896 8084 27948 8090
rect 27896 8026 27948 8032
rect 25964 7948 26016 7954
rect 25964 7890 26016 7896
rect 27804 7948 27856 7954
rect 27804 7890 27856 7896
rect 25976 7342 26004 7890
rect 26698 7848 26754 7857
rect 26698 7783 26700 7792
rect 26752 7783 26754 7792
rect 26700 7754 26752 7760
rect 27365 7644 27673 7653
rect 27365 7642 27371 7644
rect 27427 7642 27451 7644
rect 27507 7642 27531 7644
rect 27587 7642 27611 7644
rect 27667 7642 27673 7644
rect 27427 7590 27429 7642
rect 27609 7590 27611 7642
rect 27365 7588 27371 7590
rect 27427 7588 27451 7590
rect 27507 7588 27531 7590
rect 27587 7588 27611 7590
rect 27667 7588 27673 7590
rect 27365 7579 27673 7588
rect 27816 7546 27844 7890
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 27908 7410 27936 8026
rect 27896 7404 27948 7410
rect 27896 7346 27948 7352
rect 25964 7336 26016 7342
rect 25964 7278 26016 7284
rect 25976 6934 26004 7278
rect 27528 7268 27580 7274
rect 27528 7210 27580 7216
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 25964 6928 26016 6934
rect 25964 6870 26016 6876
rect 26068 6254 26096 7142
rect 27540 7002 27568 7210
rect 27908 7002 27936 7346
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 27712 6996 27764 7002
rect 27712 6938 27764 6944
rect 27896 6996 27948 7002
rect 27896 6938 27948 6944
rect 26240 6860 26292 6866
rect 26240 6802 26292 6808
rect 26252 6390 26280 6802
rect 27160 6656 27212 6662
rect 27160 6598 27212 6604
rect 26240 6384 26292 6390
rect 26240 6326 26292 6332
rect 25780 6248 25832 6254
rect 25780 6190 25832 6196
rect 26056 6248 26108 6254
rect 26056 6190 26108 6196
rect 26068 5846 26096 6190
rect 26252 5846 26280 6326
rect 27172 6254 27200 6598
rect 27365 6556 27673 6565
rect 27365 6554 27371 6556
rect 27427 6554 27451 6556
rect 27507 6554 27531 6556
rect 27587 6554 27611 6556
rect 27667 6554 27673 6556
rect 27427 6502 27429 6554
rect 27609 6502 27611 6554
rect 27365 6500 27371 6502
rect 27427 6500 27451 6502
rect 27507 6500 27531 6502
rect 27587 6500 27611 6502
rect 27667 6500 27673 6502
rect 27365 6491 27673 6500
rect 27724 6338 27752 6938
rect 27804 6860 27856 6866
rect 27804 6802 27856 6808
rect 27632 6310 27752 6338
rect 27632 6254 27660 6310
rect 26332 6248 26384 6254
rect 26332 6190 26384 6196
rect 27160 6248 27212 6254
rect 27160 6190 27212 6196
rect 27436 6248 27488 6254
rect 27436 6190 27488 6196
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 26344 5914 26372 6190
rect 26332 5908 26384 5914
rect 26332 5850 26384 5856
rect 26056 5840 26108 5846
rect 26056 5782 26108 5788
rect 26240 5840 26292 5846
rect 26240 5782 26292 5788
rect 27172 5778 27200 6190
rect 27448 6118 27476 6190
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 27816 5914 27844 6802
rect 28172 6656 28224 6662
rect 28172 6598 28224 6604
rect 28184 6254 28212 6598
rect 28172 6248 28224 6254
rect 28172 6190 28224 6196
rect 27804 5908 27856 5914
rect 27804 5850 27856 5856
rect 27988 5840 28040 5846
rect 27988 5782 28040 5788
rect 27160 5772 27212 5778
rect 27160 5714 27212 5720
rect 25412 5228 25464 5234
rect 25412 5170 25464 5176
rect 24952 5160 25004 5166
rect 24952 5102 25004 5108
rect 24860 5092 24912 5098
rect 24860 5034 24912 5040
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 24780 4282 24808 4626
rect 24768 4276 24820 4282
rect 24768 4218 24820 4224
rect 25424 4154 25452 5170
rect 27172 5166 27200 5714
rect 27365 5468 27673 5477
rect 27365 5466 27371 5468
rect 27427 5466 27451 5468
rect 27507 5466 27531 5468
rect 27587 5466 27611 5468
rect 27667 5466 27673 5468
rect 27427 5414 27429 5466
rect 27609 5414 27611 5466
rect 27365 5412 27371 5414
rect 27427 5412 27451 5414
rect 27507 5412 27531 5414
rect 27587 5412 27611 5414
rect 27667 5412 27673 5414
rect 27365 5403 27673 5412
rect 28000 5166 28028 5782
rect 27160 5160 27212 5166
rect 27160 5102 27212 5108
rect 27988 5160 28040 5166
rect 27988 5102 28040 5108
rect 27712 4684 27764 4690
rect 27712 4626 27764 4632
rect 27365 4380 27673 4389
rect 27365 4378 27371 4380
rect 27427 4378 27451 4380
rect 27507 4378 27531 4380
rect 27587 4378 27611 4380
rect 27667 4378 27673 4380
rect 27427 4326 27429 4378
rect 27609 4326 27611 4378
rect 27365 4324 27371 4326
rect 27427 4324 27451 4326
rect 27507 4324 27531 4326
rect 27587 4324 27611 4326
rect 27667 4324 27673 4326
rect 27365 4315 27673 4324
rect 25240 4126 25452 4154
rect 24584 4004 24636 4010
rect 24584 3946 24636 3952
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24504 3670 24532 3878
rect 24596 3738 24624 3946
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24492 3664 24544 3670
rect 24492 3606 24544 3612
rect 25240 3398 25268 4126
rect 26056 4072 26108 4078
rect 26056 4014 26108 4020
rect 26606 4040 26662 4049
rect 25596 3664 25648 3670
rect 25596 3606 25648 3612
rect 25412 3596 25464 3602
rect 25412 3538 25464 3544
rect 25228 3392 25280 3398
rect 25148 3340 25228 3346
rect 25148 3334 25280 3340
rect 25148 3318 25268 3334
rect 25148 2990 25176 3318
rect 25424 3126 25452 3538
rect 25412 3120 25464 3126
rect 25412 3062 25464 3068
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 24032 2916 24084 2922
rect 24032 2858 24084 2864
rect 24952 2916 25004 2922
rect 24952 2858 25004 2864
rect 24044 2650 24072 2858
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24136 2106 24164 2450
rect 24964 2310 24992 2858
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24952 2304 25004 2310
rect 24952 2246 25004 2252
rect 24504 2106 24532 2246
rect 24124 2100 24176 2106
rect 24124 2042 24176 2048
rect 24492 2100 24544 2106
rect 24492 2042 24544 2048
rect 25148 1970 25176 2926
rect 25608 2854 25636 3606
rect 26068 3534 26096 4014
rect 26332 4004 26384 4010
rect 26606 3975 26662 3984
rect 27252 4004 27304 4010
rect 26332 3946 26384 3952
rect 26056 3528 26108 3534
rect 26056 3470 26108 3476
rect 26344 2990 26372 3946
rect 26620 3942 26648 3975
rect 27252 3946 27304 3952
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 27264 3738 27292 3946
rect 27724 3924 27752 4626
rect 28000 4622 28028 5102
rect 28276 4758 28304 16390
rect 28736 16250 28764 16594
rect 29196 16250 29224 16594
rect 30024 16590 30052 16934
rect 31217 16892 31525 16901
rect 31217 16890 31223 16892
rect 31279 16890 31303 16892
rect 31359 16890 31383 16892
rect 31439 16890 31463 16892
rect 31519 16890 31525 16892
rect 31279 16838 31281 16890
rect 31461 16838 31463 16890
rect 31217 16836 31223 16838
rect 31279 16836 31303 16838
rect 31359 16836 31383 16838
rect 31439 16836 31463 16838
rect 31519 16836 31525 16838
rect 31217 16827 31525 16836
rect 30012 16584 30064 16590
rect 30012 16526 30064 16532
rect 28724 16244 28776 16250
rect 28724 16186 28776 16192
rect 29184 16244 29236 16250
rect 29184 16186 29236 16192
rect 29000 15972 29052 15978
rect 29000 15914 29052 15920
rect 28448 15904 28500 15910
rect 28448 15846 28500 15852
rect 28632 15904 28684 15910
rect 28632 15846 28684 15852
rect 28460 15706 28488 15846
rect 28448 15700 28500 15706
rect 28448 15642 28500 15648
rect 28644 15570 28672 15846
rect 29012 15706 29040 15914
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 28632 15564 28684 15570
rect 28632 15506 28684 15512
rect 28644 15450 28672 15506
rect 28644 15422 28764 15450
rect 29196 15434 29224 16186
rect 29276 15904 29328 15910
rect 29276 15846 29328 15852
rect 28736 15162 28764 15422
rect 28816 15428 28868 15434
rect 28816 15370 28868 15376
rect 29184 15428 29236 15434
rect 29184 15370 29236 15376
rect 28724 15156 28776 15162
rect 28724 15098 28776 15104
rect 28724 15020 28776 15026
rect 28828 15008 28856 15370
rect 29288 15162 29316 15846
rect 30024 15706 30052 16526
rect 31217 15804 31525 15813
rect 31217 15802 31223 15804
rect 31279 15802 31303 15804
rect 31359 15802 31383 15804
rect 31439 15802 31463 15804
rect 31519 15802 31525 15804
rect 31279 15750 31281 15802
rect 31461 15750 31463 15802
rect 31217 15748 31223 15750
rect 31279 15748 31303 15750
rect 31359 15748 31383 15750
rect 31439 15748 31463 15750
rect 31519 15748 31525 15750
rect 31217 15739 31525 15748
rect 30012 15700 30064 15706
rect 30012 15642 30064 15648
rect 29552 15564 29604 15570
rect 29552 15506 29604 15512
rect 29276 15156 29328 15162
rect 29276 15098 29328 15104
rect 28776 14980 28856 15008
rect 28724 14962 28776 14968
rect 29184 14952 29236 14958
rect 29184 14894 29236 14900
rect 29460 14952 29512 14958
rect 29460 14894 29512 14900
rect 29196 14618 29224 14894
rect 29368 14816 29420 14822
rect 29368 14758 29420 14764
rect 29184 14612 29236 14618
rect 29184 14554 29236 14560
rect 28908 14544 28960 14550
rect 28908 14486 28960 14492
rect 28920 14385 28948 14486
rect 28906 14376 28962 14385
rect 28906 14311 28962 14320
rect 29196 13938 29224 14554
rect 29276 14340 29328 14346
rect 29276 14282 29328 14288
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 29288 13870 29316 14282
rect 29380 14074 29408 14758
rect 29472 14278 29500 14894
rect 29564 14550 29592 15506
rect 30932 15360 30984 15366
rect 30932 15302 30984 15308
rect 29644 15088 29696 15094
rect 29644 15030 29696 15036
rect 29656 14822 29684 15030
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 29656 14550 29684 14758
rect 29552 14544 29604 14550
rect 29552 14486 29604 14492
rect 29644 14544 29696 14550
rect 29644 14486 29696 14492
rect 29460 14272 29512 14278
rect 29460 14214 29512 14220
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 29288 13462 29316 13806
rect 29472 13734 29500 14214
rect 30944 14074 30972 15302
rect 31217 14716 31525 14725
rect 31217 14714 31223 14716
rect 31279 14714 31303 14716
rect 31359 14714 31383 14716
rect 31439 14714 31463 14716
rect 31519 14714 31525 14716
rect 31279 14662 31281 14714
rect 31461 14662 31463 14714
rect 31217 14660 31223 14662
rect 31279 14660 31303 14662
rect 31359 14660 31383 14662
rect 31439 14660 31463 14662
rect 31519 14660 31525 14662
rect 31217 14651 31525 14660
rect 30932 14068 30984 14074
rect 30932 14010 30984 14016
rect 29460 13728 29512 13734
rect 29460 13670 29512 13676
rect 29276 13456 29328 13462
rect 29276 13398 29328 13404
rect 29092 13184 29144 13190
rect 29092 13126 29144 13132
rect 29104 12782 29132 13126
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 29000 12776 29052 12782
rect 29000 12718 29052 12724
rect 29092 12776 29144 12782
rect 29092 12718 29144 12724
rect 28632 12436 28684 12442
rect 28632 12378 28684 12384
rect 28644 12345 28672 12378
rect 28630 12336 28686 12345
rect 28630 12271 28686 12280
rect 29012 11898 29040 12718
rect 29104 12374 29132 12718
rect 29092 12368 29144 12374
rect 29092 12310 29144 12316
rect 29196 11898 29224 12786
rect 29472 12782 29500 13670
rect 31217 13628 31525 13637
rect 31217 13626 31223 13628
rect 31279 13626 31303 13628
rect 31359 13626 31383 13628
rect 31439 13626 31463 13628
rect 31519 13626 31525 13628
rect 31279 13574 31281 13626
rect 31461 13574 31463 13626
rect 31217 13572 31223 13574
rect 31279 13572 31303 13574
rect 31359 13572 31383 13574
rect 31439 13572 31463 13574
rect 31519 13572 31525 13574
rect 31217 13563 31525 13572
rect 30746 13424 30802 13433
rect 30746 13359 30802 13368
rect 30760 12986 30788 13359
rect 30748 12980 30800 12986
rect 30748 12922 30800 12928
rect 29460 12776 29512 12782
rect 29460 12718 29512 12724
rect 29276 12640 29328 12646
rect 29276 12582 29328 12588
rect 29920 12640 29972 12646
rect 29920 12582 29972 12588
rect 29288 12306 29316 12582
rect 29932 12306 29960 12582
rect 31217 12540 31525 12549
rect 31217 12538 31223 12540
rect 31279 12538 31303 12540
rect 31359 12538 31383 12540
rect 31439 12538 31463 12540
rect 31519 12538 31525 12540
rect 31279 12486 31281 12538
rect 31461 12486 31463 12538
rect 31217 12484 31223 12486
rect 31279 12484 31303 12486
rect 31359 12484 31383 12486
rect 31439 12484 31463 12486
rect 31519 12484 31525 12486
rect 31217 12475 31525 12484
rect 29276 12300 29328 12306
rect 29276 12242 29328 12248
rect 29828 12300 29880 12306
rect 29828 12242 29880 12248
rect 29920 12300 29972 12306
rect 29920 12242 29972 12248
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 29184 11892 29236 11898
rect 29184 11834 29236 11840
rect 29288 11762 29316 12242
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 28448 11552 28500 11558
rect 28448 11494 28500 11500
rect 29000 11552 29052 11558
rect 29000 11494 29052 11500
rect 28460 11354 28488 11494
rect 28448 11348 28500 11354
rect 28448 11290 28500 11296
rect 28448 11008 28500 11014
rect 28448 10950 28500 10956
rect 28460 10606 28488 10950
rect 28816 10804 28868 10810
rect 28816 10746 28868 10752
rect 28448 10600 28500 10606
rect 28448 10542 28500 10548
rect 28828 10130 28856 10746
rect 29012 10538 29040 11494
rect 29288 11354 29316 11698
rect 29840 11694 29868 12242
rect 30380 12096 30432 12102
rect 30380 12038 30432 12044
rect 29828 11688 29880 11694
rect 29828 11630 29880 11636
rect 30288 11688 30340 11694
rect 30288 11630 30340 11636
rect 29276 11348 29328 11354
rect 29276 11290 29328 11296
rect 29288 11054 29316 11290
rect 30300 11218 30328 11630
rect 30392 11626 30420 12038
rect 30380 11620 30432 11626
rect 30380 11562 30432 11568
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 29104 11026 29316 11054
rect 29104 10606 29132 11026
rect 29460 10804 29512 10810
rect 29460 10746 29512 10752
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29276 10600 29328 10606
rect 29276 10542 29328 10548
rect 29000 10532 29052 10538
rect 29000 10474 29052 10480
rect 29288 10266 29316 10542
rect 29276 10260 29328 10266
rect 29276 10202 29328 10208
rect 28908 10192 28960 10198
rect 28908 10134 28960 10140
rect 28816 10124 28868 10130
rect 28816 10066 28868 10072
rect 28920 9722 28948 10134
rect 29368 10056 29420 10062
rect 29368 9998 29420 10004
rect 29184 9920 29236 9926
rect 29184 9862 29236 9868
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 29092 9648 29144 9654
rect 29092 9590 29144 9596
rect 29104 9042 29132 9590
rect 29196 9382 29224 9862
rect 29184 9376 29236 9382
rect 29184 9318 29236 9324
rect 29196 9042 29224 9318
rect 29380 9178 29408 9998
rect 29472 9518 29500 10746
rect 30392 10674 30420 11562
rect 31217 11452 31525 11461
rect 31217 11450 31223 11452
rect 31279 11450 31303 11452
rect 31359 11450 31383 11452
rect 31439 11450 31463 11452
rect 31519 11450 31525 11452
rect 31279 11398 31281 11450
rect 31461 11398 31463 11450
rect 31217 11396 31223 11398
rect 31279 11396 31303 11398
rect 31359 11396 31383 11398
rect 31439 11396 31463 11398
rect 31519 11396 31525 11398
rect 31217 11387 31525 11396
rect 30656 11212 30708 11218
rect 30656 11154 30708 11160
rect 30668 10810 30696 11154
rect 30656 10804 30708 10810
rect 30656 10746 30708 10752
rect 30380 10668 30432 10674
rect 30380 10610 30432 10616
rect 29920 10532 29972 10538
rect 29920 10474 29972 10480
rect 29932 10130 29960 10474
rect 30392 10266 30420 10610
rect 31668 10600 31720 10606
rect 31668 10542 31720 10548
rect 31217 10364 31525 10373
rect 31217 10362 31223 10364
rect 31279 10362 31303 10364
rect 31359 10362 31383 10364
rect 31439 10362 31463 10364
rect 31519 10362 31525 10364
rect 31279 10310 31281 10362
rect 31461 10310 31463 10362
rect 31217 10308 31223 10310
rect 31279 10308 31303 10310
rect 31359 10308 31383 10310
rect 31439 10308 31463 10310
rect 31519 10308 31525 10310
rect 31217 10299 31525 10308
rect 31680 10305 31708 10542
rect 31666 10296 31722 10305
rect 30380 10260 30432 10266
rect 31666 10231 31722 10240
rect 30380 10202 30432 10208
rect 30288 10192 30340 10198
rect 30288 10134 30340 10140
rect 29920 10124 29972 10130
rect 29920 10066 29972 10072
rect 30300 9722 30328 10134
rect 30288 9716 30340 9722
rect 30288 9658 30340 9664
rect 30300 9602 30328 9658
rect 30024 9574 30328 9602
rect 29460 9512 29512 9518
rect 29460 9454 29512 9460
rect 29368 9172 29420 9178
rect 29368 9114 29420 9120
rect 28724 9036 28776 9042
rect 29092 9036 29144 9042
rect 28776 8996 29092 9024
rect 28724 8978 28776 8984
rect 29092 8978 29144 8984
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 28448 8832 28500 8838
rect 28448 8774 28500 8780
rect 28724 8832 28776 8838
rect 28724 8774 28776 8780
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 28460 8634 28488 8774
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 28736 8498 28764 8774
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 29196 8430 29224 8774
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 28540 8356 28592 8362
rect 28540 8298 28592 8304
rect 29000 8356 29052 8362
rect 29000 8298 29052 8304
rect 28552 8090 28580 8298
rect 28540 8084 28592 8090
rect 28540 8026 28592 8032
rect 29012 7954 29040 8298
rect 29380 7954 29408 9114
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 29748 8430 29776 8570
rect 30024 8566 30052 9574
rect 30288 9512 30340 9518
rect 30392 9500 30420 10202
rect 30340 9472 30420 9500
rect 30288 9454 30340 9460
rect 31217 9276 31525 9285
rect 31217 9274 31223 9276
rect 31279 9274 31303 9276
rect 31359 9274 31383 9276
rect 31439 9274 31463 9276
rect 31519 9274 31525 9276
rect 31279 9222 31281 9274
rect 31461 9222 31463 9274
rect 31217 9220 31223 9222
rect 31279 9220 31303 9222
rect 31359 9220 31383 9222
rect 31439 9220 31463 9222
rect 31519 9220 31525 9222
rect 30930 9208 30986 9217
rect 31217 9211 31525 9220
rect 30930 9143 30932 9152
rect 30984 9143 30986 9152
rect 30932 9114 30984 9120
rect 30012 8560 30064 8566
rect 30012 8502 30064 8508
rect 29736 8424 29788 8430
rect 29736 8366 29788 8372
rect 30472 8424 30524 8430
rect 30472 8366 30524 8372
rect 29736 8288 29788 8294
rect 29736 8230 29788 8236
rect 30196 8288 30248 8294
rect 30196 8230 30248 8236
rect 30380 8288 30432 8294
rect 30380 8230 30432 8236
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 29368 7948 29420 7954
rect 29368 7890 29420 7896
rect 28448 7812 28500 7818
rect 28448 7754 28500 7760
rect 28460 7342 28488 7754
rect 28632 7744 28684 7750
rect 28632 7686 28684 7692
rect 29184 7744 29236 7750
rect 29184 7686 29236 7692
rect 28448 7336 28500 7342
rect 28448 7278 28500 7284
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28552 6322 28580 7142
rect 28644 6934 28672 7686
rect 28908 7404 28960 7410
rect 28908 7346 28960 7352
rect 28632 6928 28684 6934
rect 28632 6870 28684 6876
rect 28644 6458 28672 6870
rect 28920 6866 28948 7346
rect 29196 7002 29224 7686
rect 29748 7342 29776 8230
rect 30208 8022 30236 8230
rect 30288 8084 30340 8090
rect 30288 8026 30340 8032
rect 30196 8016 30248 8022
rect 30196 7958 30248 7964
rect 30300 7546 30328 8026
rect 30288 7540 30340 7546
rect 30288 7482 30340 7488
rect 29736 7336 29788 7342
rect 29736 7278 29788 7284
rect 29276 7200 29328 7206
rect 29276 7142 29328 7148
rect 29184 6996 29236 7002
rect 29184 6938 29236 6944
rect 28724 6860 28776 6866
rect 28724 6802 28776 6808
rect 28908 6860 28960 6866
rect 28908 6802 28960 6808
rect 28632 6452 28684 6458
rect 28632 6394 28684 6400
rect 28540 6316 28592 6322
rect 28540 6258 28592 6264
rect 28448 6248 28500 6254
rect 28448 6190 28500 6196
rect 28460 5914 28488 6190
rect 28448 5908 28500 5914
rect 28448 5850 28500 5856
rect 28552 5778 28580 6258
rect 28540 5772 28592 5778
rect 28540 5714 28592 5720
rect 28644 5166 28672 6394
rect 28736 5370 28764 6802
rect 28816 6656 28868 6662
rect 28816 6598 28868 6604
rect 28828 6390 28856 6598
rect 28816 6384 28868 6390
rect 28816 6326 28868 6332
rect 28724 5364 28776 5370
rect 28724 5306 28776 5312
rect 28632 5160 28684 5166
rect 28632 5102 28684 5108
rect 28736 4758 28764 5306
rect 28920 5302 28948 6802
rect 29184 6316 29236 6322
rect 29184 6258 29236 6264
rect 29196 5914 29224 6258
rect 29184 5908 29236 5914
rect 29184 5850 29236 5856
rect 29196 5778 29224 5850
rect 29092 5772 29144 5778
rect 29092 5714 29144 5720
rect 29184 5772 29236 5778
rect 29184 5714 29236 5720
rect 28908 5296 28960 5302
rect 28908 5238 28960 5244
rect 28920 5166 28948 5238
rect 28908 5160 28960 5166
rect 28908 5102 28960 5108
rect 29104 4758 29132 5714
rect 29288 5166 29316 7142
rect 29748 6866 29776 7278
rect 29828 7200 29880 7206
rect 29828 7142 29880 7148
rect 29840 6866 29868 7142
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 29828 6860 29880 6866
rect 29828 6802 29880 6808
rect 29736 6656 29788 6662
rect 29736 6598 29788 6604
rect 29748 6254 29776 6598
rect 30392 6254 30420 8230
rect 30484 7342 30512 8366
rect 30748 8288 30800 8294
rect 30748 8230 30800 8236
rect 30564 8016 30616 8022
rect 30564 7958 30616 7964
rect 30576 7342 30604 7958
rect 30760 7818 30788 8230
rect 31217 8188 31525 8197
rect 31217 8186 31223 8188
rect 31279 8186 31303 8188
rect 31359 8186 31383 8188
rect 31439 8186 31463 8188
rect 31519 8186 31525 8188
rect 31279 8134 31281 8186
rect 31461 8134 31463 8186
rect 31217 8132 31223 8134
rect 31279 8132 31303 8134
rect 31359 8132 31383 8134
rect 31439 8132 31463 8134
rect 31519 8132 31525 8134
rect 31217 8123 31525 8132
rect 30932 8084 30984 8090
rect 30932 8026 30984 8032
rect 30944 7993 30972 8026
rect 30930 7984 30986 7993
rect 30930 7919 30986 7928
rect 30748 7812 30800 7818
rect 30748 7754 30800 7760
rect 30760 7546 30788 7754
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 30472 7336 30524 7342
rect 30472 7278 30524 7284
rect 30564 7336 30616 7342
rect 30564 7278 30616 7284
rect 30484 7188 30512 7278
rect 30748 7268 30800 7274
rect 30748 7210 30800 7216
rect 30656 7200 30708 7206
rect 30484 7160 30604 7188
rect 30576 7002 30604 7160
rect 30656 7142 30708 7148
rect 30668 7002 30696 7142
rect 30564 6996 30616 7002
rect 30564 6938 30616 6944
rect 30656 6996 30708 7002
rect 30656 6938 30708 6944
rect 30576 6882 30604 6938
rect 30760 6882 30788 7210
rect 31217 7100 31525 7109
rect 31217 7098 31223 7100
rect 31279 7098 31303 7100
rect 31359 7098 31383 7100
rect 31439 7098 31463 7100
rect 31519 7098 31525 7100
rect 31279 7046 31281 7098
rect 31461 7046 31463 7098
rect 31217 7044 31223 7046
rect 31279 7044 31303 7046
rect 31359 7044 31383 7046
rect 31439 7044 31463 7046
rect 31519 7044 31525 7046
rect 31217 7035 31525 7044
rect 30576 6854 30788 6882
rect 31022 6896 31078 6905
rect 31022 6831 31078 6840
rect 30656 6656 30708 6662
rect 30656 6598 30708 6604
rect 30932 6656 30984 6662
rect 30932 6598 30984 6604
rect 29644 6248 29696 6254
rect 29644 6190 29696 6196
rect 29736 6248 29788 6254
rect 29736 6190 29788 6196
rect 30380 6248 30432 6254
rect 30380 6190 30432 6196
rect 29368 6112 29420 6118
rect 29368 6054 29420 6060
rect 29380 5778 29408 6054
rect 29656 5846 29684 6190
rect 29644 5840 29696 5846
rect 29644 5782 29696 5788
rect 29368 5772 29420 5778
rect 29368 5714 29420 5720
rect 29366 5672 29422 5681
rect 29366 5607 29368 5616
rect 29420 5607 29422 5616
rect 29368 5578 29420 5584
rect 30392 5302 30420 6190
rect 30564 5908 30616 5914
rect 30564 5850 30616 5856
rect 30576 5370 30604 5850
rect 30668 5778 30696 6598
rect 30944 5914 30972 6598
rect 31036 6458 31064 6831
rect 31024 6452 31076 6458
rect 31024 6394 31076 6400
rect 31217 6012 31525 6021
rect 31217 6010 31223 6012
rect 31279 6010 31303 6012
rect 31359 6010 31383 6012
rect 31439 6010 31463 6012
rect 31519 6010 31525 6012
rect 31279 5958 31281 6010
rect 31461 5958 31463 6010
rect 31217 5956 31223 5958
rect 31279 5956 31303 5958
rect 31359 5956 31383 5958
rect 31439 5956 31463 5958
rect 31519 5956 31525 5958
rect 31217 5947 31525 5956
rect 30932 5908 30984 5914
rect 30932 5850 30984 5856
rect 30656 5772 30708 5778
rect 30656 5714 30708 5720
rect 30748 5772 30800 5778
rect 30748 5714 30800 5720
rect 30564 5364 30616 5370
rect 30564 5306 30616 5312
rect 30380 5296 30432 5302
rect 30380 5238 30432 5244
rect 29276 5160 29328 5166
rect 29276 5102 29328 5108
rect 28264 4752 28316 4758
rect 28264 4694 28316 4700
rect 28724 4752 28776 4758
rect 28724 4694 28776 4700
rect 29092 4752 29144 4758
rect 29092 4694 29144 4700
rect 30760 4690 30788 5714
rect 31217 4924 31525 4933
rect 31217 4922 31223 4924
rect 31279 4922 31303 4924
rect 31359 4922 31383 4924
rect 31439 4922 31463 4924
rect 31519 4922 31525 4924
rect 31279 4870 31281 4922
rect 31461 4870 31463 4922
rect 31217 4868 31223 4870
rect 31279 4868 31303 4870
rect 31359 4868 31383 4870
rect 31439 4868 31463 4870
rect 31519 4868 31525 4870
rect 31217 4859 31525 4868
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 30564 4684 30616 4690
rect 30564 4626 30616 4632
rect 30748 4684 30800 4690
rect 30748 4626 30800 4632
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 28000 4078 28028 4558
rect 27988 4072 28040 4078
rect 27988 4014 28040 4020
rect 27804 3936 27856 3942
rect 27724 3896 27804 3924
rect 27724 3738 27752 3896
rect 27804 3878 27856 3884
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 27712 3732 27764 3738
rect 27712 3674 27764 3680
rect 28000 3602 28028 4014
rect 28264 4004 28316 4010
rect 28264 3946 28316 3952
rect 28276 3738 28304 3946
rect 28920 3738 28948 4626
rect 29828 4616 29880 4622
rect 29828 4558 29880 4564
rect 29840 4282 29868 4558
rect 29828 4276 29880 4282
rect 29828 4218 29880 4224
rect 29644 4072 29696 4078
rect 29644 4014 29696 4020
rect 29656 3942 29684 4014
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 29656 3738 29684 3878
rect 28264 3732 28316 3738
rect 28264 3674 28316 3680
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 29644 3732 29696 3738
rect 29644 3674 29696 3680
rect 27160 3596 27212 3602
rect 27160 3538 27212 3544
rect 27252 3596 27304 3602
rect 27252 3538 27304 3544
rect 27988 3596 28040 3602
rect 27988 3538 28040 3544
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 25688 2984 25740 2990
rect 25688 2926 25740 2932
rect 26332 2984 26384 2990
rect 26332 2926 26384 2932
rect 25320 2848 25372 2854
rect 25320 2790 25372 2796
rect 25596 2848 25648 2854
rect 25596 2790 25648 2796
rect 25332 2514 25360 2790
rect 25608 2650 25636 2790
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 25596 2508 25648 2514
rect 25596 2450 25648 2456
rect 25608 2310 25636 2450
rect 25700 2446 25728 2926
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 26160 2582 26188 2790
rect 26148 2576 26200 2582
rect 26148 2518 26200 2524
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 26344 2378 26372 2926
rect 26700 2916 26752 2922
rect 26700 2858 26752 2864
rect 26608 2848 26660 2854
rect 26608 2790 26660 2796
rect 26620 2650 26648 2790
rect 26712 2650 26740 2858
rect 27172 2650 27200 3538
rect 27264 3126 27292 3538
rect 27365 3292 27673 3301
rect 27365 3290 27371 3292
rect 27427 3290 27451 3292
rect 27507 3290 27531 3292
rect 27587 3290 27611 3292
rect 27667 3290 27673 3292
rect 27427 3238 27429 3290
rect 27609 3238 27611 3290
rect 27365 3236 27371 3238
rect 27427 3236 27451 3238
rect 27507 3236 27531 3238
rect 27587 3236 27611 3238
rect 27667 3236 27673 3238
rect 27365 3227 27673 3236
rect 27252 3120 27304 3126
rect 27252 3062 27304 3068
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 27264 2514 27292 3062
rect 28000 2990 28028 3538
rect 29104 3194 29132 3538
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 29840 2990 29868 4218
rect 30576 4146 30604 4626
rect 30564 4140 30616 4146
rect 30564 4082 30616 4088
rect 29920 3936 29972 3942
rect 29920 3878 29972 3884
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 29932 3670 29960 3878
rect 29920 3664 29972 3670
rect 29920 3606 29972 3612
rect 30484 3194 30512 3878
rect 31217 3836 31525 3845
rect 31217 3834 31223 3836
rect 31279 3834 31303 3836
rect 31359 3834 31383 3836
rect 31439 3834 31463 3836
rect 31519 3834 31525 3836
rect 31279 3782 31281 3834
rect 31461 3782 31463 3834
rect 31217 3780 31223 3782
rect 31279 3780 31303 3782
rect 31359 3780 31383 3782
rect 31439 3780 31463 3782
rect 31519 3780 31525 3782
rect 31217 3771 31525 3780
rect 30932 3392 30984 3398
rect 30932 3334 30984 3340
rect 30944 3194 30972 3334
rect 30472 3188 30524 3194
rect 30472 3130 30524 3136
rect 30932 3188 30984 3194
rect 30932 3130 30984 3136
rect 27988 2984 28040 2990
rect 27988 2926 28040 2932
rect 29828 2984 29880 2990
rect 29828 2926 29880 2932
rect 31576 2984 31628 2990
rect 31628 2944 31708 2972
rect 31576 2926 31628 2932
rect 27528 2916 27580 2922
rect 27528 2858 27580 2864
rect 27540 2650 27568 2858
rect 31680 2825 31708 2944
rect 31666 2816 31722 2825
rect 31217 2748 31525 2757
rect 31666 2751 31722 2760
rect 31217 2746 31223 2748
rect 31279 2746 31303 2748
rect 31359 2746 31383 2748
rect 31439 2746 31463 2748
rect 31519 2746 31525 2748
rect 31279 2694 31281 2746
rect 31461 2694 31463 2746
rect 31217 2692 31223 2694
rect 31279 2692 31303 2694
rect 31359 2692 31383 2694
rect 31439 2692 31463 2694
rect 31519 2692 31525 2694
rect 31217 2683 31525 2692
rect 27528 2644 27580 2650
rect 27528 2586 27580 2592
rect 27252 2508 27304 2514
rect 27252 2450 27304 2456
rect 26332 2372 26384 2378
rect 26332 2314 26384 2320
rect 25412 2304 25464 2310
rect 25412 2246 25464 2252
rect 25596 2304 25648 2310
rect 25596 2246 25648 2252
rect 31024 2304 31076 2310
rect 31024 2246 31076 2252
rect 24492 1964 24544 1970
rect 24492 1906 24544 1912
rect 25136 1964 25188 1970
rect 25136 1906 25188 1912
rect 24216 1760 24268 1766
rect 24216 1702 24268 1708
rect 24228 1494 24256 1702
rect 24216 1488 24268 1494
rect 24216 1430 24268 1436
rect 24228 1018 24256 1430
rect 24504 1018 24532 1906
rect 25148 1426 25176 1906
rect 25424 1562 25452 2246
rect 27365 2204 27673 2213
rect 27365 2202 27371 2204
rect 27427 2202 27451 2204
rect 27507 2202 27531 2204
rect 27587 2202 27611 2204
rect 27667 2202 27673 2204
rect 27427 2150 27429 2202
rect 27609 2150 27611 2202
rect 27365 2148 27371 2150
rect 27427 2148 27451 2150
rect 27507 2148 27531 2150
rect 27587 2148 27611 2150
rect 27667 2148 27673 2150
rect 27365 2139 27673 2148
rect 31036 2145 31064 2246
rect 31022 2136 31078 2145
rect 31022 2071 31078 2080
rect 31024 1896 31076 1902
rect 31024 1838 31076 1844
rect 25412 1556 25464 1562
rect 25412 1498 25464 1504
rect 31036 1465 31064 1838
rect 31217 1660 31525 1669
rect 31217 1658 31223 1660
rect 31279 1658 31303 1660
rect 31359 1658 31383 1660
rect 31439 1658 31463 1660
rect 31519 1658 31525 1660
rect 31279 1606 31281 1658
rect 31461 1606 31463 1658
rect 31217 1604 31223 1606
rect 31279 1604 31303 1606
rect 31359 1604 31383 1606
rect 31439 1604 31463 1606
rect 31519 1604 31525 1606
rect 31217 1595 31525 1604
rect 31022 1456 31078 1465
rect 24584 1420 24636 1426
rect 24584 1362 24636 1368
rect 25136 1420 25188 1426
rect 31022 1391 31078 1400
rect 25136 1362 25188 1368
rect 24216 1012 24268 1018
rect 24216 954 24268 960
rect 24492 1012 24544 1018
rect 24492 954 24544 960
rect 23900 904 23980 932
rect 23848 886 23900 892
rect 24596 814 24624 1362
rect 27365 1116 27673 1125
rect 27365 1114 27371 1116
rect 27427 1114 27451 1116
rect 27507 1114 27531 1116
rect 27587 1114 27611 1116
rect 27667 1114 27673 1116
rect 27427 1062 27429 1114
rect 27609 1062 27611 1114
rect 27365 1060 27371 1062
rect 27427 1060 27451 1062
rect 27507 1060 27531 1062
rect 27587 1060 27611 1062
rect 27667 1060 27673 1062
rect 27365 1051 27673 1060
rect 19524 808 19576 814
rect 19524 750 19576 756
rect 21272 808 21324 814
rect 21272 750 21324 756
rect 21732 808 21784 814
rect 21732 750 21784 756
rect 22928 808 22980 814
rect 22928 750 22980 756
rect 24584 808 24636 814
rect 31024 808 31076 814
rect 24584 750 24636 756
rect 31022 776 31024 785
rect 31076 776 31078 785
rect 31022 711 31078 720
rect 23512 572 23820 581
rect 23512 570 23518 572
rect 23574 570 23598 572
rect 23654 570 23678 572
rect 23734 570 23758 572
rect 23814 570 23820 572
rect 23574 518 23576 570
rect 23756 518 23758 570
rect 23512 516 23518 518
rect 23574 516 23598 518
rect 23654 516 23678 518
rect 23734 516 23758 518
rect 23814 516 23820 518
rect 23512 507 23820 516
rect 31217 572 31525 581
rect 31217 570 31223 572
rect 31279 570 31303 572
rect 31359 570 31383 572
rect 31439 570 31463 572
rect 31519 570 31525 572
rect 31279 518 31281 570
rect 31461 518 31463 570
rect 31217 516 31223 518
rect 31279 516 31303 518
rect 31359 516 31383 518
rect 31439 516 31463 518
rect 31519 516 31525 518
rect 31217 507 31525 516
rect 18 0 74 400
rect 662 0 718 400
rect 1306 0 1362 400
rect 1950 0 2006 400
rect 2594 0 2650 400
rect 3238 0 3294 400
rect 3882 0 3938 400
rect 4526 0 4582 400
rect 5170 0 5226 400
rect 5814 0 5870 400
rect 6458 0 6514 400
rect 7102 0 7158 400
rect 7746 0 7802 400
rect 15474 0 15530 400
rect 16118 348 16120 400
rect 16172 348 16174 400
rect 16118 0 16174 348
rect 16304 342 16356 348
rect 16762 0 16818 400
rect 17406 0 17462 400
rect 18050 0 18106 400
<< via2 >>
rect 1122 19760 1178 19816
rect 754 19080 810 19136
rect 8108 19066 8164 19068
rect 8188 19066 8244 19068
rect 8268 19066 8324 19068
rect 8348 19066 8404 19068
rect 8108 19014 8154 19066
rect 8154 19014 8164 19066
rect 8188 19014 8218 19066
rect 8218 19014 8230 19066
rect 8230 19014 8244 19066
rect 8268 19014 8282 19066
rect 8282 19014 8294 19066
rect 8294 19014 8324 19066
rect 8348 19014 8358 19066
rect 8358 19014 8404 19066
rect 8108 19012 8164 19014
rect 8188 19012 8244 19014
rect 8268 19012 8324 19014
rect 8348 19012 8404 19014
rect 15813 19066 15869 19068
rect 15893 19066 15949 19068
rect 15973 19066 16029 19068
rect 16053 19066 16109 19068
rect 15813 19014 15859 19066
rect 15859 19014 15869 19066
rect 15893 19014 15923 19066
rect 15923 19014 15935 19066
rect 15935 19014 15949 19066
rect 15973 19014 15987 19066
rect 15987 19014 15999 19066
rect 15999 19014 16029 19066
rect 16053 19014 16063 19066
rect 16063 19014 16109 19066
rect 15813 19012 15869 19014
rect 15893 19012 15949 19014
rect 15973 19012 16029 19014
rect 16053 19012 16109 19014
rect 4256 18522 4312 18524
rect 4336 18522 4392 18524
rect 4416 18522 4472 18524
rect 4496 18522 4552 18524
rect 4256 18470 4302 18522
rect 4302 18470 4312 18522
rect 4336 18470 4366 18522
rect 4366 18470 4378 18522
rect 4378 18470 4392 18522
rect 4416 18470 4430 18522
rect 4430 18470 4442 18522
rect 4442 18470 4472 18522
rect 4496 18470 4506 18522
rect 4506 18470 4552 18522
rect 4256 18468 4312 18470
rect 4336 18468 4392 18470
rect 4416 18468 4472 18470
rect 4496 18468 4552 18470
rect 846 18400 902 18456
rect 846 17720 902 17776
rect 4256 17434 4312 17436
rect 4336 17434 4392 17436
rect 4416 17434 4472 17436
rect 4496 17434 4552 17436
rect 4256 17382 4302 17434
rect 4302 17382 4312 17434
rect 4336 17382 4366 17434
rect 4366 17382 4378 17434
rect 4378 17382 4392 17434
rect 4416 17382 4430 17434
rect 4430 17382 4442 17434
rect 4442 17382 4472 17434
rect 4496 17382 4506 17434
rect 4506 17382 4552 17434
rect 4256 17380 4312 17382
rect 4336 17380 4392 17382
rect 4416 17380 4472 17382
rect 4496 17380 4552 17382
rect 846 17076 848 17096
rect 848 17076 900 17096
rect 900 17076 902 17096
rect 846 17040 902 17076
rect 4256 16346 4312 16348
rect 4336 16346 4392 16348
rect 4416 16346 4472 16348
rect 4496 16346 4552 16348
rect 4256 16294 4302 16346
rect 4302 16294 4312 16346
rect 4336 16294 4366 16346
rect 4366 16294 4378 16346
rect 4378 16294 4392 16346
rect 4416 16294 4430 16346
rect 4430 16294 4442 16346
rect 4442 16294 4472 16346
rect 4496 16294 4506 16346
rect 4506 16294 4552 16346
rect 4256 16292 4312 16294
rect 4336 16292 4392 16294
rect 4416 16292 4472 16294
rect 4496 16292 4552 16294
rect 3054 13252 3110 13288
rect 3054 13232 3056 13252
rect 3056 13232 3108 13252
rect 3108 13232 3110 13252
rect 3054 12280 3110 12336
rect 4256 15258 4312 15260
rect 4336 15258 4392 15260
rect 4416 15258 4472 15260
rect 4496 15258 4552 15260
rect 4256 15206 4302 15258
rect 4302 15206 4312 15258
rect 4336 15206 4366 15258
rect 4366 15206 4378 15258
rect 4378 15206 4392 15258
rect 4416 15206 4430 15258
rect 4430 15206 4442 15258
rect 4442 15206 4472 15258
rect 4496 15206 4506 15258
rect 4506 15206 4552 15258
rect 4256 15204 4312 15206
rect 4336 15204 4392 15206
rect 4416 15204 4472 15206
rect 4496 15204 4552 15206
rect 4256 14170 4312 14172
rect 4336 14170 4392 14172
rect 4416 14170 4472 14172
rect 4496 14170 4552 14172
rect 4256 14118 4302 14170
rect 4302 14118 4312 14170
rect 4336 14118 4366 14170
rect 4366 14118 4378 14170
rect 4378 14118 4392 14170
rect 4416 14118 4430 14170
rect 4430 14118 4442 14170
rect 4442 14118 4472 14170
rect 4496 14118 4506 14170
rect 4506 14118 4552 14170
rect 4256 14116 4312 14118
rect 4336 14116 4392 14118
rect 4416 14116 4472 14118
rect 4496 14116 4552 14118
rect 4066 13368 4122 13424
rect 4256 13082 4312 13084
rect 4336 13082 4392 13084
rect 4416 13082 4472 13084
rect 4496 13082 4552 13084
rect 4256 13030 4302 13082
rect 4302 13030 4312 13082
rect 4336 13030 4366 13082
rect 4366 13030 4378 13082
rect 4378 13030 4392 13082
rect 4416 13030 4430 13082
rect 4430 13030 4442 13082
rect 4442 13030 4472 13082
rect 4496 13030 4506 13082
rect 4506 13030 4552 13082
rect 4256 13028 4312 13030
rect 4336 13028 4392 13030
rect 4416 13028 4472 13030
rect 4496 13028 4552 13030
rect 3974 12144 4030 12200
rect 4256 11994 4312 11996
rect 4336 11994 4392 11996
rect 4416 11994 4472 11996
rect 4496 11994 4552 11996
rect 4256 11942 4302 11994
rect 4302 11942 4312 11994
rect 4336 11942 4366 11994
rect 4366 11942 4378 11994
rect 4378 11942 4392 11994
rect 4416 11942 4430 11994
rect 4430 11942 4442 11994
rect 4442 11942 4472 11994
rect 4496 11942 4506 11994
rect 4506 11942 4552 11994
rect 4256 11940 4312 11942
rect 4336 11940 4392 11942
rect 4416 11940 4472 11942
rect 4496 11940 4552 11942
rect 4256 10906 4312 10908
rect 4336 10906 4392 10908
rect 4416 10906 4472 10908
rect 4496 10906 4552 10908
rect 4256 10854 4302 10906
rect 4302 10854 4312 10906
rect 4336 10854 4366 10906
rect 4366 10854 4378 10906
rect 4378 10854 4392 10906
rect 4416 10854 4430 10906
rect 4430 10854 4442 10906
rect 4442 10854 4472 10906
rect 4496 10854 4506 10906
rect 4506 10854 4552 10906
rect 4256 10852 4312 10854
rect 4336 10852 4392 10854
rect 4416 10852 4472 10854
rect 4496 10852 4552 10854
rect 4256 9818 4312 9820
rect 4336 9818 4392 9820
rect 4416 9818 4472 9820
rect 4496 9818 4552 9820
rect 4256 9766 4302 9818
rect 4302 9766 4312 9818
rect 4336 9766 4366 9818
rect 4366 9766 4378 9818
rect 4378 9766 4392 9818
rect 4416 9766 4430 9818
rect 4430 9766 4442 9818
rect 4442 9766 4472 9818
rect 4496 9766 4506 9818
rect 4506 9766 4552 9818
rect 4256 9764 4312 9766
rect 4336 9764 4392 9766
rect 4416 9764 4472 9766
rect 4496 9764 4552 9766
rect 5998 14864 6054 14920
rect 8108 17978 8164 17980
rect 8188 17978 8244 17980
rect 8268 17978 8324 17980
rect 8348 17978 8404 17980
rect 8108 17926 8154 17978
rect 8154 17926 8164 17978
rect 8188 17926 8218 17978
rect 8218 17926 8230 17978
rect 8230 17926 8244 17978
rect 8268 17926 8282 17978
rect 8282 17926 8294 17978
rect 8294 17926 8324 17978
rect 8348 17926 8358 17978
rect 8358 17926 8404 17978
rect 8108 17924 8164 17926
rect 8188 17924 8244 17926
rect 8268 17924 8324 17926
rect 8348 17924 8404 17926
rect 11961 18522 12017 18524
rect 12041 18522 12097 18524
rect 12121 18522 12177 18524
rect 12201 18522 12257 18524
rect 11961 18470 12007 18522
rect 12007 18470 12017 18522
rect 12041 18470 12071 18522
rect 12071 18470 12083 18522
rect 12083 18470 12097 18522
rect 12121 18470 12135 18522
rect 12135 18470 12147 18522
rect 12147 18470 12177 18522
rect 12201 18470 12211 18522
rect 12211 18470 12257 18522
rect 11961 18468 12017 18470
rect 12041 18468 12097 18470
rect 12121 18468 12177 18470
rect 12201 18468 12257 18470
rect 8108 16890 8164 16892
rect 8188 16890 8244 16892
rect 8268 16890 8324 16892
rect 8348 16890 8404 16892
rect 8108 16838 8154 16890
rect 8154 16838 8164 16890
rect 8188 16838 8218 16890
rect 8218 16838 8230 16890
rect 8230 16838 8244 16890
rect 8268 16838 8282 16890
rect 8282 16838 8294 16890
rect 8294 16838 8324 16890
rect 8348 16838 8358 16890
rect 8358 16838 8404 16890
rect 8108 16836 8164 16838
rect 8188 16836 8244 16838
rect 8268 16836 8324 16838
rect 8348 16836 8404 16838
rect 6826 12824 6882 12880
rect 6458 12144 6514 12200
rect 6274 11600 6330 11656
rect 4256 8730 4312 8732
rect 4336 8730 4392 8732
rect 4416 8730 4472 8732
rect 4496 8730 4552 8732
rect 4256 8678 4302 8730
rect 4302 8678 4312 8730
rect 4336 8678 4366 8730
rect 4366 8678 4378 8730
rect 4378 8678 4392 8730
rect 4416 8678 4430 8730
rect 4430 8678 4442 8730
rect 4442 8678 4472 8730
rect 4496 8678 4506 8730
rect 4506 8678 4552 8730
rect 4256 8676 4312 8678
rect 4336 8676 4392 8678
rect 4416 8676 4472 8678
rect 4496 8676 4552 8678
rect 8108 15802 8164 15804
rect 8188 15802 8244 15804
rect 8268 15802 8324 15804
rect 8348 15802 8404 15804
rect 8108 15750 8154 15802
rect 8154 15750 8164 15802
rect 8188 15750 8218 15802
rect 8218 15750 8230 15802
rect 8230 15750 8244 15802
rect 8268 15750 8282 15802
rect 8282 15750 8294 15802
rect 8294 15750 8324 15802
rect 8348 15750 8358 15802
rect 8358 15750 8404 15802
rect 8108 15748 8164 15750
rect 8188 15748 8244 15750
rect 8268 15748 8324 15750
rect 8348 15748 8404 15750
rect 8206 15036 8208 15056
rect 8208 15036 8260 15056
rect 8260 15036 8262 15056
rect 8206 15000 8262 15036
rect 8108 14714 8164 14716
rect 8188 14714 8244 14716
rect 8268 14714 8324 14716
rect 8348 14714 8404 14716
rect 8108 14662 8154 14714
rect 8154 14662 8164 14714
rect 8188 14662 8218 14714
rect 8218 14662 8230 14714
rect 8230 14662 8244 14714
rect 8268 14662 8282 14714
rect 8282 14662 8294 14714
rect 8294 14662 8324 14714
rect 8348 14662 8358 14714
rect 8358 14662 8404 14714
rect 8108 14660 8164 14662
rect 8188 14660 8244 14662
rect 8268 14660 8324 14662
rect 8348 14660 8404 14662
rect 8108 13626 8164 13628
rect 8188 13626 8244 13628
rect 8268 13626 8324 13628
rect 8348 13626 8404 13628
rect 8108 13574 8154 13626
rect 8154 13574 8164 13626
rect 8188 13574 8218 13626
rect 8218 13574 8230 13626
rect 8230 13574 8244 13626
rect 8268 13574 8282 13626
rect 8282 13574 8294 13626
rect 8294 13574 8324 13626
rect 8348 13574 8358 13626
rect 8358 13574 8404 13626
rect 8108 13572 8164 13574
rect 8188 13572 8244 13574
rect 8268 13572 8324 13574
rect 8348 13572 8404 13574
rect 8108 12538 8164 12540
rect 8188 12538 8244 12540
rect 8268 12538 8324 12540
rect 8348 12538 8404 12540
rect 8108 12486 8154 12538
rect 8154 12486 8164 12538
rect 8188 12486 8218 12538
rect 8218 12486 8230 12538
rect 8230 12486 8244 12538
rect 8268 12486 8282 12538
rect 8282 12486 8294 12538
rect 8294 12486 8324 12538
rect 8348 12486 8358 12538
rect 8358 12486 8404 12538
rect 8108 12484 8164 12486
rect 8188 12484 8244 12486
rect 8268 12484 8324 12486
rect 8348 12484 8404 12486
rect 8114 11600 8170 11656
rect 8108 11450 8164 11452
rect 8188 11450 8244 11452
rect 8268 11450 8324 11452
rect 8348 11450 8404 11452
rect 8108 11398 8154 11450
rect 8154 11398 8164 11450
rect 8188 11398 8218 11450
rect 8218 11398 8230 11450
rect 8230 11398 8244 11450
rect 8268 11398 8282 11450
rect 8282 11398 8294 11450
rect 8294 11398 8324 11450
rect 8348 11398 8358 11450
rect 8358 11398 8404 11450
rect 8108 11396 8164 11398
rect 8188 11396 8244 11398
rect 8268 11396 8324 11398
rect 8348 11396 8404 11398
rect 7930 10648 7986 10704
rect 11961 17434 12017 17436
rect 12041 17434 12097 17436
rect 12121 17434 12177 17436
rect 12201 17434 12257 17436
rect 11961 17382 12007 17434
rect 12007 17382 12017 17434
rect 12041 17382 12071 17434
rect 12071 17382 12083 17434
rect 12083 17382 12097 17434
rect 12121 17382 12135 17434
rect 12135 17382 12147 17434
rect 12147 17382 12177 17434
rect 12201 17382 12211 17434
rect 12211 17382 12257 17434
rect 11961 17380 12017 17382
rect 12041 17380 12097 17382
rect 12121 17380 12177 17382
rect 12201 17380 12257 17382
rect 11961 16346 12017 16348
rect 12041 16346 12097 16348
rect 12121 16346 12177 16348
rect 12201 16346 12257 16348
rect 11961 16294 12007 16346
rect 12007 16294 12017 16346
rect 12041 16294 12071 16346
rect 12071 16294 12083 16346
rect 12083 16294 12097 16346
rect 12121 16294 12135 16346
rect 12135 16294 12147 16346
rect 12147 16294 12177 16346
rect 12201 16294 12211 16346
rect 12211 16294 12257 16346
rect 11961 16292 12017 16294
rect 12041 16292 12097 16294
rect 12121 16292 12177 16294
rect 12201 16292 12257 16294
rect 11961 15258 12017 15260
rect 12041 15258 12097 15260
rect 12121 15258 12177 15260
rect 12201 15258 12257 15260
rect 11961 15206 12007 15258
rect 12007 15206 12017 15258
rect 12041 15206 12071 15258
rect 12071 15206 12083 15258
rect 12083 15206 12097 15258
rect 12121 15206 12135 15258
rect 12135 15206 12147 15258
rect 12147 15206 12177 15258
rect 12201 15206 12211 15258
rect 12211 15206 12257 15258
rect 11961 15204 12017 15206
rect 12041 15204 12097 15206
rect 12121 15204 12177 15206
rect 12201 15204 12257 15206
rect 11242 13676 11244 13696
rect 11244 13676 11296 13696
rect 11296 13676 11298 13696
rect 11242 13640 11298 13676
rect 10874 12688 10930 12744
rect 10046 12416 10102 12472
rect 11961 14170 12017 14172
rect 12041 14170 12097 14172
rect 12121 14170 12177 14172
rect 12201 14170 12257 14172
rect 11961 14118 12007 14170
rect 12007 14118 12017 14170
rect 12041 14118 12071 14170
rect 12071 14118 12083 14170
rect 12083 14118 12097 14170
rect 12121 14118 12135 14170
rect 12135 14118 12147 14170
rect 12147 14118 12177 14170
rect 12201 14118 12211 14170
rect 12211 14118 12257 14170
rect 11961 14116 12017 14118
rect 12041 14116 12097 14118
rect 12121 14116 12177 14118
rect 12201 14116 12257 14118
rect 11794 13504 11850 13560
rect 9678 11056 9734 11112
rect 7746 9016 7802 9072
rect 7378 8472 7434 8528
rect 4256 7642 4312 7644
rect 4336 7642 4392 7644
rect 4416 7642 4472 7644
rect 4496 7642 4552 7644
rect 4256 7590 4302 7642
rect 4302 7590 4312 7642
rect 4336 7590 4366 7642
rect 4366 7590 4378 7642
rect 4378 7590 4392 7642
rect 4416 7590 4430 7642
rect 4430 7590 4442 7642
rect 4442 7590 4472 7642
rect 4496 7590 4506 7642
rect 4506 7590 4552 7642
rect 4256 7588 4312 7590
rect 4336 7588 4392 7590
rect 4416 7588 4472 7590
rect 4496 7588 4552 7590
rect 4256 6554 4312 6556
rect 4336 6554 4392 6556
rect 4416 6554 4472 6556
rect 4496 6554 4552 6556
rect 4256 6502 4302 6554
rect 4302 6502 4312 6554
rect 4336 6502 4366 6554
rect 4366 6502 4378 6554
rect 4378 6502 4392 6554
rect 4416 6502 4430 6554
rect 4430 6502 4442 6554
rect 4442 6502 4472 6554
rect 4496 6502 4506 6554
rect 4506 6502 4552 6554
rect 4256 6500 4312 6502
rect 4336 6500 4392 6502
rect 4416 6500 4472 6502
rect 4496 6500 4552 6502
rect 4618 6160 4674 6216
rect 4256 5466 4312 5468
rect 4336 5466 4392 5468
rect 4416 5466 4472 5468
rect 4496 5466 4552 5468
rect 4256 5414 4302 5466
rect 4302 5414 4312 5466
rect 4336 5414 4366 5466
rect 4366 5414 4378 5466
rect 4378 5414 4392 5466
rect 4416 5414 4430 5466
rect 4430 5414 4442 5466
rect 4442 5414 4472 5466
rect 4496 5414 4506 5466
rect 4506 5414 4552 5466
rect 4256 5412 4312 5414
rect 4336 5412 4392 5414
rect 4416 5412 4472 5414
rect 4496 5412 4552 5414
rect 8108 10362 8164 10364
rect 8188 10362 8244 10364
rect 8268 10362 8324 10364
rect 8348 10362 8404 10364
rect 8108 10310 8154 10362
rect 8154 10310 8164 10362
rect 8188 10310 8218 10362
rect 8218 10310 8230 10362
rect 8230 10310 8244 10362
rect 8268 10310 8282 10362
rect 8282 10310 8294 10362
rect 8294 10310 8324 10362
rect 8348 10310 8358 10362
rect 8358 10310 8404 10362
rect 8108 10308 8164 10310
rect 8188 10308 8244 10310
rect 8268 10308 8324 10310
rect 8348 10308 8404 10310
rect 8108 9274 8164 9276
rect 8188 9274 8244 9276
rect 8268 9274 8324 9276
rect 8348 9274 8404 9276
rect 8108 9222 8154 9274
rect 8154 9222 8164 9274
rect 8188 9222 8218 9274
rect 8218 9222 8230 9274
rect 8230 9222 8244 9274
rect 8268 9222 8282 9274
rect 8282 9222 8294 9274
rect 8294 9222 8324 9274
rect 8348 9222 8358 9274
rect 8358 9222 8404 9274
rect 8108 9220 8164 9222
rect 8188 9220 8244 9222
rect 8268 9220 8324 9222
rect 8348 9220 8404 9222
rect 8108 8186 8164 8188
rect 8188 8186 8244 8188
rect 8268 8186 8324 8188
rect 8348 8186 8404 8188
rect 8108 8134 8154 8186
rect 8154 8134 8164 8186
rect 8188 8134 8218 8186
rect 8218 8134 8230 8186
rect 8230 8134 8244 8186
rect 8268 8134 8282 8186
rect 8282 8134 8294 8186
rect 8294 8134 8324 8186
rect 8348 8134 8358 8186
rect 8358 8134 8404 8186
rect 8108 8132 8164 8134
rect 8188 8132 8244 8134
rect 8268 8132 8324 8134
rect 8348 8132 8404 8134
rect 8108 7098 8164 7100
rect 8188 7098 8244 7100
rect 8268 7098 8324 7100
rect 8348 7098 8404 7100
rect 8108 7046 8154 7098
rect 8154 7046 8164 7098
rect 8188 7046 8218 7098
rect 8218 7046 8230 7098
rect 8230 7046 8244 7098
rect 8268 7046 8282 7098
rect 8282 7046 8294 7098
rect 8294 7046 8324 7098
rect 8348 7046 8358 7098
rect 8358 7046 8404 7098
rect 8108 7044 8164 7046
rect 8188 7044 8244 7046
rect 8268 7044 8324 7046
rect 8348 7044 8404 7046
rect 11961 13082 12017 13084
rect 12041 13082 12097 13084
rect 12121 13082 12177 13084
rect 12201 13082 12257 13084
rect 11961 13030 12007 13082
rect 12007 13030 12017 13082
rect 12041 13030 12071 13082
rect 12071 13030 12083 13082
rect 12083 13030 12097 13082
rect 12121 13030 12135 13082
rect 12135 13030 12147 13082
rect 12147 13030 12177 13082
rect 12201 13030 12211 13082
rect 12211 13030 12257 13082
rect 11961 13028 12017 13030
rect 12041 13028 12097 13030
rect 12121 13028 12177 13030
rect 12201 13028 12257 13030
rect 11242 10512 11298 10568
rect 10046 10376 10102 10432
rect 11961 11994 12017 11996
rect 12041 11994 12097 11996
rect 12121 11994 12177 11996
rect 12201 11994 12257 11996
rect 11961 11942 12007 11994
rect 12007 11942 12017 11994
rect 12041 11942 12071 11994
rect 12071 11942 12083 11994
rect 12083 11942 12097 11994
rect 12121 11942 12135 11994
rect 12135 11942 12147 11994
rect 12147 11942 12177 11994
rect 12201 11942 12211 11994
rect 12211 11942 12257 11994
rect 11961 11940 12017 11942
rect 12041 11940 12097 11942
rect 12121 11940 12177 11942
rect 12201 11940 12257 11942
rect 11978 11464 12034 11520
rect 11961 10906 12017 10908
rect 12041 10906 12097 10908
rect 12121 10906 12177 10908
rect 12201 10906 12257 10908
rect 11961 10854 12007 10906
rect 12007 10854 12017 10906
rect 12041 10854 12071 10906
rect 12071 10854 12083 10906
rect 12083 10854 12097 10906
rect 12121 10854 12135 10906
rect 12135 10854 12147 10906
rect 12147 10854 12177 10906
rect 12201 10854 12211 10906
rect 12211 10854 12257 10906
rect 11961 10852 12017 10854
rect 12041 10852 12097 10854
rect 12121 10852 12177 10854
rect 12201 10852 12257 10854
rect 11961 9818 12017 9820
rect 12041 9818 12097 9820
rect 12121 9818 12177 9820
rect 12201 9818 12257 9820
rect 11961 9766 12007 9818
rect 12007 9766 12017 9818
rect 12041 9766 12071 9818
rect 12071 9766 12083 9818
rect 12083 9766 12097 9818
rect 12121 9766 12135 9818
rect 12135 9766 12147 9818
rect 12147 9766 12177 9818
rect 12201 9766 12211 9818
rect 12211 9766 12257 9818
rect 11961 9764 12017 9766
rect 12041 9764 12097 9766
rect 12121 9764 12177 9766
rect 12201 9764 12257 9766
rect 15014 17992 15070 18048
rect 15813 17978 15869 17980
rect 15893 17978 15949 17980
rect 15973 17978 16029 17980
rect 16053 17978 16109 17980
rect 15813 17926 15859 17978
rect 15859 17926 15869 17978
rect 15893 17926 15923 17978
rect 15923 17926 15935 17978
rect 15935 17926 15949 17978
rect 15973 17926 15987 17978
rect 15987 17926 15999 17978
rect 15999 17926 16029 17978
rect 16053 17926 16063 17978
rect 16063 17926 16109 17978
rect 15813 17924 15869 17926
rect 15893 17924 15949 17926
rect 15973 17924 16029 17926
rect 16053 17924 16109 17926
rect 12438 9832 12494 9888
rect 8108 6010 8164 6012
rect 8188 6010 8244 6012
rect 8268 6010 8324 6012
rect 8348 6010 8404 6012
rect 8108 5958 8154 6010
rect 8154 5958 8164 6010
rect 8188 5958 8218 6010
rect 8218 5958 8230 6010
rect 8230 5958 8244 6010
rect 8268 5958 8282 6010
rect 8282 5958 8294 6010
rect 8294 5958 8324 6010
rect 8348 5958 8358 6010
rect 8358 5958 8404 6010
rect 8108 5956 8164 5958
rect 8188 5956 8244 5958
rect 8268 5956 8324 5958
rect 8348 5956 8404 5958
rect 9218 5364 9274 5400
rect 9218 5344 9220 5364
rect 9220 5344 9272 5364
rect 9272 5344 9274 5364
rect 8108 4922 8164 4924
rect 8188 4922 8244 4924
rect 8268 4922 8324 4924
rect 8348 4922 8404 4924
rect 8108 4870 8154 4922
rect 8154 4870 8164 4922
rect 8188 4870 8218 4922
rect 8218 4870 8230 4922
rect 8230 4870 8244 4922
rect 8268 4870 8282 4922
rect 8282 4870 8294 4922
rect 8294 4870 8324 4922
rect 8348 4870 8358 4922
rect 8358 4870 8404 4922
rect 8108 4868 8164 4870
rect 8188 4868 8244 4870
rect 8268 4868 8324 4870
rect 8348 4868 8404 4870
rect 7194 4664 7250 4720
rect 4894 4548 4950 4584
rect 4894 4528 4896 4548
rect 4896 4528 4948 4548
rect 4948 4528 4950 4548
rect 4256 4378 4312 4380
rect 4336 4378 4392 4380
rect 4416 4378 4472 4380
rect 4496 4378 4552 4380
rect 4256 4326 4302 4378
rect 4302 4326 4312 4378
rect 4336 4326 4366 4378
rect 4366 4326 4378 4378
rect 4378 4326 4392 4378
rect 4416 4326 4430 4378
rect 4430 4326 4442 4378
rect 4442 4326 4472 4378
rect 4496 4326 4506 4378
rect 4506 4326 4552 4378
rect 4256 4324 4312 4326
rect 4336 4324 4392 4326
rect 4416 4324 4472 4326
rect 4496 4324 4552 4326
rect 4256 3290 4312 3292
rect 4336 3290 4392 3292
rect 4416 3290 4472 3292
rect 4496 3290 4552 3292
rect 4256 3238 4302 3290
rect 4302 3238 4312 3290
rect 4336 3238 4366 3290
rect 4366 3238 4378 3290
rect 4378 3238 4392 3290
rect 4416 3238 4430 3290
rect 4430 3238 4442 3290
rect 4442 3238 4472 3290
rect 4496 3238 4506 3290
rect 4506 3238 4552 3290
rect 4256 3236 4312 3238
rect 4336 3236 4392 3238
rect 4416 3236 4472 3238
rect 4496 3236 4552 3238
rect 10414 5364 10470 5400
rect 10414 5344 10416 5364
rect 10416 5344 10468 5364
rect 10468 5344 10470 5364
rect 8108 3834 8164 3836
rect 8188 3834 8244 3836
rect 8268 3834 8324 3836
rect 8348 3834 8404 3836
rect 8108 3782 8154 3834
rect 8154 3782 8164 3834
rect 8188 3782 8218 3834
rect 8218 3782 8230 3834
rect 8230 3782 8244 3834
rect 8268 3782 8282 3834
rect 8282 3782 8294 3834
rect 8294 3782 8324 3834
rect 8348 3782 8358 3834
rect 8358 3782 8404 3834
rect 8108 3780 8164 3782
rect 8188 3780 8244 3782
rect 8268 3780 8324 3782
rect 8348 3780 8404 3782
rect 5262 2896 5318 2952
rect 4256 2202 4312 2204
rect 4336 2202 4392 2204
rect 4416 2202 4472 2204
rect 4496 2202 4552 2204
rect 4256 2150 4302 2202
rect 4302 2150 4312 2202
rect 4336 2150 4366 2202
rect 4366 2150 4378 2202
rect 4378 2150 4392 2202
rect 4416 2150 4430 2202
rect 4430 2150 4442 2202
rect 4442 2150 4472 2202
rect 4496 2150 4506 2202
rect 4506 2150 4552 2202
rect 4256 2148 4312 2150
rect 4336 2148 4392 2150
rect 4416 2148 4472 2150
rect 4496 2148 4552 2150
rect 8108 2746 8164 2748
rect 8188 2746 8244 2748
rect 8268 2746 8324 2748
rect 8348 2746 8404 2748
rect 8108 2694 8154 2746
rect 8154 2694 8164 2746
rect 8188 2694 8218 2746
rect 8218 2694 8230 2746
rect 8230 2694 8244 2746
rect 8268 2694 8282 2746
rect 8282 2694 8294 2746
rect 8294 2694 8324 2746
rect 8348 2694 8358 2746
rect 8358 2694 8404 2746
rect 8108 2692 8164 2694
rect 8188 2692 8244 2694
rect 8268 2692 8324 2694
rect 8348 2692 8404 2694
rect 11610 5888 11666 5944
rect 11961 8730 12017 8732
rect 12041 8730 12097 8732
rect 12121 8730 12177 8732
rect 12201 8730 12257 8732
rect 11961 8678 12007 8730
rect 12007 8678 12017 8730
rect 12041 8678 12071 8730
rect 12071 8678 12083 8730
rect 12083 8678 12097 8730
rect 12121 8678 12135 8730
rect 12135 8678 12147 8730
rect 12147 8678 12177 8730
rect 12201 8678 12211 8730
rect 12211 8678 12257 8730
rect 11961 8676 12017 8678
rect 12041 8676 12097 8678
rect 12121 8676 12177 8678
rect 12201 8676 12257 8678
rect 11961 7642 12017 7644
rect 12041 7642 12097 7644
rect 12121 7642 12177 7644
rect 12201 7642 12257 7644
rect 11961 7590 12007 7642
rect 12007 7590 12017 7642
rect 12041 7590 12071 7642
rect 12071 7590 12083 7642
rect 12083 7590 12097 7642
rect 12121 7590 12135 7642
rect 12135 7590 12147 7642
rect 12147 7590 12177 7642
rect 12201 7590 12211 7642
rect 12211 7590 12257 7642
rect 11961 7588 12017 7590
rect 12041 7588 12097 7590
rect 12121 7588 12177 7590
rect 12201 7588 12257 7590
rect 12714 8608 12770 8664
rect 12714 8372 12716 8392
rect 12716 8372 12768 8392
rect 12768 8372 12770 8392
rect 12714 8336 12770 8372
rect 13634 13096 13690 13152
rect 13266 9696 13322 9752
rect 12254 6724 12310 6760
rect 12254 6704 12256 6724
rect 12256 6704 12308 6724
rect 12308 6704 12310 6724
rect 11961 6554 12017 6556
rect 12041 6554 12097 6556
rect 12121 6554 12177 6556
rect 12201 6554 12257 6556
rect 11961 6502 12007 6554
rect 12007 6502 12017 6554
rect 12041 6502 12071 6554
rect 12071 6502 12083 6554
rect 12083 6502 12097 6554
rect 12121 6502 12135 6554
rect 12135 6502 12147 6554
rect 12147 6502 12177 6554
rect 12201 6502 12211 6554
rect 12211 6502 12257 6554
rect 11961 6500 12017 6502
rect 12041 6500 12097 6502
rect 12121 6500 12177 6502
rect 12201 6500 12257 6502
rect 12806 6976 12862 7032
rect 13082 6296 13138 6352
rect 12530 6160 12586 6216
rect 11961 5466 12017 5468
rect 12041 5466 12097 5468
rect 12121 5466 12177 5468
rect 12201 5466 12257 5468
rect 11961 5414 12007 5466
rect 12007 5414 12017 5466
rect 12041 5414 12071 5466
rect 12071 5414 12083 5466
rect 12083 5414 12097 5466
rect 12121 5414 12135 5466
rect 12135 5414 12147 5466
rect 12147 5414 12177 5466
rect 12201 5414 12211 5466
rect 12211 5414 12257 5466
rect 11961 5412 12017 5414
rect 12041 5412 12097 5414
rect 12121 5412 12177 5414
rect 12201 5412 12257 5414
rect 11961 4378 12017 4380
rect 12041 4378 12097 4380
rect 12121 4378 12177 4380
rect 12201 4378 12257 4380
rect 11961 4326 12007 4378
rect 12007 4326 12017 4378
rect 12041 4326 12071 4378
rect 12071 4326 12083 4378
rect 12083 4326 12097 4378
rect 12121 4326 12135 4378
rect 12135 4326 12147 4378
rect 12147 4326 12177 4378
rect 12201 4326 12211 4378
rect 12211 4326 12257 4378
rect 11961 4324 12017 4326
rect 12041 4324 12097 4326
rect 12121 4324 12177 4326
rect 12201 4324 12257 4326
rect 11978 3712 12034 3768
rect 4256 1114 4312 1116
rect 4336 1114 4392 1116
rect 4416 1114 4472 1116
rect 4496 1114 4552 1116
rect 4256 1062 4302 1114
rect 4302 1062 4312 1114
rect 4336 1062 4366 1114
rect 4366 1062 4378 1114
rect 4378 1062 4392 1114
rect 4416 1062 4430 1114
rect 4430 1062 4442 1114
rect 4442 1062 4472 1114
rect 4496 1062 4506 1114
rect 4506 1062 4552 1114
rect 4256 1060 4312 1062
rect 4336 1060 4392 1062
rect 4416 1060 4472 1062
rect 4496 1060 4552 1062
rect 8108 1658 8164 1660
rect 8188 1658 8244 1660
rect 8268 1658 8324 1660
rect 8348 1658 8404 1660
rect 8108 1606 8154 1658
rect 8154 1606 8164 1658
rect 8188 1606 8218 1658
rect 8218 1606 8230 1658
rect 8230 1606 8244 1658
rect 8268 1606 8282 1658
rect 8282 1606 8294 1658
rect 8294 1606 8324 1658
rect 8348 1606 8358 1658
rect 8358 1606 8404 1658
rect 8108 1604 8164 1606
rect 8188 1604 8244 1606
rect 8268 1604 8324 1606
rect 8348 1604 8404 1606
rect 11961 3290 12017 3292
rect 12041 3290 12097 3292
rect 12121 3290 12177 3292
rect 12201 3290 12257 3292
rect 11961 3238 12007 3290
rect 12007 3238 12017 3290
rect 12041 3238 12071 3290
rect 12071 3238 12083 3290
rect 12083 3238 12097 3290
rect 12121 3238 12135 3290
rect 12135 3238 12147 3290
rect 12147 3238 12177 3290
rect 12201 3238 12211 3290
rect 12211 3238 12257 3290
rect 11961 3236 12017 3238
rect 12041 3236 12097 3238
rect 12121 3236 12177 3238
rect 12201 3236 12257 3238
rect 12530 3576 12586 3632
rect 11961 2202 12017 2204
rect 12041 2202 12097 2204
rect 12121 2202 12177 2204
rect 12201 2202 12257 2204
rect 11961 2150 12007 2202
rect 12007 2150 12017 2202
rect 12041 2150 12071 2202
rect 12071 2150 12083 2202
rect 12083 2150 12097 2202
rect 12121 2150 12135 2202
rect 12135 2150 12147 2202
rect 12147 2150 12177 2202
rect 12201 2150 12211 2202
rect 12211 2150 12257 2202
rect 11961 2148 12017 2150
rect 12041 2148 12097 2150
rect 12121 2148 12177 2150
rect 12201 2148 12257 2150
rect 11961 1114 12017 1116
rect 12041 1114 12097 1116
rect 12121 1114 12177 1116
rect 12201 1114 12257 1116
rect 11961 1062 12007 1114
rect 12007 1062 12017 1114
rect 12041 1062 12071 1114
rect 12071 1062 12083 1114
rect 12083 1062 12097 1114
rect 12121 1062 12135 1114
rect 12135 1062 12147 1114
rect 12147 1062 12177 1114
rect 12201 1062 12211 1114
rect 12211 1062 12257 1114
rect 11961 1060 12017 1062
rect 12041 1060 12097 1062
rect 12121 1060 12177 1062
rect 12201 1060 12257 1062
rect 13450 8900 13506 8936
rect 13450 8880 13452 8900
rect 13452 8880 13504 8900
rect 13504 8880 13506 8900
rect 13450 8064 13506 8120
rect 13266 4392 13322 4448
rect 13910 13640 13966 13696
rect 13910 12552 13966 12608
rect 13910 12416 13966 12472
rect 14278 12824 14334 12880
rect 13818 11736 13874 11792
rect 14186 11464 14242 11520
rect 15014 14492 15016 14512
rect 15016 14492 15068 14512
rect 15068 14492 15070 14512
rect 15014 14456 15070 14492
rect 14738 10648 14794 10704
rect 14002 10240 14058 10296
rect 13726 6840 13782 6896
rect 13634 5072 13690 5128
rect 14186 10376 14242 10432
rect 14278 10124 14334 10160
rect 15014 11736 15070 11792
rect 14278 10104 14280 10124
rect 14280 10104 14332 10124
rect 14332 10104 14334 10124
rect 14278 9968 14334 10024
rect 14278 9424 14334 9480
rect 14002 6452 14058 6488
rect 14002 6432 14004 6452
rect 14004 6432 14056 6452
rect 14056 6432 14058 6452
rect 14278 7928 14334 7984
rect 14646 9868 14648 9888
rect 14648 9868 14700 9888
rect 14700 9868 14702 9888
rect 14646 9832 14702 9868
rect 14554 8628 14610 8664
rect 14554 8608 14556 8628
rect 14556 8608 14608 8628
rect 14608 8608 14610 8628
rect 14554 8064 14610 8120
rect 14922 9716 14978 9752
rect 14922 9696 14924 9716
rect 14924 9696 14976 9716
rect 14976 9696 14978 9716
rect 14922 9560 14978 9616
rect 15813 16890 15869 16892
rect 15893 16890 15949 16892
rect 15973 16890 16029 16892
rect 16053 16890 16109 16892
rect 15813 16838 15859 16890
rect 15859 16838 15869 16890
rect 15893 16838 15923 16890
rect 15923 16838 15935 16890
rect 15935 16838 15949 16890
rect 15973 16838 15987 16890
rect 15987 16838 15999 16890
rect 15999 16838 16029 16890
rect 16053 16838 16063 16890
rect 16063 16838 16109 16890
rect 15813 16836 15869 16838
rect 15893 16836 15949 16838
rect 15973 16836 16029 16838
rect 16053 16836 16109 16838
rect 16026 15952 16082 16008
rect 15813 15802 15869 15804
rect 15893 15802 15949 15804
rect 15973 15802 16029 15804
rect 16053 15802 16109 15804
rect 15813 15750 15859 15802
rect 15859 15750 15869 15802
rect 15893 15750 15923 15802
rect 15923 15750 15935 15802
rect 15935 15750 15949 15802
rect 15973 15750 15987 15802
rect 15987 15750 15999 15802
rect 15999 15750 16029 15802
rect 16053 15750 16063 15802
rect 16063 15750 16109 15802
rect 15813 15748 15869 15750
rect 15893 15748 15949 15750
rect 15973 15748 16029 15750
rect 16053 15748 16109 15750
rect 15813 14714 15869 14716
rect 15893 14714 15949 14716
rect 15973 14714 16029 14716
rect 16053 14714 16109 14716
rect 15813 14662 15859 14714
rect 15859 14662 15869 14714
rect 15893 14662 15923 14714
rect 15923 14662 15935 14714
rect 15935 14662 15949 14714
rect 15973 14662 15987 14714
rect 15987 14662 15999 14714
rect 15999 14662 16029 14714
rect 16053 14662 16063 14714
rect 16063 14662 16109 14714
rect 15813 14660 15869 14662
rect 15893 14660 15949 14662
rect 15973 14660 16029 14662
rect 16053 14660 16109 14662
rect 15813 13626 15869 13628
rect 15893 13626 15949 13628
rect 15973 13626 16029 13628
rect 16053 13626 16109 13628
rect 15813 13574 15859 13626
rect 15859 13574 15869 13626
rect 15893 13574 15923 13626
rect 15923 13574 15935 13626
rect 15935 13574 15949 13626
rect 15973 13574 15987 13626
rect 15987 13574 15999 13626
rect 15999 13574 16029 13626
rect 16053 13574 16063 13626
rect 16063 13574 16109 13626
rect 15813 13572 15869 13574
rect 15893 13572 15949 13574
rect 15973 13572 16029 13574
rect 16053 13572 16109 13574
rect 15566 13232 15622 13288
rect 15658 13096 15714 13152
rect 15474 12436 15530 12472
rect 15474 12416 15476 12436
rect 15476 12416 15528 12436
rect 15528 12416 15530 12436
rect 15813 12538 15869 12540
rect 15893 12538 15949 12540
rect 15973 12538 16029 12540
rect 16053 12538 16109 12540
rect 15813 12486 15859 12538
rect 15859 12486 15869 12538
rect 15893 12486 15923 12538
rect 15923 12486 15935 12538
rect 15935 12486 15949 12538
rect 15973 12486 15987 12538
rect 15987 12486 15999 12538
rect 15999 12486 16029 12538
rect 16053 12486 16063 12538
rect 16063 12486 16109 12538
rect 15813 12484 15869 12486
rect 15893 12484 15949 12486
rect 15973 12484 16029 12486
rect 16053 12484 16109 12486
rect 16026 12280 16082 12336
rect 15198 12008 15254 12064
rect 15290 9696 15346 9752
rect 15198 9444 15254 9480
rect 15198 9424 15200 9444
rect 15200 9424 15252 9444
rect 15252 9424 15254 9444
rect 15934 12164 15990 12200
rect 15934 12144 15936 12164
rect 15936 12144 15988 12164
rect 15988 12144 15990 12164
rect 16026 11736 16082 11792
rect 16210 11464 16266 11520
rect 15813 11450 15869 11452
rect 15893 11450 15949 11452
rect 15973 11450 16029 11452
rect 16053 11450 16109 11452
rect 15813 11398 15859 11450
rect 15859 11398 15869 11450
rect 15893 11398 15923 11450
rect 15923 11398 15935 11450
rect 15935 11398 15949 11450
rect 15973 11398 15987 11450
rect 15987 11398 15999 11450
rect 15999 11398 16029 11450
rect 16053 11398 16063 11450
rect 16063 11398 16109 11450
rect 15813 11396 15869 11398
rect 15893 11396 15949 11398
rect 15973 11396 16029 11398
rect 16053 11396 16109 11398
rect 15658 11328 15714 11384
rect 16762 13812 16764 13832
rect 16764 13812 16816 13832
rect 16816 13812 16818 13832
rect 16762 13776 16818 13812
rect 16486 13096 16542 13152
rect 16486 12416 16542 12472
rect 15750 10784 15806 10840
rect 15750 10512 15806 10568
rect 15934 10548 15936 10568
rect 15936 10548 15988 10568
rect 15988 10548 15990 10568
rect 15934 10512 15990 10548
rect 16762 13368 16818 13424
rect 16854 12960 16910 13016
rect 16210 10376 16266 10432
rect 15813 10362 15869 10364
rect 15893 10362 15949 10364
rect 15973 10362 16029 10364
rect 16053 10362 16109 10364
rect 15813 10310 15859 10362
rect 15859 10310 15869 10362
rect 15893 10310 15923 10362
rect 15923 10310 15935 10362
rect 15935 10310 15949 10362
rect 15973 10310 15987 10362
rect 15987 10310 15999 10362
rect 15999 10310 16029 10362
rect 16053 10310 16063 10362
rect 16063 10310 16109 10362
rect 15813 10308 15869 10310
rect 15893 10308 15949 10310
rect 15973 10308 16029 10310
rect 16053 10308 16109 10310
rect 16302 10240 16358 10296
rect 15750 9832 15806 9888
rect 15474 8372 15476 8392
rect 15476 8372 15528 8392
rect 15528 8372 15530 8392
rect 14922 7792 14978 7848
rect 14462 6160 14518 6216
rect 14370 5888 14426 5944
rect 14278 3712 14334 3768
rect 15106 6976 15162 7032
rect 14646 4120 14702 4176
rect 15474 8336 15530 8372
rect 16118 9560 16174 9616
rect 15750 9444 15806 9480
rect 15750 9424 15752 9444
rect 15752 9424 15804 9444
rect 15804 9424 15806 9444
rect 16578 11464 16634 11520
rect 16854 11736 16910 11792
rect 16762 11464 16818 11520
rect 16854 11056 16910 11112
rect 16578 10784 16634 10840
rect 16762 10784 16818 10840
rect 16670 9560 16726 9616
rect 15813 9274 15869 9276
rect 15893 9274 15949 9276
rect 15973 9274 16029 9276
rect 16053 9274 16109 9276
rect 15813 9222 15859 9274
rect 15859 9222 15869 9274
rect 15893 9222 15923 9274
rect 15923 9222 15935 9274
rect 15935 9222 15949 9274
rect 15973 9222 15987 9274
rect 15987 9222 15999 9274
rect 15999 9222 16029 9274
rect 16053 9222 16063 9274
rect 16063 9222 16109 9274
rect 15813 9220 15869 9222
rect 15893 9220 15949 9222
rect 15973 9220 16029 9222
rect 16053 9220 16109 9222
rect 15813 8186 15869 8188
rect 15893 8186 15949 8188
rect 15973 8186 16029 8188
rect 16053 8186 16109 8188
rect 15813 8134 15859 8186
rect 15859 8134 15869 8186
rect 15893 8134 15923 8186
rect 15923 8134 15935 8186
rect 15935 8134 15949 8186
rect 15973 8134 15987 8186
rect 15987 8134 15999 8186
rect 15999 8134 16029 8186
rect 16053 8134 16063 8186
rect 16063 8134 16109 8186
rect 15813 8132 15869 8134
rect 15893 8132 15949 8134
rect 15973 8132 16029 8134
rect 16053 8132 16109 8134
rect 16394 9152 16450 9208
rect 16670 8744 16726 8800
rect 16578 8608 16634 8664
rect 17038 11212 17094 11248
rect 17038 11192 17040 11212
rect 17040 11192 17092 11212
rect 17092 11192 17094 11212
rect 17222 10920 17278 10976
rect 17774 16632 17830 16688
rect 17682 15000 17738 15056
rect 17866 14592 17922 14648
rect 17406 11328 17462 11384
rect 17774 13096 17830 13152
rect 18694 14900 18696 14920
rect 18696 14900 18748 14920
rect 18748 14900 18750 14920
rect 18694 14864 18750 14900
rect 18878 14456 18934 14512
rect 17774 12724 17776 12744
rect 17776 12724 17828 12744
rect 17828 12724 17830 12744
rect 17774 12688 17830 12724
rect 17682 11464 17738 11520
rect 17406 10920 17462 10976
rect 17222 10104 17278 10160
rect 17590 9560 17646 9616
rect 17774 10104 17830 10160
rect 18142 12280 18198 12336
rect 18142 10240 18198 10296
rect 18694 13640 18750 13696
rect 18602 12416 18658 12472
rect 18418 11872 18474 11928
rect 18326 10648 18382 10704
rect 16578 7792 16634 7848
rect 15813 7098 15869 7100
rect 15893 7098 15949 7100
rect 15973 7098 16029 7100
rect 16053 7098 16109 7100
rect 15813 7046 15859 7098
rect 15859 7046 15869 7098
rect 15893 7046 15923 7098
rect 15923 7046 15935 7098
rect 15935 7046 15949 7098
rect 15973 7046 15987 7098
rect 15987 7046 15999 7098
rect 15999 7046 16029 7098
rect 16053 7046 16063 7098
rect 16063 7046 16109 7098
rect 15813 7044 15869 7046
rect 15893 7044 15949 7046
rect 15973 7044 16029 7046
rect 16053 7044 16109 7046
rect 15813 6010 15869 6012
rect 15893 6010 15949 6012
rect 15973 6010 16029 6012
rect 16053 6010 16109 6012
rect 15813 5958 15859 6010
rect 15859 5958 15869 6010
rect 15893 5958 15923 6010
rect 15923 5958 15935 6010
rect 15935 5958 15949 6010
rect 15973 5958 15987 6010
rect 15987 5958 15999 6010
rect 15999 5958 16029 6010
rect 16053 5958 16063 6010
rect 16063 5958 16109 6010
rect 15813 5956 15869 5958
rect 15893 5956 15949 5958
rect 15973 5956 16029 5958
rect 16053 5956 16109 5958
rect 15934 5364 15990 5400
rect 15934 5344 15936 5364
rect 15936 5344 15988 5364
rect 15988 5344 15990 5364
rect 15290 5208 15346 5264
rect 15813 4922 15869 4924
rect 15893 4922 15949 4924
rect 15973 4922 16029 4924
rect 16053 4922 16109 4924
rect 15813 4870 15859 4922
rect 15859 4870 15869 4922
rect 15893 4870 15923 4922
rect 15923 4870 15935 4922
rect 15935 4870 15949 4922
rect 15973 4870 15987 4922
rect 15987 4870 15999 4922
rect 15999 4870 16029 4922
rect 16053 4870 16063 4922
rect 16063 4870 16109 4922
rect 15813 4868 15869 4870
rect 15893 4868 15949 4870
rect 15973 4868 16029 4870
rect 16053 4868 16109 4870
rect 15566 4256 15622 4312
rect 15842 4428 15844 4448
rect 15844 4428 15896 4448
rect 15896 4428 15898 4448
rect 15842 4392 15898 4428
rect 15566 4120 15622 4176
rect 15813 3834 15869 3836
rect 15893 3834 15949 3836
rect 15973 3834 16029 3836
rect 16053 3834 16109 3836
rect 15813 3782 15859 3834
rect 15859 3782 15869 3834
rect 15893 3782 15923 3834
rect 15923 3782 15935 3834
rect 15935 3782 15949 3834
rect 15973 3782 15987 3834
rect 15987 3782 15999 3834
rect 15999 3782 16029 3834
rect 16053 3782 16063 3834
rect 16063 3782 16109 3834
rect 15813 3780 15869 3782
rect 15893 3780 15949 3782
rect 15973 3780 16029 3782
rect 16053 3780 16109 3782
rect 15813 2746 15869 2748
rect 15893 2746 15949 2748
rect 15973 2746 16029 2748
rect 16053 2746 16109 2748
rect 15813 2694 15859 2746
rect 15859 2694 15869 2746
rect 15893 2694 15923 2746
rect 15923 2694 15935 2746
rect 15935 2694 15949 2746
rect 15973 2694 15987 2746
rect 15987 2694 15999 2746
rect 15999 2694 16029 2746
rect 16053 2694 16063 2746
rect 16063 2694 16109 2746
rect 15813 2692 15869 2694
rect 15893 2692 15949 2694
rect 15973 2692 16029 2694
rect 16053 2692 16109 2694
rect 15813 1658 15869 1660
rect 15893 1658 15949 1660
rect 15973 1658 16029 1660
rect 16053 1658 16109 1660
rect 15813 1606 15859 1658
rect 15859 1606 15869 1658
rect 15893 1606 15923 1658
rect 15923 1606 15935 1658
rect 15935 1606 15949 1658
rect 15973 1606 15987 1658
rect 15987 1606 15999 1658
rect 15999 1606 16029 1658
rect 16053 1606 16063 1658
rect 16063 1606 16109 1658
rect 15813 1604 15869 1606
rect 15893 1604 15949 1606
rect 15973 1604 16029 1606
rect 16053 1604 16109 1606
rect 16578 3984 16634 4040
rect 17038 9016 17094 9072
rect 17314 8372 17316 8392
rect 17316 8372 17368 8392
rect 17368 8372 17370 8392
rect 17314 8336 17370 8372
rect 16946 8064 17002 8120
rect 16946 4256 17002 4312
rect 17590 9052 17592 9072
rect 17592 9052 17644 9072
rect 17644 9052 17646 9072
rect 17590 9016 17646 9052
rect 18050 9288 18106 9344
rect 17682 8744 17738 8800
rect 18234 7928 18290 7984
rect 17590 6704 17646 6760
rect 8108 570 8164 572
rect 8188 570 8244 572
rect 8268 570 8324 572
rect 8348 570 8404 572
rect 8108 518 8154 570
rect 8154 518 8164 570
rect 8188 518 8218 570
rect 8218 518 8230 570
rect 8230 518 8244 570
rect 8268 518 8282 570
rect 8282 518 8294 570
rect 8294 518 8324 570
rect 8348 518 8358 570
rect 8358 518 8404 570
rect 8108 516 8164 518
rect 8188 516 8244 518
rect 8268 516 8324 518
rect 8348 516 8404 518
rect 15813 570 15869 572
rect 15893 570 15949 572
rect 15973 570 16029 572
rect 16053 570 16109 572
rect 15813 518 15859 570
rect 15859 518 15869 570
rect 15893 518 15923 570
rect 15923 518 15935 570
rect 15935 518 15949 570
rect 15973 518 15987 570
rect 15987 518 15999 570
rect 15999 518 16029 570
rect 16053 518 16063 570
rect 16063 518 16109 570
rect 15813 516 15869 518
rect 15893 516 15949 518
rect 15973 516 16029 518
rect 16053 516 16109 518
rect 17222 3576 17278 3632
rect 17958 6432 18014 6488
rect 17866 6160 17922 6216
rect 18510 9052 18512 9072
rect 18512 9052 18564 9072
rect 18564 9052 18566 9072
rect 18510 9016 18566 9052
rect 18510 8336 18566 8392
rect 18050 4528 18106 4584
rect 19666 18522 19722 18524
rect 19746 18522 19802 18524
rect 19826 18522 19882 18524
rect 19906 18522 19962 18524
rect 19666 18470 19712 18522
rect 19712 18470 19722 18522
rect 19746 18470 19776 18522
rect 19776 18470 19788 18522
rect 19788 18470 19802 18522
rect 19826 18470 19840 18522
rect 19840 18470 19852 18522
rect 19852 18470 19882 18522
rect 19906 18470 19916 18522
rect 19916 18470 19962 18522
rect 19666 18468 19722 18470
rect 19746 18468 19802 18470
rect 19826 18468 19882 18470
rect 19906 18468 19962 18470
rect 19666 17434 19722 17436
rect 19746 17434 19802 17436
rect 19826 17434 19882 17436
rect 19906 17434 19962 17436
rect 19666 17382 19712 17434
rect 19712 17382 19722 17434
rect 19746 17382 19776 17434
rect 19776 17382 19788 17434
rect 19788 17382 19802 17434
rect 19826 17382 19840 17434
rect 19840 17382 19852 17434
rect 19852 17382 19882 17434
rect 19906 17382 19916 17434
rect 19916 17382 19962 17434
rect 19666 17380 19722 17382
rect 19746 17380 19802 17382
rect 19826 17380 19882 17382
rect 19906 17380 19962 17382
rect 19666 16346 19722 16348
rect 19746 16346 19802 16348
rect 19826 16346 19882 16348
rect 19906 16346 19962 16348
rect 19666 16294 19712 16346
rect 19712 16294 19722 16346
rect 19746 16294 19776 16346
rect 19776 16294 19788 16346
rect 19788 16294 19802 16346
rect 19826 16294 19840 16346
rect 19840 16294 19852 16346
rect 19852 16294 19882 16346
rect 19906 16294 19916 16346
rect 19916 16294 19962 16346
rect 19666 16292 19722 16294
rect 19746 16292 19802 16294
rect 19826 16292 19882 16294
rect 19906 16292 19962 16294
rect 19430 14340 19486 14376
rect 19430 14320 19432 14340
rect 19432 14320 19484 14340
rect 19484 14320 19486 14340
rect 19338 13232 19394 13288
rect 18786 12008 18842 12064
rect 18878 11736 18934 11792
rect 19062 11736 19118 11792
rect 18878 10784 18934 10840
rect 18694 9560 18750 9616
rect 19338 11600 19394 11656
rect 19246 9832 19302 9888
rect 19154 8472 19210 8528
rect 18970 7792 19026 7848
rect 18878 6196 18880 6216
rect 18880 6196 18932 6216
rect 18932 6196 18934 6216
rect 18878 6160 18934 6196
rect 19338 5616 19394 5672
rect 18970 4664 19026 4720
rect 19666 15258 19722 15260
rect 19746 15258 19802 15260
rect 19826 15258 19882 15260
rect 19906 15258 19962 15260
rect 19666 15206 19712 15258
rect 19712 15206 19722 15258
rect 19746 15206 19776 15258
rect 19776 15206 19788 15258
rect 19788 15206 19802 15258
rect 19826 15206 19840 15258
rect 19840 15206 19852 15258
rect 19852 15206 19882 15258
rect 19906 15206 19916 15258
rect 19916 15206 19962 15258
rect 19666 15204 19722 15206
rect 19746 15204 19802 15206
rect 19826 15204 19882 15206
rect 19906 15204 19962 15206
rect 19666 14170 19722 14172
rect 19746 14170 19802 14172
rect 19826 14170 19882 14172
rect 19906 14170 19962 14172
rect 19666 14118 19712 14170
rect 19712 14118 19722 14170
rect 19746 14118 19776 14170
rect 19776 14118 19788 14170
rect 19788 14118 19802 14170
rect 19826 14118 19840 14170
rect 19840 14118 19852 14170
rect 19852 14118 19882 14170
rect 19906 14118 19916 14170
rect 19916 14118 19962 14170
rect 19666 14116 19722 14118
rect 19746 14116 19802 14118
rect 19826 14116 19882 14118
rect 19906 14116 19962 14118
rect 19982 13912 20038 13968
rect 19666 13082 19722 13084
rect 19746 13082 19802 13084
rect 19826 13082 19882 13084
rect 19906 13082 19962 13084
rect 19666 13030 19712 13082
rect 19712 13030 19722 13082
rect 19746 13030 19776 13082
rect 19776 13030 19788 13082
rect 19788 13030 19802 13082
rect 19826 13030 19840 13082
rect 19840 13030 19852 13082
rect 19852 13030 19882 13082
rect 19906 13030 19916 13082
rect 19916 13030 19962 13082
rect 19666 13028 19722 13030
rect 19746 13028 19802 13030
rect 19826 13028 19882 13030
rect 19906 13028 19962 13030
rect 19890 12280 19946 12336
rect 19666 11994 19722 11996
rect 19746 11994 19802 11996
rect 19826 11994 19882 11996
rect 19906 11994 19962 11996
rect 19666 11942 19712 11994
rect 19712 11942 19722 11994
rect 19746 11942 19776 11994
rect 19776 11942 19788 11994
rect 19788 11942 19802 11994
rect 19826 11942 19840 11994
rect 19840 11942 19852 11994
rect 19852 11942 19882 11994
rect 19906 11942 19916 11994
rect 19916 11942 19962 11994
rect 19666 11940 19722 11942
rect 19746 11940 19802 11942
rect 19826 11940 19882 11942
rect 19906 11940 19962 11942
rect 19798 11736 19854 11792
rect 19706 11636 19708 11656
rect 19708 11636 19760 11656
rect 19760 11636 19762 11656
rect 19706 11600 19762 11636
rect 19666 10906 19722 10908
rect 19746 10906 19802 10908
rect 19826 10906 19882 10908
rect 19906 10906 19962 10908
rect 19666 10854 19712 10906
rect 19712 10854 19722 10906
rect 19746 10854 19776 10906
rect 19776 10854 19788 10906
rect 19788 10854 19802 10906
rect 19826 10854 19840 10906
rect 19840 10854 19852 10906
rect 19852 10854 19882 10906
rect 19906 10854 19916 10906
rect 19916 10854 19962 10906
rect 19666 10852 19722 10854
rect 19746 10852 19802 10854
rect 19826 10852 19882 10854
rect 19906 10852 19962 10854
rect 19890 10648 19946 10704
rect 19706 10376 19762 10432
rect 19798 10104 19854 10160
rect 20442 14456 20498 14512
rect 20350 13368 20406 13424
rect 20166 12824 20222 12880
rect 20074 11736 20130 11792
rect 20074 11348 20130 11384
rect 20074 11328 20076 11348
rect 20076 11328 20128 11348
rect 20128 11328 20130 11348
rect 19666 9818 19722 9820
rect 19746 9818 19802 9820
rect 19826 9818 19882 9820
rect 19906 9818 19962 9820
rect 19666 9766 19712 9818
rect 19712 9766 19722 9818
rect 19746 9766 19776 9818
rect 19776 9766 19788 9818
rect 19788 9766 19802 9818
rect 19826 9766 19840 9818
rect 19840 9766 19852 9818
rect 19852 9766 19882 9818
rect 19906 9766 19916 9818
rect 19916 9766 19962 9818
rect 19666 9764 19722 9766
rect 19746 9764 19802 9766
rect 19826 9764 19882 9766
rect 19906 9764 19962 9766
rect 19890 9016 19946 9072
rect 19666 8730 19722 8732
rect 19746 8730 19802 8732
rect 19826 8730 19882 8732
rect 19906 8730 19962 8732
rect 19666 8678 19712 8730
rect 19712 8678 19722 8730
rect 19746 8678 19776 8730
rect 19776 8678 19788 8730
rect 19788 8678 19802 8730
rect 19826 8678 19840 8730
rect 19840 8678 19852 8730
rect 19852 8678 19882 8730
rect 19906 8678 19916 8730
rect 19916 8678 19962 8730
rect 19666 8676 19722 8678
rect 19746 8676 19802 8678
rect 19826 8676 19882 8678
rect 19906 8676 19962 8678
rect 19706 7964 19708 7984
rect 19708 7964 19760 7984
rect 19760 7964 19762 7984
rect 19706 7928 19762 7964
rect 19666 7642 19722 7644
rect 19746 7642 19802 7644
rect 19826 7642 19882 7644
rect 19906 7642 19962 7644
rect 19666 7590 19712 7642
rect 19712 7590 19722 7642
rect 19746 7590 19776 7642
rect 19776 7590 19788 7642
rect 19788 7590 19802 7642
rect 19826 7590 19840 7642
rect 19840 7590 19852 7642
rect 19852 7590 19882 7642
rect 19906 7590 19916 7642
rect 19916 7590 19962 7642
rect 19666 7588 19722 7590
rect 19746 7588 19802 7590
rect 19826 7588 19882 7590
rect 19906 7588 19962 7590
rect 19706 6876 19708 6896
rect 19708 6876 19760 6896
rect 19760 6876 19762 6896
rect 19706 6840 19762 6876
rect 19666 6554 19722 6556
rect 19746 6554 19802 6556
rect 19826 6554 19882 6556
rect 19906 6554 19962 6556
rect 19666 6502 19712 6554
rect 19712 6502 19722 6554
rect 19746 6502 19776 6554
rect 19776 6502 19788 6554
rect 19788 6502 19802 6554
rect 19826 6502 19840 6554
rect 19840 6502 19852 6554
rect 19852 6502 19882 6554
rect 19906 6502 19916 6554
rect 19916 6502 19962 6554
rect 19666 6500 19722 6502
rect 19746 6500 19802 6502
rect 19826 6500 19882 6502
rect 19906 6500 19962 6502
rect 19890 5888 19946 5944
rect 19890 5788 19892 5808
rect 19892 5788 19944 5808
rect 19944 5788 19946 5808
rect 19890 5752 19946 5788
rect 19614 5636 19670 5672
rect 19614 5616 19616 5636
rect 19616 5616 19668 5636
rect 19668 5616 19670 5636
rect 19666 5466 19722 5468
rect 19746 5466 19802 5468
rect 19826 5466 19882 5468
rect 19906 5466 19962 5468
rect 19666 5414 19712 5466
rect 19712 5414 19722 5466
rect 19746 5414 19776 5466
rect 19776 5414 19788 5466
rect 19788 5414 19802 5466
rect 19826 5414 19840 5466
rect 19840 5414 19852 5466
rect 19852 5414 19882 5466
rect 19906 5414 19916 5466
rect 19916 5414 19962 5466
rect 19666 5412 19722 5414
rect 19746 5412 19802 5414
rect 19826 5412 19882 5414
rect 19906 5412 19962 5414
rect 19062 4528 19118 4584
rect 18878 4392 18934 4448
rect 19666 4378 19722 4380
rect 19746 4378 19802 4380
rect 19826 4378 19882 4380
rect 19906 4378 19962 4380
rect 19666 4326 19712 4378
rect 19712 4326 19722 4378
rect 19746 4326 19776 4378
rect 19776 4326 19788 4378
rect 19788 4326 19802 4378
rect 19826 4326 19840 4378
rect 19840 4326 19852 4378
rect 19852 4326 19882 4378
rect 19906 4326 19916 4378
rect 19916 4326 19962 4378
rect 19666 4324 19722 4326
rect 19746 4324 19802 4326
rect 19826 4324 19882 4326
rect 19906 4324 19962 4326
rect 20350 12008 20406 12064
rect 23518 19066 23574 19068
rect 23598 19066 23654 19068
rect 23678 19066 23734 19068
rect 23758 19066 23814 19068
rect 23518 19014 23564 19066
rect 23564 19014 23574 19066
rect 23598 19014 23628 19066
rect 23628 19014 23640 19066
rect 23640 19014 23654 19066
rect 23678 19014 23692 19066
rect 23692 19014 23704 19066
rect 23704 19014 23734 19066
rect 23758 19014 23768 19066
rect 23768 19014 23814 19066
rect 23518 19012 23574 19014
rect 23598 19012 23654 19014
rect 23678 19012 23734 19014
rect 23758 19012 23814 19014
rect 31666 19080 31722 19136
rect 31223 19066 31279 19068
rect 31303 19066 31359 19068
rect 31383 19066 31439 19068
rect 31463 19066 31519 19068
rect 31223 19014 31269 19066
rect 31269 19014 31279 19066
rect 31303 19014 31333 19066
rect 31333 19014 31345 19066
rect 31345 19014 31359 19066
rect 31383 19014 31397 19066
rect 31397 19014 31409 19066
rect 31409 19014 31439 19066
rect 31463 19014 31473 19066
rect 31473 19014 31519 19066
rect 31223 19012 31279 19014
rect 31303 19012 31359 19014
rect 31383 19012 31439 19014
rect 31463 19012 31519 19014
rect 23518 17978 23574 17980
rect 23598 17978 23654 17980
rect 23678 17978 23734 17980
rect 23758 17978 23814 17980
rect 23518 17926 23564 17978
rect 23564 17926 23574 17978
rect 23598 17926 23628 17978
rect 23628 17926 23640 17978
rect 23640 17926 23654 17978
rect 23678 17926 23692 17978
rect 23692 17926 23704 17978
rect 23704 17926 23734 17978
rect 23758 17926 23768 17978
rect 23768 17926 23814 17978
rect 23518 17924 23574 17926
rect 23598 17924 23654 17926
rect 23678 17924 23734 17926
rect 23758 17924 23814 17926
rect 20534 9560 20590 9616
rect 20442 9152 20498 9208
rect 20902 14320 20958 14376
rect 21178 13912 21234 13968
rect 20810 11600 20866 11656
rect 20810 11328 20866 11384
rect 21362 13912 21418 13968
rect 21546 13812 21548 13832
rect 21548 13812 21600 13832
rect 21600 13812 21602 13832
rect 21362 13268 21364 13288
rect 21364 13268 21416 13288
rect 21416 13268 21418 13288
rect 21362 13232 21418 13268
rect 21546 13776 21602 13812
rect 22190 13232 22246 13288
rect 21638 12008 21694 12064
rect 21546 10104 21602 10160
rect 21362 9696 21418 9752
rect 20442 8744 20498 8800
rect 20442 8200 20498 8256
rect 20626 8200 20682 8256
rect 20718 5208 20774 5264
rect 22006 11772 22008 11792
rect 22008 11772 22060 11792
rect 22060 11772 22062 11792
rect 22006 11736 22062 11772
rect 22926 14320 22982 14376
rect 22834 13524 22890 13560
rect 22834 13504 22836 13524
rect 22836 13504 22888 13524
rect 22888 13504 22890 13524
rect 22374 9560 22430 9616
rect 23518 16890 23574 16892
rect 23598 16890 23654 16892
rect 23678 16890 23734 16892
rect 23758 16890 23814 16892
rect 23518 16838 23564 16890
rect 23564 16838 23574 16890
rect 23598 16838 23628 16890
rect 23628 16838 23640 16890
rect 23640 16838 23654 16890
rect 23678 16838 23692 16890
rect 23692 16838 23704 16890
rect 23704 16838 23734 16890
rect 23758 16838 23768 16890
rect 23768 16838 23814 16890
rect 23518 16836 23574 16838
rect 23598 16836 23654 16838
rect 23678 16836 23734 16838
rect 23758 16836 23814 16838
rect 23518 15802 23574 15804
rect 23598 15802 23654 15804
rect 23678 15802 23734 15804
rect 23758 15802 23814 15804
rect 23518 15750 23564 15802
rect 23564 15750 23574 15802
rect 23598 15750 23628 15802
rect 23628 15750 23640 15802
rect 23640 15750 23654 15802
rect 23678 15750 23692 15802
rect 23692 15750 23704 15802
rect 23704 15750 23734 15802
rect 23758 15750 23768 15802
rect 23768 15750 23814 15802
rect 23518 15748 23574 15750
rect 23598 15748 23654 15750
rect 23678 15748 23734 15750
rect 23758 15748 23814 15750
rect 23518 14714 23574 14716
rect 23598 14714 23654 14716
rect 23678 14714 23734 14716
rect 23758 14714 23814 14716
rect 23518 14662 23564 14714
rect 23564 14662 23574 14714
rect 23598 14662 23628 14714
rect 23628 14662 23640 14714
rect 23640 14662 23654 14714
rect 23678 14662 23692 14714
rect 23692 14662 23704 14714
rect 23704 14662 23734 14714
rect 23758 14662 23768 14714
rect 23768 14662 23814 14714
rect 23518 14660 23574 14662
rect 23598 14660 23654 14662
rect 23678 14660 23734 14662
rect 23758 14660 23814 14662
rect 23662 14320 23718 14376
rect 23570 13912 23626 13968
rect 23478 13776 23534 13832
rect 23938 14476 23994 14512
rect 27371 18522 27427 18524
rect 27451 18522 27507 18524
rect 27531 18522 27587 18524
rect 27611 18522 27667 18524
rect 27371 18470 27417 18522
rect 27417 18470 27427 18522
rect 27451 18470 27481 18522
rect 27481 18470 27493 18522
rect 27493 18470 27507 18522
rect 27531 18470 27545 18522
rect 27545 18470 27557 18522
rect 27557 18470 27587 18522
rect 27611 18470 27621 18522
rect 27621 18470 27667 18522
rect 27371 18468 27427 18470
rect 27451 18468 27507 18470
rect 27531 18468 27587 18470
rect 27611 18468 27667 18470
rect 31022 18400 31078 18456
rect 31223 17978 31279 17980
rect 31303 17978 31359 17980
rect 31383 17978 31439 17980
rect 31463 17978 31519 17980
rect 31223 17926 31269 17978
rect 31269 17926 31279 17978
rect 31303 17926 31333 17978
rect 31333 17926 31345 17978
rect 31345 17926 31359 17978
rect 31383 17926 31397 17978
rect 31397 17926 31409 17978
rect 31409 17926 31439 17978
rect 31463 17926 31473 17978
rect 31473 17926 31519 17978
rect 31223 17924 31279 17926
rect 31303 17924 31359 17926
rect 31383 17924 31439 17926
rect 31463 17924 31519 17926
rect 27371 17434 27427 17436
rect 27451 17434 27507 17436
rect 27531 17434 27587 17436
rect 27611 17434 27667 17436
rect 27371 17382 27417 17434
rect 27417 17382 27427 17434
rect 27451 17382 27481 17434
rect 27481 17382 27493 17434
rect 27493 17382 27507 17434
rect 27531 17382 27545 17434
rect 27545 17382 27557 17434
rect 27557 17382 27587 17434
rect 27611 17382 27621 17434
rect 27621 17382 27667 17434
rect 27371 17380 27427 17382
rect 27451 17380 27507 17382
rect 27531 17380 27587 17382
rect 27611 17380 27667 17382
rect 23938 14456 23940 14476
rect 23940 14456 23992 14476
rect 23992 14456 23994 14476
rect 23294 13504 23350 13560
rect 23518 13626 23574 13628
rect 23598 13626 23654 13628
rect 23678 13626 23734 13628
rect 23758 13626 23814 13628
rect 23518 13574 23564 13626
rect 23564 13574 23574 13626
rect 23598 13574 23628 13626
rect 23628 13574 23640 13626
rect 23640 13574 23654 13626
rect 23678 13574 23692 13626
rect 23692 13574 23704 13626
rect 23704 13574 23734 13626
rect 23758 13574 23768 13626
rect 23768 13574 23814 13626
rect 23518 13572 23574 13574
rect 23598 13572 23654 13574
rect 23678 13572 23734 13574
rect 23758 13572 23814 13574
rect 23478 13268 23480 13288
rect 23480 13268 23532 13288
rect 23532 13268 23534 13288
rect 23478 13232 23534 13268
rect 22742 11328 22798 11384
rect 23018 11328 23074 11384
rect 23018 10512 23074 10568
rect 19062 3476 19064 3496
rect 19064 3476 19116 3496
rect 19116 3476 19118 3496
rect 19062 3440 19118 3476
rect 19666 3290 19722 3292
rect 19746 3290 19802 3292
rect 19826 3290 19882 3292
rect 19906 3290 19962 3292
rect 19666 3238 19712 3290
rect 19712 3238 19722 3290
rect 19746 3238 19776 3290
rect 19776 3238 19788 3290
rect 19788 3238 19802 3290
rect 19826 3238 19840 3290
rect 19840 3238 19852 3290
rect 19852 3238 19882 3290
rect 19906 3238 19916 3290
rect 19916 3238 19962 3290
rect 19666 3236 19722 3238
rect 19746 3236 19802 3238
rect 19826 3236 19882 3238
rect 19906 3236 19962 3238
rect 19666 2202 19722 2204
rect 19746 2202 19802 2204
rect 19826 2202 19882 2204
rect 19906 2202 19962 2204
rect 19666 2150 19712 2202
rect 19712 2150 19722 2202
rect 19746 2150 19776 2202
rect 19776 2150 19788 2202
rect 19788 2150 19802 2202
rect 19826 2150 19840 2202
rect 19840 2150 19852 2202
rect 19852 2150 19882 2202
rect 19906 2150 19916 2202
rect 19916 2150 19962 2202
rect 19666 2148 19722 2150
rect 19746 2148 19802 2150
rect 19826 2148 19882 2150
rect 19906 2148 19962 2150
rect 19666 1114 19722 1116
rect 19746 1114 19802 1116
rect 19826 1114 19882 1116
rect 19906 1114 19962 1116
rect 19666 1062 19712 1114
rect 19712 1062 19722 1114
rect 19746 1062 19776 1114
rect 19776 1062 19788 1114
rect 19788 1062 19802 1114
rect 19826 1062 19840 1114
rect 19840 1062 19852 1114
rect 19852 1062 19882 1114
rect 19906 1062 19916 1114
rect 19916 1062 19962 1114
rect 19666 1060 19722 1062
rect 19746 1060 19802 1062
rect 19826 1060 19882 1062
rect 19906 1060 19962 1062
rect 20718 3440 20774 3496
rect 22834 6604 22836 6624
rect 22836 6604 22888 6624
rect 22888 6604 22890 6624
rect 22834 6568 22890 6604
rect 22926 5888 22982 5944
rect 23202 11464 23258 11520
rect 23294 10376 23350 10432
rect 23518 12538 23574 12540
rect 23598 12538 23654 12540
rect 23678 12538 23734 12540
rect 23758 12538 23814 12540
rect 23518 12486 23564 12538
rect 23564 12486 23574 12538
rect 23598 12486 23628 12538
rect 23628 12486 23640 12538
rect 23640 12486 23654 12538
rect 23678 12486 23692 12538
rect 23692 12486 23704 12538
rect 23704 12486 23734 12538
rect 23758 12486 23768 12538
rect 23768 12486 23814 12538
rect 23518 12484 23574 12486
rect 23598 12484 23654 12486
rect 23678 12484 23734 12486
rect 23758 12484 23814 12486
rect 24030 11772 24032 11792
rect 24032 11772 24084 11792
rect 24084 11772 24086 11792
rect 24030 11736 24086 11772
rect 23518 11450 23574 11452
rect 23598 11450 23654 11452
rect 23678 11450 23734 11452
rect 23758 11450 23814 11452
rect 23518 11398 23564 11450
rect 23564 11398 23574 11450
rect 23598 11398 23628 11450
rect 23628 11398 23640 11450
rect 23640 11398 23654 11450
rect 23678 11398 23692 11450
rect 23692 11398 23704 11450
rect 23704 11398 23734 11450
rect 23758 11398 23768 11450
rect 23768 11398 23814 11450
rect 23518 11396 23574 11398
rect 23598 11396 23654 11398
rect 23678 11396 23734 11398
rect 23758 11396 23814 11398
rect 23518 10362 23574 10364
rect 23598 10362 23654 10364
rect 23678 10362 23734 10364
rect 23758 10362 23814 10364
rect 23518 10310 23564 10362
rect 23564 10310 23574 10362
rect 23598 10310 23628 10362
rect 23628 10310 23640 10362
rect 23640 10310 23654 10362
rect 23678 10310 23692 10362
rect 23692 10310 23704 10362
rect 23704 10310 23734 10362
rect 23758 10310 23768 10362
rect 23768 10310 23814 10362
rect 23518 10308 23574 10310
rect 23598 10308 23654 10310
rect 23678 10308 23734 10310
rect 23758 10308 23814 10310
rect 23202 9988 23258 10024
rect 23202 9968 23204 9988
rect 23204 9968 23256 9988
rect 23256 9968 23258 9988
rect 23518 9274 23574 9276
rect 23598 9274 23654 9276
rect 23678 9274 23734 9276
rect 23758 9274 23814 9276
rect 23518 9222 23564 9274
rect 23564 9222 23574 9274
rect 23598 9222 23628 9274
rect 23628 9222 23640 9274
rect 23640 9222 23654 9274
rect 23678 9222 23692 9274
rect 23692 9222 23704 9274
rect 23704 9222 23734 9274
rect 23758 9222 23768 9274
rect 23768 9222 23814 9274
rect 23518 9220 23574 9222
rect 23598 9220 23654 9222
rect 23678 9220 23734 9222
rect 23758 9220 23814 9222
rect 23110 8200 23166 8256
rect 23518 8186 23574 8188
rect 23598 8186 23654 8188
rect 23678 8186 23734 8188
rect 23758 8186 23814 8188
rect 23518 8134 23564 8186
rect 23564 8134 23574 8186
rect 23598 8134 23628 8186
rect 23628 8134 23640 8186
rect 23640 8134 23654 8186
rect 23678 8134 23692 8186
rect 23692 8134 23704 8186
rect 23704 8134 23734 8186
rect 23758 8134 23768 8186
rect 23768 8134 23814 8186
rect 23518 8132 23574 8134
rect 23598 8132 23654 8134
rect 23678 8132 23734 8134
rect 23758 8132 23814 8134
rect 23518 7098 23574 7100
rect 23598 7098 23654 7100
rect 23678 7098 23734 7100
rect 23758 7098 23814 7100
rect 23518 7046 23564 7098
rect 23564 7046 23574 7098
rect 23598 7046 23628 7098
rect 23628 7046 23640 7098
rect 23640 7046 23654 7098
rect 23678 7046 23692 7098
rect 23692 7046 23704 7098
rect 23704 7046 23734 7098
rect 23758 7046 23768 7098
rect 23768 7046 23814 7098
rect 23518 7044 23574 7046
rect 23598 7044 23654 7046
rect 23678 7044 23734 7046
rect 23758 7044 23814 7046
rect 23518 6010 23574 6012
rect 23598 6010 23654 6012
rect 23678 6010 23734 6012
rect 23758 6010 23814 6012
rect 23518 5958 23564 6010
rect 23564 5958 23574 6010
rect 23598 5958 23628 6010
rect 23628 5958 23640 6010
rect 23640 5958 23654 6010
rect 23678 5958 23692 6010
rect 23692 5958 23704 6010
rect 23704 5958 23734 6010
rect 23758 5958 23768 6010
rect 23768 5958 23814 6010
rect 23518 5956 23574 5958
rect 23598 5956 23654 5958
rect 23678 5956 23734 5958
rect 23758 5956 23814 5958
rect 22742 5072 22798 5128
rect 21638 4528 21694 4584
rect 23018 4528 23074 4584
rect 22926 4004 22982 4040
rect 22926 3984 22928 4004
rect 22928 3984 22980 4004
rect 22980 3984 22982 4004
rect 23518 4922 23574 4924
rect 23598 4922 23654 4924
rect 23678 4922 23734 4924
rect 23758 4922 23814 4924
rect 23518 4870 23564 4922
rect 23564 4870 23574 4922
rect 23598 4870 23628 4922
rect 23628 4870 23640 4922
rect 23640 4870 23654 4922
rect 23678 4870 23692 4922
rect 23692 4870 23704 4922
rect 23704 4870 23734 4922
rect 23758 4870 23768 4922
rect 23768 4870 23814 4922
rect 23518 4868 23574 4870
rect 23598 4868 23654 4870
rect 23678 4868 23734 4870
rect 23758 4868 23814 4870
rect 23518 3834 23574 3836
rect 23598 3834 23654 3836
rect 23678 3834 23734 3836
rect 23758 3834 23814 3836
rect 23518 3782 23564 3834
rect 23564 3782 23574 3834
rect 23598 3782 23628 3834
rect 23628 3782 23640 3834
rect 23640 3782 23654 3834
rect 23678 3782 23692 3834
rect 23692 3782 23704 3834
rect 23704 3782 23734 3834
rect 23758 3782 23768 3834
rect 23768 3782 23814 3834
rect 23518 3780 23574 3782
rect 23598 3780 23654 3782
rect 23678 3780 23734 3782
rect 23758 3780 23814 3782
rect 23518 2746 23574 2748
rect 23598 2746 23654 2748
rect 23678 2746 23734 2748
rect 23758 2746 23814 2748
rect 23518 2694 23564 2746
rect 23564 2694 23574 2746
rect 23598 2694 23628 2746
rect 23628 2694 23640 2746
rect 23640 2694 23654 2746
rect 23678 2694 23692 2746
rect 23692 2694 23704 2746
rect 23704 2694 23734 2746
rect 23758 2694 23768 2746
rect 23768 2694 23814 2746
rect 23518 2692 23574 2694
rect 23598 2692 23654 2694
rect 23678 2692 23734 2694
rect 23758 2692 23814 2694
rect 23518 1658 23574 1660
rect 23598 1658 23654 1660
rect 23678 1658 23734 1660
rect 23758 1658 23814 1660
rect 23518 1606 23564 1658
rect 23564 1606 23574 1658
rect 23598 1606 23628 1658
rect 23628 1606 23640 1658
rect 23640 1606 23654 1658
rect 23678 1606 23692 1658
rect 23692 1606 23704 1658
rect 23704 1606 23734 1658
rect 23758 1606 23768 1658
rect 23768 1606 23814 1658
rect 23518 1604 23574 1606
rect 23598 1604 23654 1606
rect 23678 1604 23734 1606
rect 23758 1604 23814 1606
rect 24122 9152 24178 9208
rect 24398 12144 24454 12200
rect 24582 11736 24638 11792
rect 25318 12280 25374 12336
rect 24490 9016 24546 9072
rect 25686 9580 25742 9616
rect 25686 9560 25688 9580
rect 25688 9560 25740 9580
rect 25740 9560 25742 9580
rect 27371 16346 27427 16348
rect 27451 16346 27507 16348
rect 27531 16346 27587 16348
rect 27611 16346 27667 16348
rect 27371 16294 27417 16346
rect 27417 16294 27427 16346
rect 27451 16294 27481 16346
rect 27481 16294 27493 16346
rect 27493 16294 27507 16346
rect 27531 16294 27545 16346
rect 27545 16294 27557 16346
rect 27557 16294 27587 16346
rect 27611 16294 27621 16346
rect 27621 16294 27667 16346
rect 27371 16292 27427 16294
rect 27451 16292 27507 16294
rect 27531 16292 27587 16294
rect 27611 16292 27667 16294
rect 27371 15258 27427 15260
rect 27451 15258 27507 15260
rect 27531 15258 27587 15260
rect 27611 15258 27667 15260
rect 27371 15206 27417 15258
rect 27417 15206 27427 15258
rect 27451 15206 27481 15258
rect 27481 15206 27493 15258
rect 27493 15206 27507 15258
rect 27531 15206 27545 15258
rect 27545 15206 27557 15258
rect 27557 15206 27587 15258
rect 27611 15206 27621 15258
rect 27621 15206 27667 15258
rect 27371 15204 27427 15206
rect 27451 15204 27507 15206
rect 27531 15204 27587 15206
rect 27611 15204 27667 15206
rect 27371 14170 27427 14172
rect 27451 14170 27507 14172
rect 27531 14170 27587 14172
rect 27611 14170 27667 14172
rect 27371 14118 27417 14170
rect 27417 14118 27427 14170
rect 27451 14118 27481 14170
rect 27481 14118 27493 14170
rect 27493 14118 27507 14170
rect 27531 14118 27545 14170
rect 27545 14118 27557 14170
rect 27557 14118 27587 14170
rect 27611 14118 27621 14170
rect 27621 14118 27667 14170
rect 27371 14116 27427 14118
rect 27451 14116 27507 14118
rect 27531 14116 27587 14118
rect 27611 14116 27667 14118
rect 27371 13082 27427 13084
rect 27451 13082 27507 13084
rect 27531 13082 27587 13084
rect 27611 13082 27667 13084
rect 27371 13030 27417 13082
rect 27417 13030 27427 13082
rect 27451 13030 27481 13082
rect 27481 13030 27493 13082
rect 27493 13030 27507 13082
rect 27531 13030 27545 13082
rect 27545 13030 27557 13082
rect 27557 13030 27587 13082
rect 27611 13030 27621 13082
rect 27621 13030 27667 13082
rect 27371 13028 27427 13030
rect 27451 13028 27507 13030
rect 27531 13028 27587 13030
rect 27611 13028 27667 13030
rect 27371 11994 27427 11996
rect 27451 11994 27507 11996
rect 27531 11994 27587 11996
rect 27611 11994 27667 11996
rect 27371 11942 27417 11994
rect 27417 11942 27427 11994
rect 27451 11942 27481 11994
rect 27481 11942 27493 11994
rect 27493 11942 27507 11994
rect 27531 11942 27545 11994
rect 27545 11942 27557 11994
rect 27557 11942 27587 11994
rect 27611 11942 27621 11994
rect 27621 11942 27667 11994
rect 27371 11940 27427 11942
rect 27451 11940 27507 11942
rect 27531 11940 27587 11942
rect 27611 11940 27667 11942
rect 27710 11192 27766 11248
rect 27371 10906 27427 10908
rect 27451 10906 27507 10908
rect 27531 10906 27587 10908
rect 27611 10906 27667 10908
rect 27371 10854 27417 10906
rect 27417 10854 27427 10906
rect 27451 10854 27481 10906
rect 27481 10854 27493 10906
rect 27493 10854 27507 10906
rect 27531 10854 27545 10906
rect 27545 10854 27557 10906
rect 27557 10854 27587 10906
rect 27611 10854 27621 10906
rect 27621 10854 27667 10906
rect 27371 10852 27427 10854
rect 27451 10852 27507 10854
rect 27531 10852 27587 10854
rect 27611 10852 27667 10854
rect 26330 9424 26386 9480
rect 26882 10104 26938 10160
rect 27371 9818 27427 9820
rect 27451 9818 27507 9820
rect 27531 9818 27587 9820
rect 27611 9818 27667 9820
rect 27371 9766 27417 9818
rect 27417 9766 27427 9818
rect 27451 9766 27481 9818
rect 27481 9766 27493 9818
rect 27493 9766 27507 9818
rect 27531 9766 27545 9818
rect 27545 9766 27557 9818
rect 27557 9766 27587 9818
rect 27611 9766 27621 9818
rect 27621 9766 27667 9818
rect 27371 9764 27427 9766
rect 27451 9764 27507 9766
rect 27531 9764 27587 9766
rect 27611 9764 27667 9766
rect 24766 8880 24822 8936
rect 24858 8744 24914 8800
rect 27371 8730 27427 8732
rect 27451 8730 27507 8732
rect 27531 8730 27587 8732
rect 27611 8730 27667 8732
rect 27371 8678 27417 8730
rect 27417 8678 27427 8730
rect 27451 8678 27481 8730
rect 27481 8678 27493 8730
rect 27493 8678 27507 8730
rect 27531 8678 27545 8730
rect 27545 8678 27557 8730
rect 27557 8678 27587 8730
rect 27611 8678 27621 8730
rect 27621 8678 27667 8730
rect 27371 8676 27427 8678
rect 27451 8676 27507 8678
rect 27531 8676 27587 8678
rect 27611 8676 27667 8678
rect 26698 7812 26754 7848
rect 26698 7792 26700 7812
rect 26700 7792 26752 7812
rect 26752 7792 26754 7812
rect 27371 7642 27427 7644
rect 27451 7642 27507 7644
rect 27531 7642 27587 7644
rect 27611 7642 27667 7644
rect 27371 7590 27417 7642
rect 27417 7590 27427 7642
rect 27451 7590 27481 7642
rect 27481 7590 27493 7642
rect 27493 7590 27507 7642
rect 27531 7590 27545 7642
rect 27545 7590 27557 7642
rect 27557 7590 27587 7642
rect 27611 7590 27621 7642
rect 27621 7590 27667 7642
rect 27371 7588 27427 7590
rect 27451 7588 27507 7590
rect 27531 7588 27587 7590
rect 27611 7588 27667 7590
rect 27371 6554 27427 6556
rect 27451 6554 27507 6556
rect 27531 6554 27587 6556
rect 27611 6554 27667 6556
rect 27371 6502 27417 6554
rect 27417 6502 27427 6554
rect 27451 6502 27481 6554
rect 27481 6502 27493 6554
rect 27493 6502 27507 6554
rect 27531 6502 27545 6554
rect 27545 6502 27557 6554
rect 27557 6502 27587 6554
rect 27611 6502 27621 6554
rect 27621 6502 27667 6554
rect 27371 6500 27427 6502
rect 27451 6500 27507 6502
rect 27531 6500 27587 6502
rect 27611 6500 27667 6502
rect 27371 5466 27427 5468
rect 27451 5466 27507 5468
rect 27531 5466 27587 5468
rect 27611 5466 27667 5468
rect 27371 5414 27417 5466
rect 27417 5414 27427 5466
rect 27451 5414 27481 5466
rect 27481 5414 27493 5466
rect 27493 5414 27507 5466
rect 27531 5414 27545 5466
rect 27545 5414 27557 5466
rect 27557 5414 27587 5466
rect 27611 5414 27621 5466
rect 27621 5414 27667 5466
rect 27371 5412 27427 5414
rect 27451 5412 27507 5414
rect 27531 5412 27587 5414
rect 27611 5412 27667 5414
rect 27371 4378 27427 4380
rect 27451 4378 27507 4380
rect 27531 4378 27587 4380
rect 27611 4378 27667 4380
rect 27371 4326 27417 4378
rect 27417 4326 27427 4378
rect 27451 4326 27481 4378
rect 27481 4326 27493 4378
rect 27493 4326 27507 4378
rect 27531 4326 27545 4378
rect 27545 4326 27557 4378
rect 27557 4326 27587 4378
rect 27611 4326 27621 4378
rect 27621 4326 27667 4378
rect 27371 4324 27427 4326
rect 27451 4324 27507 4326
rect 27531 4324 27587 4326
rect 27611 4324 27667 4326
rect 26606 3984 26662 4040
rect 31223 16890 31279 16892
rect 31303 16890 31359 16892
rect 31383 16890 31439 16892
rect 31463 16890 31519 16892
rect 31223 16838 31269 16890
rect 31269 16838 31279 16890
rect 31303 16838 31333 16890
rect 31333 16838 31345 16890
rect 31345 16838 31359 16890
rect 31383 16838 31397 16890
rect 31397 16838 31409 16890
rect 31409 16838 31439 16890
rect 31463 16838 31473 16890
rect 31473 16838 31519 16890
rect 31223 16836 31279 16838
rect 31303 16836 31359 16838
rect 31383 16836 31439 16838
rect 31463 16836 31519 16838
rect 31223 15802 31279 15804
rect 31303 15802 31359 15804
rect 31383 15802 31439 15804
rect 31463 15802 31519 15804
rect 31223 15750 31269 15802
rect 31269 15750 31279 15802
rect 31303 15750 31333 15802
rect 31333 15750 31345 15802
rect 31345 15750 31359 15802
rect 31383 15750 31397 15802
rect 31397 15750 31409 15802
rect 31409 15750 31439 15802
rect 31463 15750 31473 15802
rect 31473 15750 31519 15802
rect 31223 15748 31279 15750
rect 31303 15748 31359 15750
rect 31383 15748 31439 15750
rect 31463 15748 31519 15750
rect 28906 14320 28962 14376
rect 31223 14714 31279 14716
rect 31303 14714 31359 14716
rect 31383 14714 31439 14716
rect 31463 14714 31519 14716
rect 31223 14662 31269 14714
rect 31269 14662 31279 14714
rect 31303 14662 31333 14714
rect 31333 14662 31345 14714
rect 31345 14662 31359 14714
rect 31383 14662 31397 14714
rect 31397 14662 31409 14714
rect 31409 14662 31439 14714
rect 31463 14662 31473 14714
rect 31473 14662 31519 14714
rect 31223 14660 31279 14662
rect 31303 14660 31359 14662
rect 31383 14660 31439 14662
rect 31463 14660 31519 14662
rect 28630 12280 28686 12336
rect 31223 13626 31279 13628
rect 31303 13626 31359 13628
rect 31383 13626 31439 13628
rect 31463 13626 31519 13628
rect 31223 13574 31269 13626
rect 31269 13574 31279 13626
rect 31303 13574 31333 13626
rect 31333 13574 31345 13626
rect 31345 13574 31359 13626
rect 31383 13574 31397 13626
rect 31397 13574 31409 13626
rect 31409 13574 31439 13626
rect 31463 13574 31473 13626
rect 31473 13574 31519 13626
rect 31223 13572 31279 13574
rect 31303 13572 31359 13574
rect 31383 13572 31439 13574
rect 31463 13572 31519 13574
rect 30746 13368 30802 13424
rect 31223 12538 31279 12540
rect 31303 12538 31359 12540
rect 31383 12538 31439 12540
rect 31463 12538 31519 12540
rect 31223 12486 31269 12538
rect 31269 12486 31279 12538
rect 31303 12486 31333 12538
rect 31333 12486 31345 12538
rect 31345 12486 31359 12538
rect 31383 12486 31397 12538
rect 31397 12486 31409 12538
rect 31409 12486 31439 12538
rect 31463 12486 31473 12538
rect 31473 12486 31519 12538
rect 31223 12484 31279 12486
rect 31303 12484 31359 12486
rect 31383 12484 31439 12486
rect 31463 12484 31519 12486
rect 31223 11450 31279 11452
rect 31303 11450 31359 11452
rect 31383 11450 31439 11452
rect 31463 11450 31519 11452
rect 31223 11398 31269 11450
rect 31269 11398 31279 11450
rect 31303 11398 31333 11450
rect 31333 11398 31345 11450
rect 31345 11398 31359 11450
rect 31383 11398 31397 11450
rect 31397 11398 31409 11450
rect 31409 11398 31439 11450
rect 31463 11398 31473 11450
rect 31473 11398 31519 11450
rect 31223 11396 31279 11398
rect 31303 11396 31359 11398
rect 31383 11396 31439 11398
rect 31463 11396 31519 11398
rect 31223 10362 31279 10364
rect 31303 10362 31359 10364
rect 31383 10362 31439 10364
rect 31463 10362 31519 10364
rect 31223 10310 31269 10362
rect 31269 10310 31279 10362
rect 31303 10310 31333 10362
rect 31333 10310 31345 10362
rect 31345 10310 31359 10362
rect 31383 10310 31397 10362
rect 31397 10310 31409 10362
rect 31409 10310 31439 10362
rect 31463 10310 31473 10362
rect 31473 10310 31519 10362
rect 31223 10308 31279 10310
rect 31303 10308 31359 10310
rect 31383 10308 31439 10310
rect 31463 10308 31519 10310
rect 31666 10240 31722 10296
rect 31223 9274 31279 9276
rect 31303 9274 31359 9276
rect 31383 9274 31439 9276
rect 31463 9274 31519 9276
rect 31223 9222 31269 9274
rect 31269 9222 31279 9274
rect 31303 9222 31333 9274
rect 31333 9222 31345 9274
rect 31345 9222 31359 9274
rect 31383 9222 31397 9274
rect 31397 9222 31409 9274
rect 31409 9222 31439 9274
rect 31463 9222 31473 9274
rect 31473 9222 31519 9274
rect 31223 9220 31279 9222
rect 31303 9220 31359 9222
rect 31383 9220 31439 9222
rect 31463 9220 31519 9222
rect 30930 9172 30986 9208
rect 30930 9152 30932 9172
rect 30932 9152 30984 9172
rect 30984 9152 30986 9172
rect 31223 8186 31279 8188
rect 31303 8186 31359 8188
rect 31383 8186 31439 8188
rect 31463 8186 31519 8188
rect 31223 8134 31269 8186
rect 31269 8134 31279 8186
rect 31303 8134 31333 8186
rect 31333 8134 31345 8186
rect 31345 8134 31359 8186
rect 31383 8134 31397 8186
rect 31397 8134 31409 8186
rect 31409 8134 31439 8186
rect 31463 8134 31473 8186
rect 31473 8134 31519 8186
rect 31223 8132 31279 8134
rect 31303 8132 31359 8134
rect 31383 8132 31439 8134
rect 31463 8132 31519 8134
rect 30930 7928 30986 7984
rect 31223 7098 31279 7100
rect 31303 7098 31359 7100
rect 31383 7098 31439 7100
rect 31463 7098 31519 7100
rect 31223 7046 31269 7098
rect 31269 7046 31279 7098
rect 31303 7046 31333 7098
rect 31333 7046 31345 7098
rect 31345 7046 31359 7098
rect 31383 7046 31397 7098
rect 31397 7046 31409 7098
rect 31409 7046 31439 7098
rect 31463 7046 31473 7098
rect 31473 7046 31519 7098
rect 31223 7044 31279 7046
rect 31303 7044 31359 7046
rect 31383 7044 31439 7046
rect 31463 7044 31519 7046
rect 31022 6840 31078 6896
rect 29366 5636 29422 5672
rect 29366 5616 29368 5636
rect 29368 5616 29420 5636
rect 29420 5616 29422 5636
rect 31223 6010 31279 6012
rect 31303 6010 31359 6012
rect 31383 6010 31439 6012
rect 31463 6010 31519 6012
rect 31223 5958 31269 6010
rect 31269 5958 31279 6010
rect 31303 5958 31333 6010
rect 31333 5958 31345 6010
rect 31345 5958 31359 6010
rect 31383 5958 31397 6010
rect 31397 5958 31409 6010
rect 31409 5958 31439 6010
rect 31463 5958 31473 6010
rect 31473 5958 31519 6010
rect 31223 5956 31279 5958
rect 31303 5956 31359 5958
rect 31383 5956 31439 5958
rect 31463 5956 31519 5958
rect 31223 4922 31279 4924
rect 31303 4922 31359 4924
rect 31383 4922 31439 4924
rect 31463 4922 31519 4924
rect 31223 4870 31269 4922
rect 31269 4870 31279 4922
rect 31303 4870 31333 4922
rect 31333 4870 31345 4922
rect 31345 4870 31359 4922
rect 31383 4870 31397 4922
rect 31397 4870 31409 4922
rect 31409 4870 31439 4922
rect 31463 4870 31473 4922
rect 31473 4870 31519 4922
rect 31223 4868 31279 4870
rect 31303 4868 31359 4870
rect 31383 4868 31439 4870
rect 31463 4868 31519 4870
rect 27371 3290 27427 3292
rect 27451 3290 27507 3292
rect 27531 3290 27587 3292
rect 27611 3290 27667 3292
rect 27371 3238 27417 3290
rect 27417 3238 27427 3290
rect 27451 3238 27481 3290
rect 27481 3238 27493 3290
rect 27493 3238 27507 3290
rect 27531 3238 27545 3290
rect 27545 3238 27557 3290
rect 27557 3238 27587 3290
rect 27611 3238 27621 3290
rect 27621 3238 27667 3290
rect 27371 3236 27427 3238
rect 27451 3236 27507 3238
rect 27531 3236 27587 3238
rect 27611 3236 27667 3238
rect 31223 3834 31279 3836
rect 31303 3834 31359 3836
rect 31383 3834 31439 3836
rect 31463 3834 31519 3836
rect 31223 3782 31269 3834
rect 31269 3782 31279 3834
rect 31303 3782 31333 3834
rect 31333 3782 31345 3834
rect 31345 3782 31359 3834
rect 31383 3782 31397 3834
rect 31397 3782 31409 3834
rect 31409 3782 31439 3834
rect 31463 3782 31473 3834
rect 31473 3782 31519 3834
rect 31223 3780 31279 3782
rect 31303 3780 31359 3782
rect 31383 3780 31439 3782
rect 31463 3780 31519 3782
rect 31666 2760 31722 2816
rect 31223 2746 31279 2748
rect 31303 2746 31359 2748
rect 31383 2746 31439 2748
rect 31463 2746 31519 2748
rect 31223 2694 31269 2746
rect 31269 2694 31279 2746
rect 31303 2694 31333 2746
rect 31333 2694 31345 2746
rect 31345 2694 31359 2746
rect 31383 2694 31397 2746
rect 31397 2694 31409 2746
rect 31409 2694 31439 2746
rect 31463 2694 31473 2746
rect 31473 2694 31519 2746
rect 31223 2692 31279 2694
rect 31303 2692 31359 2694
rect 31383 2692 31439 2694
rect 31463 2692 31519 2694
rect 27371 2202 27427 2204
rect 27451 2202 27507 2204
rect 27531 2202 27587 2204
rect 27611 2202 27667 2204
rect 27371 2150 27417 2202
rect 27417 2150 27427 2202
rect 27451 2150 27481 2202
rect 27481 2150 27493 2202
rect 27493 2150 27507 2202
rect 27531 2150 27545 2202
rect 27545 2150 27557 2202
rect 27557 2150 27587 2202
rect 27611 2150 27621 2202
rect 27621 2150 27667 2202
rect 27371 2148 27427 2150
rect 27451 2148 27507 2150
rect 27531 2148 27587 2150
rect 27611 2148 27667 2150
rect 31022 2080 31078 2136
rect 31223 1658 31279 1660
rect 31303 1658 31359 1660
rect 31383 1658 31439 1660
rect 31463 1658 31519 1660
rect 31223 1606 31269 1658
rect 31269 1606 31279 1658
rect 31303 1606 31333 1658
rect 31333 1606 31345 1658
rect 31345 1606 31359 1658
rect 31383 1606 31397 1658
rect 31397 1606 31409 1658
rect 31409 1606 31439 1658
rect 31463 1606 31473 1658
rect 31473 1606 31519 1658
rect 31223 1604 31279 1606
rect 31303 1604 31359 1606
rect 31383 1604 31439 1606
rect 31463 1604 31519 1606
rect 31022 1400 31078 1456
rect 27371 1114 27427 1116
rect 27451 1114 27507 1116
rect 27531 1114 27587 1116
rect 27611 1114 27667 1116
rect 27371 1062 27417 1114
rect 27417 1062 27427 1114
rect 27451 1062 27481 1114
rect 27481 1062 27493 1114
rect 27493 1062 27507 1114
rect 27531 1062 27545 1114
rect 27545 1062 27557 1114
rect 27557 1062 27587 1114
rect 27611 1062 27621 1114
rect 27621 1062 27667 1114
rect 27371 1060 27427 1062
rect 27451 1060 27507 1062
rect 27531 1060 27587 1062
rect 27611 1060 27667 1062
rect 31022 756 31024 776
rect 31024 756 31076 776
rect 31076 756 31078 776
rect 31022 720 31078 756
rect 23518 570 23574 572
rect 23598 570 23654 572
rect 23678 570 23734 572
rect 23758 570 23814 572
rect 23518 518 23564 570
rect 23564 518 23574 570
rect 23598 518 23628 570
rect 23628 518 23640 570
rect 23640 518 23654 570
rect 23678 518 23692 570
rect 23692 518 23704 570
rect 23704 518 23734 570
rect 23758 518 23768 570
rect 23768 518 23814 570
rect 23518 516 23574 518
rect 23598 516 23654 518
rect 23678 516 23734 518
rect 23758 516 23814 518
rect 31223 570 31279 572
rect 31303 570 31359 572
rect 31383 570 31439 572
rect 31463 570 31519 572
rect 31223 518 31269 570
rect 31269 518 31279 570
rect 31303 518 31333 570
rect 31333 518 31345 570
rect 31345 518 31359 570
rect 31383 518 31397 570
rect 31397 518 31409 570
rect 31409 518 31439 570
rect 31463 518 31473 570
rect 31473 518 31519 570
rect 31223 516 31279 518
rect 31303 516 31359 518
rect 31383 516 31439 518
rect 31463 516 31519 518
<< metal3 >>
rect 0 19818 400 19848
rect 1117 19818 1183 19821
rect 0 19816 1183 19818
rect 0 19760 1122 19816
rect 1178 19760 1183 19816
rect 0 19758 1183 19760
rect 0 19728 400 19758
rect 1117 19755 1183 19758
rect 0 19138 400 19168
rect 749 19138 815 19141
rect 0 19136 815 19138
rect 0 19080 754 19136
rect 810 19080 815 19136
rect 0 19078 815 19080
rect 0 19048 400 19078
rect 749 19075 815 19078
rect 31600 19136 32000 19168
rect 31600 19080 31666 19136
rect 31722 19080 32000 19136
rect 8098 19072 8414 19073
rect 8098 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8414 19072
rect 8098 19007 8414 19008
rect 15803 19072 16119 19073
rect 15803 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16119 19072
rect 15803 19007 16119 19008
rect 23508 19072 23824 19073
rect 23508 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23824 19072
rect 23508 19007 23824 19008
rect 31213 19072 31529 19073
rect 31213 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31529 19072
rect 31600 19048 32000 19080
rect 31213 19007 31529 19008
rect 4246 18528 4562 18529
rect 0 18458 400 18488
rect 4246 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4562 18528
rect 4246 18463 4562 18464
rect 11951 18528 12267 18529
rect 11951 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12267 18528
rect 11951 18463 12267 18464
rect 19656 18528 19972 18529
rect 19656 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19972 18528
rect 19656 18463 19972 18464
rect 27361 18528 27677 18529
rect 27361 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27677 18528
rect 27361 18463 27677 18464
rect 841 18458 907 18461
rect 0 18456 907 18458
rect 0 18400 846 18456
rect 902 18400 907 18456
rect 0 18398 907 18400
rect 0 18368 400 18398
rect 841 18395 907 18398
rect 31017 18458 31083 18461
rect 31600 18458 32000 18488
rect 31017 18456 32000 18458
rect 31017 18400 31022 18456
rect 31078 18400 32000 18456
rect 31017 18398 32000 18400
rect 31017 18395 31083 18398
rect 31600 18368 32000 18398
rect 15009 18052 15075 18053
rect 14958 18050 14964 18052
rect 14918 17990 14964 18050
rect 15028 18048 15075 18052
rect 15070 17992 15075 18048
rect 14958 17988 14964 17990
rect 15028 17988 15075 17992
rect 15009 17987 15075 17988
rect 8098 17984 8414 17985
rect 8098 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8414 17984
rect 8098 17919 8414 17920
rect 15803 17984 16119 17985
rect 15803 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16119 17984
rect 15803 17919 16119 17920
rect 23508 17984 23824 17985
rect 23508 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23824 17984
rect 23508 17919 23824 17920
rect 31213 17984 31529 17985
rect 31213 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31529 17984
rect 31213 17919 31529 17920
rect 0 17778 400 17808
rect 841 17778 907 17781
rect 0 17776 907 17778
rect 0 17720 846 17776
rect 902 17720 907 17776
rect 0 17718 907 17720
rect 0 17688 400 17718
rect 841 17715 907 17718
rect 4246 17440 4562 17441
rect 4246 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4562 17440
rect 4246 17375 4562 17376
rect 11951 17440 12267 17441
rect 11951 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12267 17440
rect 11951 17375 12267 17376
rect 19656 17440 19972 17441
rect 19656 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19972 17440
rect 19656 17375 19972 17376
rect 27361 17440 27677 17441
rect 27361 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27677 17440
rect 27361 17375 27677 17376
rect 0 17098 400 17128
rect 841 17098 907 17101
rect 0 17096 907 17098
rect 0 17040 846 17096
rect 902 17040 907 17096
rect 0 17038 907 17040
rect 0 17008 400 17038
rect 841 17035 907 17038
rect 8098 16896 8414 16897
rect 8098 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8414 16896
rect 8098 16831 8414 16832
rect 15803 16896 16119 16897
rect 15803 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16119 16896
rect 15803 16831 16119 16832
rect 23508 16896 23824 16897
rect 23508 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23824 16896
rect 23508 16831 23824 16832
rect 31213 16896 31529 16897
rect 31213 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31529 16896
rect 31213 16831 31529 16832
rect 17769 16690 17835 16693
rect 18822 16690 18828 16692
rect 17769 16688 18828 16690
rect 17769 16632 17774 16688
rect 17830 16632 18828 16688
rect 17769 16630 18828 16632
rect 17769 16627 17835 16630
rect 18822 16628 18828 16630
rect 18892 16628 18898 16692
rect 4246 16352 4562 16353
rect 4246 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4562 16352
rect 4246 16287 4562 16288
rect 11951 16352 12267 16353
rect 11951 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12267 16352
rect 11951 16287 12267 16288
rect 19656 16352 19972 16353
rect 19656 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19972 16352
rect 19656 16287 19972 16288
rect 27361 16352 27677 16353
rect 27361 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27677 16352
rect 27361 16287 27677 16288
rect 16021 16010 16087 16013
rect 16614 16010 16620 16012
rect 16021 16008 16620 16010
rect 16021 15952 16026 16008
rect 16082 15952 16620 16008
rect 16021 15950 16620 15952
rect 16021 15947 16087 15950
rect 16614 15948 16620 15950
rect 16684 15948 16690 16012
rect 8098 15808 8414 15809
rect 8098 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8414 15808
rect 8098 15743 8414 15744
rect 15803 15808 16119 15809
rect 15803 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16119 15808
rect 15803 15743 16119 15744
rect 23508 15808 23824 15809
rect 23508 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23824 15808
rect 23508 15743 23824 15744
rect 31213 15808 31529 15809
rect 31213 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31529 15808
rect 31213 15743 31529 15744
rect 4246 15264 4562 15265
rect 4246 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4562 15264
rect 4246 15199 4562 15200
rect 11951 15264 12267 15265
rect 11951 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12267 15264
rect 11951 15199 12267 15200
rect 19656 15264 19972 15265
rect 19656 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19972 15264
rect 19656 15199 19972 15200
rect 27361 15264 27677 15265
rect 27361 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27677 15264
rect 27361 15199 27677 15200
rect 8201 15058 8267 15061
rect 17677 15058 17743 15061
rect 8201 15056 17743 15058
rect 8201 15000 8206 15056
rect 8262 15000 17682 15056
rect 17738 15000 17743 15056
rect 8201 14998 17743 15000
rect 8201 14995 8267 14998
rect 17677 14995 17743 14998
rect 5993 14922 6059 14925
rect 18689 14922 18755 14925
rect 5993 14920 18755 14922
rect 5993 14864 5998 14920
rect 6054 14864 18694 14920
rect 18750 14864 18755 14920
rect 5993 14862 18755 14864
rect 5993 14859 6059 14862
rect 18689 14859 18755 14862
rect 8098 14720 8414 14721
rect 8098 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8414 14720
rect 8098 14655 8414 14656
rect 15803 14720 16119 14721
rect 15803 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16119 14720
rect 15803 14655 16119 14656
rect 23508 14720 23824 14721
rect 23508 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23824 14720
rect 23508 14655 23824 14656
rect 31213 14720 31529 14721
rect 31213 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31529 14720
rect 31213 14655 31529 14656
rect 16982 14588 16988 14652
rect 17052 14650 17058 14652
rect 17861 14650 17927 14653
rect 17052 14648 17927 14650
rect 17052 14592 17866 14648
rect 17922 14592 17927 14648
rect 17052 14590 17927 14592
rect 17052 14588 17058 14590
rect 17861 14587 17927 14590
rect 15009 14514 15075 14517
rect 18873 14514 18939 14517
rect 15009 14512 18939 14514
rect 15009 14456 15014 14512
rect 15070 14456 18878 14512
rect 18934 14456 18939 14512
rect 15009 14454 18939 14456
rect 15009 14451 15075 14454
rect 18873 14451 18939 14454
rect 20437 14514 20503 14517
rect 23933 14514 23999 14517
rect 20437 14512 23999 14514
rect 20437 14456 20442 14512
rect 20498 14456 23938 14512
rect 23994 14456 23999 14512
rect 20437 14454 23999 14456
rect 20437 14451 20503 14454
rect 23933 14451 23999 14454
rect 19425 14378 19491 14381
rect 20897 14378 20963 14381
rect 22921 14378 22987 14381
rect 19425 14376 22987 14378
rect 19425 14320 19430 14376
rect 19486 14320 20902 14376
rect 20958 14320 22926 14376
rect 22982 14320 22987 14376
rect 19425 14318 22987 14320
rect 19425 14315 19491 14318
rect 20897 14315 20963 14318
rect 22921 14315 22987 14318
rect 23657 14378 23723 14381
rect 28901 14378 28967 14381
rect 23657 14376 28967 14378
rect 23657 14320 23662 14376
rect 23718 14320 28906 14376
rect 28962 14320 28967 14376
rect 23657 14318 28967 14320
rect 23657 14315 23723 14318
rect 28901 14315 28967 14318
rect 4246 14176 4562 14177
rect 4246 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4562 14176
rect 4246 14111 4562 14112
rect 11951 14176 12267 14177
rect 11951 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12267 14176
rect 11951 14111 12267 14112
rect 19656 14176 19972 14177
rect 19656 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19972 14176
rect 19656 14111 19972 14112
rect 27361 14176 27677 14177
rect 27361 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27677 14176
rect 27361 14111 27677 14112
rect 19977 13970 20043 13973
rect 21173 13970 21239 13973
rect 19977 13968 21239 13970
rect 19977 13912 19982 13968
rect 20038 13912 21178 13968
rect 21234 13912 21239 13968
rect 19977 13910 21239 13912
rect 19977 13907 20043 13910
rect 21173 13907 21239 13910
rect 21357 13970 21423 13973
rect 23565 13970 23631 13973
rect 21357 13968 23631 13970
rect 21357 13912 21362 13968
rect 21418 13912 23570 13968
rect 23626 13912 23631 13968
rect 21357 13910 23631 13912
rect 21357 13907 21423 13910
rect 23565 13907 23631 13910
rect 16757 13836 16823 13837
rect 15518 13774 16314 13834
rect 11237 13698 11303 13701
rect 13905 13698 13971 13701
rect 11237 13696 13971 13698
rect 11237 13640 11242 13696
rect 11298 13640 13910 13696
rect 13966 13640 13971 13696
rect 11237 13638 13971 13640
rect 11237 13635 11303 13638
rect 13905 13635 13971 13638
rect 8098 13632 8414 13633
rect 8098 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8414 13632
rect 8098 13567 8414 13568
rect 11789 13562 11855 13565
rect 15518 13562 15578 13774
rect 16254 13698 16314 13774
rect 16757 13832 16804 13836
rect 16868 13834 16874 13836
rect 21541 13834 21607 13837
rect 23473 13834 23539 13837
rect 16757 13776 16762 13832
rect 16757 13772 16804 13776
rect 16868 13774 16914 13834
rect 21541 13832 23539 13834
rect 21541 13776 21546 13832
rect 21602 13776 23478 13832
rect 23534 13776 23539 13832
rect 21541 13774 23539 13776
rect 16868 13772 16874 13774
rect 16757 13771 16823 13772
rect 21541 13771 21607 13774
rect 23473 13771 23539 13774
rect 18689 13698 18755 13701
rect 16254 13696 18755 13698
rect 16254 13640 18694 13696
rect 18750 13640 18755 13696
rect 16254 13638 18755 13640
rect 18689 13635 18755 13638
rect 15803 13632 16119 13633
rect 15803 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16119 13632
rect 15803 13567 16119 13568
rect 23508 13632 23824 13633
rect 23508 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23824 13632
rect 23508 13567 23824 13568
rect 31213 13632 31529 13633
rect 31213 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31529 13632
rect 31213 13567 31529 13568
rect 11789 13560 15578 13562
rect 11789 13504 11794 13560
rect 11850 13504 15578 13560
rect 11789 13502 15578 13504
rect 22829 13562 22895 13565
rect 23289 13562 23355 13565
rect 22829 13560 23355 13562
rect 22829 13504 22834 13560
rect 22890 13504 23294 13560
rect 23350 13504 23355 13560
rect 22829 13502 23355 13504
rect 11789 13499 11855 13502
rect 22829 13499 22895 13502
rect 23289 13499 23355 13502
rect 4061 13426 4127 13429
rect 16757 13426 16823 13429
rect 4061 13424 16823 13426
rect 4061 13368 4066 13424
rect 4122 13368 16762 13424
rect 16818 13368 16823 13424
rect 4061 13366 16823 13368
rect 4061 13363 4127 13366
rect 16757 13363 16823 13366
rect 20345 13426 20411 13429
rect 30741 13426 30807 13429
rect 20345 13424 30807 13426
rect 20345 13368 20350 13424
rect 20406 13368 30746 13424
rect 30802 13368 30807 13424
rect 20345 13366 30807 13368
rect 20345 13363 20411 13366
rect 30741 13363 30807 13366
rect 3049 13290 3115 13293
rect 15561 13290 15627 13293
rect 3049 13288 15627 13290
rect 3049 13232 3054 13288
rect 3110 13232 15566 13288
rect 15622 13232 15627 13288
rect 3049 13230 15627 13232
rect 3049 13227 3115 13230
rect 15561 13227 15627 13230
rect 19333 13290 19399 13293
rect 21357 13290 21423 13293
rect 19333 13288 21423 13290
rect 19333 13232 19338 13288
rect 19394 13232 21362 13288
rect 21418 13232 21423 13288
rect 19333 13230 21423 13232
rect 19333 13227 19399 13230
rect 21357 13227 21423 13230
rect 22185 13290 22251 13293
rect 23473 13290 23539 13293
rect 22185 13288 23539 13290
rect 22185 13232 22190 13288
rect 22246 13232 23478 13288
rect 23534 13232 23539 13288
rect 22185 13230 23539 13232
rect 22185 13227 22251 13230
rect 23473 13227 23539 13230
rect 13629 13154 13695 13157
rect 15653 13154 15719 13157
rect 13629 13152 15719 13154
rect 13629 13096 13634 13152
rect 13690 13096 15658 13152
rect 15714 13096 15719 13152
rect 13629 13094 15719 13096
rect 13629 13091 13695 13094
rect 15653 13091 15719 13094
rect 16481 13154 16547 13157
rect 17769 13154 17835 13157
rect 16481 13152 17835 13154
rect 16481 13096 16486 13152
rect 16542 13096 17774 13152
rect 17830 13096 17835 13152
rect 16481 13094 17835 13096
rect 16481 13091 16547 13094
rect 17769 13091 17835 13094
rect 4246 13088 4562 13089
rect 4246 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4562 13088
rect 4246 13023 4562 13024
rect 11951 13088 12267 13089
rect 11951 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12267 13088
rect 11951 13023 12267 13024
rect 19656 13088 19972 13089
rect 19656 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19972 13088
rect 19656 13023 19972 13024
rect 27361 13088 27677 13089
rect 27361 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27677 13088
rect 27361 13023 27677 13024
rect 16849 13018 16915 13021
rect 19190 13018 19196 13020
rect 12390 12958 14658 13018
rect 6821 12882 6887 12885
rect 12390 12882 12450 12958
rect 6821 12880 12450 12882
rect 6821 12824 6826 12880
rect 6882 12824 12450 12880
rect 6821 12822 12450 12824
rect 14273 12882 14339 12885
rect 14406 12882 14412 12884
rect 14273 12880 14412 12882
rect 14273 12824 14278 12880
rect 14334 12824 14412 12880
rect 14273 12822 14412 12824
rect 6821 12819 6887 12822
rect 14273 12819 14339 12822
rect 14406 12820 14412 12822
rect 14476 12820 14482 12884
rect 14598 12882 14658 12958
rect 16849 13016 19196 13018
rect 16849 12960 16854 13016
rect 16910 12960 19196 13016
rect 16849 12958 19196 12960
rect 16849 12955 16915 12958
rect 19190 12956 19196 12958
rect 19260 12956 19266 13020
rect 20161 12882 20227 12885
rect 14598 12880 20227 12882
rect 14598 12824 20166 12880
rect 20222 12824 20227 12880
rect 14598 12822 20227 12824
rect 20161 12819 20227 12822
rect 10869 12746 10935 12749
rect 17769 12746 17835 12749
rect 10869 12744 17835 12746
rect 10869 12688 10874 12744
rect 10930 12688 17774 12744
rect 17830 12688 17835 12744
rect 10869 12686 17835 12688
rect 10869 12683 10935 12686
rect 17769 12683 17835 12686
rect 13905 12610 13971 12613
rect 14038 12610 14044 12612
rect 13905 12608 14044 12610
rect 13905 12552 13910 12608
rect 13966 12552 14044 12608
rect 13905 12550 14044 12552
rect 13905 12547 13971 12550
rect 14038 12548 14044 12550
rect 14108 12548 14114 12612
rect 8098 12544 8414 12545
rect 8098 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8414 12544
rect 8098 12479 8414 12480
rect 15803 12544 16119 12545
rect 15803 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16119 12544
rect 15803 12479 16119 12480
rect 23508 12544 23824 12545
rect 23508 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23824 12544
rect 23508 12479 23824 12480
rect 31213 12544 31529 12545
rect 31213 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31529 12544
rect 31213 12479 31529 12480
rect 10041 12474 10107 12477
rect 13905 12474 13971 12477
rect 15469 12474 15535 12477
rect 10041 12472 15535 12474
rect 10041 12416 10046 12472
rect 10102 12416 13910 12472
rect 13966 12416 15474 12472
rect 15530 12416 15535 12472
rect 10041 12414 15535 12416
rect 10041 12411 10107 12414
rect 13905 12411 13971 12414
rect 15469 12411 15535 12414
rect 16481 12474 16547 12477
rect 18597 12474 18663 12477
rect 16481 12472 18663 12474
rect 16481 12416 16486 12472
rect 16542 12416 18602 12472
rect 18658 12416 18663 12472
rect 16481 12414 18663 12416
rect 16481 12411 16547 12414
rect 18597 12411 18663 12414
rect 3049 12338 3115 12341
rect 16021 12338 16087 12341
rect 18137 12338 18203 12341
rect 3049 12336 16087 12338
rect 3049 12280 3054 12336
rect 3110 12280 16026 12336
rect 16082 12280 16087 12336
rect 3049 12278 16087 12280
rect 3049 12275 3115 12278
rect 16021 12275 16087 12278
rect 17542 12336 18203 12338
rect 17542 12280 18142 12336
rect 18198 12280 18203 12336
rect 17542 12278 18203 12280
rect 3969 12202 4035 12205
rect 6453 12202 6519 12205
rect 15929 12202 15995 12205
rect 17542 12202 17602 12278
rect 18137 12275 18203 12278
rect 19885 12338 19951 12341
rect 25313 12338 25379 12341
rect 19885 12336 25379 12338
rect 19885 12280 19890 12336
rect 19946 12280 25318 12336
rect 25374 12280 25379 12336
rect 19885 12278 25379 12280
rect 19885 12275 19951 12278
rect 25313 12275 25379 12278
rect 28625 12338 28691 12341
rect 31600 12338 32000 12368
rect 28625 12336 32000 12338
rect 28625 12280 28630 12336
rect 28686 12280 32000 12336
rect 28625 12278 32000 12280
rect 28625 12275 28691 12278
rect 31600 12248 32000 12278
rect 3969 12200 4722 12202
rect 3969 12144 3974 12200
rect 4030 12144 4722 12200
rect 3969 12142 4722 12144
rect 3969 12139 4035 12142
rect 4662 12066 4722 12142
rect 6453 12200 12450 12202
rect 6453 12144 6458 12200
rect 6514 12144 12450 12200
rect 6453 12142 12450 12144
rect 6453 12139 6519 12142
rect 4662 12006 10610 12066
rect 4246 12000 4562 12001
rect 4246 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4562 12000
rect 4246 11935 4562 11936
rect 10550 11794 10610 12006
rect 11951 12000 12267 12001
rect 11951 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12267 12000
rect 11951 11935 12267 11936
rect 12390 11930 12450 12142
rect 15929 12200 17602 12202
rect 15929 12144 15934 12200
rect 15990 12144 17602 12200
rect 15929 12142 17602 12144
rect 24393 12202 24459 12205
rect 24393 12200 24594 12202
rect 24393 12144 24398 12200
rect 24454 12144 24594 12200
rect 24393 12142 24594 12144
rect 15929 12139 15995 12142
rect 24393 12139 24459 12142
rect 15193 12066 15259 12069
rect 18781 12066 18847 12069
rect 15193 12064 18847 12066
rect 15193 12008 15198 12064
rect 15254 12008 18786 12064
rect 18842 12008 18847 12064
rect 15193 12006 18847 12008
rect 15193 12003 15259 12006
rect 18781 12003 18847 12006
rect 20345 12066 20411 12069
rect 21633 12066 21699 12069
rect 20345 12064 21699 12066
rect 20345 12008 20350 12064
rect 20406 12008 21638 12064
rect 21694 12008 21699 12064
rect 20345 12006 21699 12008
rect 20345 12003 20411 12006
rect 21633 12003 21699 12006
rect 19656 12000 19972 12001
rect 19656 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19972 12000
rect 19656 11935 19972 11936
rect 18413 11930 18479 11933
rect 12390 11928 18479 11930
rect 12390 11872 18418 11928
rect 18474 11872 18479 11928
rect 12390 11870 18479 11872
rect 18413 11867 18479 11870
rect 24534 11797 24594 12142
rect 27361 12000 27677 12001
rect 27361 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27677 12000
rect 27361 11935 27677 11936
rect 13813 11794 13879 11797
rect 7974 11734 10426 11794
rect 10550 11792 13879 11794
rect 10550 11736 13818 11792
rect 13874 11736 13879 11792
rect 10550 11734 13879 11736
rect 6269 11658 6335 11661
rect 7974 11658 8034 11734
rect 6269 11656 8034 11658
rect 6269 11600 6274 11656
rect 6330 11600 8034 11656
rect 6269 11598 8034 11600
rect 8109 11658 8175 11661
rect 10366 11658 10426 11734
rect 13813 11731 13879 11734
rect 15009 11794 15075 11797
rect 16021 11794 16087 11797
rect 15009 11792 16087 11794
rect 15009 11736 15014 11792
rect 15070 11736 16026 11792
rect 16082 11736 16087 11792
rect 15009 11734 16087 11736
rect 15009 11731 15075 11734
rect 16021 11731 16087 11734
rect 16849 11794 16915 11797
rect 17902 11794 17908 11796
rect 16849 11792 17908 11794
rect 16849 11736 16854 11792
rect 16910 11736 17908 11792
rect 16849 11734 17908 11736
rect 16849 11731 16915 11734
rect 17902 11732 17908 11734
rect 17972 11732 17978 11796
rect 18873 11794 18939 11797
rect 19057 11794 19123 11797
rect 18873 11792 19123 11794
rect 18873 11736 18878 11792
rect 18934 11736 19062 11792
rect 19118 11736 19123 11792
rect 18873 11734 19123 11736
rect 18873 11731 18939 11734
rect 19057 11731 19123 11734
rect 19793 11794 19859 11797
rect 20069 11794 20135 11797
rect 19793 11792 20135 11794
rect 19793 11736 19798 11792
rect 19854 11736 20074 11792
rect 20130 11736 20135 11792
rect 19793 11734 20135 11736
rect 19793 11731 19859 11734
rect 20069 11731 20135 11734
rect 22001 11794 22067 11797
rect 24025 11794 24091 11797
rect 22001 11792 24091 11794
rect 22001 11736 22006 11792
rect 22062 11736 24030 11792
rect 24086 11736 24091 11792
rect 22001 11734 24091 11736
rect 24534 11792 24643 11797
rect 24534 11736 24582 11792
rect 24638 11736 24643 11792
rect 24534 11734 24643 11736
rect 22001 11731 22067 11734
rect 24025 11731 24091 11734
rect 24577 11731 24643 11734
rect 19333 11658 19399 11661
rect 8109 11656 10242 11658
rect 8109 11600 8114 11656
rect 8170 11600 10242 11656
rect 8109 11598 10242 11600
rect 10366 11656 19399 11658
rect 10366 11600 19338 11656
rect 19394 11600 19399 11656
rect 10366 11598 19399 11600
rect 6269 11595 6335 11598
rect 8109 11595 8175 11598
rect 8098 11456 8414 11457
rect 8098 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8414 11456
rect 8098 11391 8414 11392
rect 10182 11250 10242 11598
rect 19333 11595 19399 11598
rect 19701 11658 19767 11661
rect 20805 11658 20871 11661
rect 19701 11656 20871 11658
rect 19701 11600 19706 11656
rect 19762 11600 20810 11656
rect 20866 11600 20871 11656
rect 19701 11598 20871 11600
rect 19701 11595 19767 11598
rect 20805 11595 20871 11598
rect 11973 11522 12039 11525
rect 14181 11522 14247 11525
rect 11973 11520 14247 11522
rect 11973 11464 11978 11520
rect 12034 11464 14186 11520
rect 14242 11464 14247 11520
rect 11973 11462 14247 11464
rect 11973 11459 12039 11462
rect 14181 11459 14247 11462
rect 16205 11522 16271 11525
rect 16573 11522 16639 11525
rect 16205 11520 16639 11522
rect 16205 11464 16210 11520
rect 16266 11464 16578 11520
rect 16634 11464 16639 11520
rect 16205 11462 16639 11464
rect 16205 11459 16271 11462
rect 16573 11459 16639 11462
rect 16757 11524 16823 11525
rect 16757 11520 16804 11524
rect 16868 11522 16874 11524
rect 17677 11522 17743 11525
rect 23197 11522 23263 11525
rect 16757 11464 16762 11520
rect 16757 11460 16804 11464
rect 16868 11462 16914 11522
rect 17677 11520 23263 11522
rect 17677 11464 17682 11520
rect 17738 11464 23202 11520
rect 23258 11464 23263 11520
rect 17677 11462 23263 11464
rect 16868 11460 16874 11462
rect 16757 11459 16823 11460
rect 17677 11459 17743 11462
rect 23197 11459 23263 11462
rect 15803 11456 16119 11457
rect 15803 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16119 11456
rect 15803 11391 16119 11392
rect 23508 11456 23824 11457
rect 23508 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23824 11456
rect 23508 11391 23824 11392
rect 31213 11456 31529 11457
rect 31213 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31529 11456
rect 31213 11391 31529 11392
rect 15142 11324 15148 11388
rect 15212 11386 15218 11388
rect 15653 11386 15719 11389
rect 17401 11386 17467 11389
rect 15212 11384 15719 11386
rect 15212 11328 15658 11384
rect 15714 11328 15719 11384
rect 15212 11326 15719 11328
rect 15212 11324 15218 11326
rect 15653 11323 15719 11326
rect 16254 11384 17467 11386
rect 16254 11328 17406 11384
rect 17462 11328 17467 11384
rect 16254 11326 17467 11328
rect 16254 11250 16314 11326
rect 17401 11323 17467 11326
rect 20069 11386 20135 11389
rect 20805 11386 20871 11389
rect 20069 11384 20871 11386
rect 20069 11328 20074 11384
rect 20130 11328 20810 11384
rect 20866 11328 20871 11384
rect 20069 11326 20871 11328
rect 20069 11323 20135 11326
rect 20805 11323 20871 11326
rect 22737 11386 22803 11389
rect 23013 11386 23079 11389
rect 22737 11384 23079 11386
rect 22737 11328 22742 11384
rect 22798 11328 23018 11384
rect 23074 11328 23079 11384
rect 22737 11326 23079 11328
rect 22737 11323 22803 11326
rect 23013 11323 23079 11326
rect 10182 11190 16314 11250
rect 17033 11250 17099 11253
rect 27705 11250 27771 11253
rect 17033 11248 27771 11250
rect 17033 11192 17038 11248
rect 17094 11192 27710 11248
rect 27766 11192 27771 11248
rect 17033 11190 27771 11192
rect 17033 11187 17099 11190
rect 27705 11187 27771 11190
rect 9673 11114 9739 11117
rect 16849 11114 16915 11117
rect 9673 11112 16915 11114
rect 9673 11056 9678 11112
rect 9734 11056 16854 11112
rect 16910 11056 16915 11112
rect 9673 11054 16915 11056
rect 9673 11051 9739 11054
rect 16849 11051 16915 11054
rect 16246 10978 16252 10980
rect 14598 10918 16252 10978
rect 4246 10912 4562 10913
rect 4246 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4562 10912
rect 4246 10847 4562 10848
rect 11951 10912 12267 10913
rect 11951 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12267 10912
rect 11951 10847 12267 10848
rect 7925 10706 7991 10709
rect 14598 10706 14658 10918
rect 16246 10916 16252 10918
rect 16316 10978 16322 10980
rect 17217 10978 17283 10981
rect 17401 10978 17467 10981
rect 16316 10976 17467 10978
rect 16316 10920 17222 10976
rect 17278 10920 17406 10976
rect 17462 10920 17467 10976
rect 16316 10918 17467 10920
rect 16316 10916 16322 10918
rect 17217 10915 17283 10918
rect 17401 10915 17467 10918
rect 19656 10912 19972 10913
rect 19656 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19972 10912
rect 19656 10847 19972 10848
rect 27361 10912 27677 10913
rect 27361 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27677 10912
rect 27361 10847 27677 10848
rect 15745 10842 15811 10845
rect 16573 10842 16639 10845
rect 15745 10840 16639 10842
rect 15745 10784 15750 10840
rect 15806 10784 16578 10840
rect 16634 10784 16639 10840
rect 15745 10782 16639 10784
rect 15745 10779 15811 10782
rect 16573 10779 16639 10782
rect 16757 10842 16823 10845
rect 18873 10842 18939 10845
rect 16757 10840 18939 10842
rect 16757 10784 16762 10840
rect 16818 10784 18878 10840
rect 18934 10784 18939 10840
rect 16757 10782 18939 10784
rect 16757 10779 16823 10782
rect 18873 10779 18939 10782
rect 7925 10704 14658 10706
rect 7925 10648 7930 10704
rect 7986 10648 14658 10704
rect 7925 10646 14658 10648
rect 14733 10706 14799 10709
rect 18321 10706 18387 10709
rect 19885 10706 19951 10709
rect 14733 10704 18387 10706
rect 14733 10648 14738 10704
rect 14794 10648 18326 10704
rect 18382 10648 18387 10704
rect 14733 10646 18387 10648
rect 7925 10643 7991 10646
rect 14733 10643 14799 10646
rect 18321 10643 18387 10646
rect 18462 10704 19951 10706
rect 18462 10648 19890 10704
rect 19946 10648 19951 10704
rect 18462 10646 19951 10648
rect 11237 10570 11303 10573
rect 15745 10570 15811 10573
rect 11237 10568 15811 10570
rect 11237 10512 11242 10568
rect 11298 10512 15750 10568
rect 15806 10512 15811 10568
rect 11237 10510 15811 10512
rect 11237 10507 11303 10510
rect 15745 10507 15811 10510
rect 15929 10570 15995 10573
rect 16430 10570 16436 10572
rect 15929 10568 16436 10570
rect 15929 10512 15934 10568
rect 15990 10512 16436 10568
rect 15929 10510 16436 10512
rect 15929 10507 15995 10510
rect 16430 10508 16436 10510
rect 16500 10508 16506 10572
rect 10041 10434 10107 10437
rect 14181 10434 14247 10437
rect 10041 10432 14247 10434
rect 10041 10376 10046 10432
rect 10102 10376 14186 10432
rect 14242 10376 14247 10432
rect 10041 10374 14247 10376
rect 10041 10371 10107 10374
rect 14181 10371 14247 10374
rect 16205 10434 16271 10437
rect 18462 10434 18522 10646
rect 19885 10643 19951 10646
rect 19190 10508 19196 10572
rect 19260 10570 19266 10572
rect 23013 10570 23079 10573
rect 19260 10568 23079 10570
rect 19260 10512 23018 10568
rect 23074 10512 23079 10568
rect 19260 10510 23079 10512
rect 19260 10508 19266 10510
rect 23013 10507 23079 10510
rect 16205 10432 18522 10434
rect 16205 10376 16210 10432
rect 16266 10376 18522 10432
rect 16205 10374 18522 10376
rect 19701 10434 19767 10437
rect 23289 10434 23355 10437
rect 19701 10432 23355 10434
rect 19701 10376 19706 10432
rect 19762 10376 23294 10432
rect 23350 10376 23355 10432
rect 19701 10374 23355 10376
rect 16205 10371 16271 10374
rect 19701 10371 19767 10374
rect 23289 10371 23355 10374
rect 8098 10368 8414 10369
rect 8098 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8414 10368
rect 8098 10303 8414 10304
rect 15803 10368 16119 10369
rect 15803 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16119 10368
rect 15803 10303 16119 10304
rect 23508 10368 23824 10369
rect 23508 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23824 10368
rect 23508 10303 23824 10304
rect 31213 10368 31529 10369
rect 31213 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31529 10368
rect 31213 10303 31529 10304
rect 13997 10298 14063 10301
rect 16297 10298 16363 10301
rect 18137 10298 18203 10301
rect 13997 10296 15716 10298
rect 13997 10240 14002 10296
rect 14058 10240 15716 10296
rect 13997 10238 15716 10240
rect 13997 10235 14063 10238
rect 14273 10162 14339 10165
rect 14774 10162 14780 10164
rect 14273 10160 14780 10162
rect 14273 10104 14278 10160
rect 14334 10104 14780 10160
rect 14273 10102 14780 10104
rect 14273 10099 14339 10102
rect 14774 10100 14780 10102
rect 14844 10100 14850 10164
rect 15656 10162 15716 10238
rect 16297 10296 18203 10298
rect 16297 10240 16302 10296
rect 16358 10240 18142 10296
rect 18198 10240 18203 10296
rect 16297 10238 18203 10240
rect 16297 10235 16363 10238
rect 18137 10235 18203 10238
rect 31600 10296 32000 10328
rect 31600 10240 31666 10296
rect 31722 10240 32000 10296
rect 31600 10208 32000 10240
rect 17217 10162 17283 10165
rect 17769 10164 17835 10165
rect 15656 10160 17283 10162
rect 15656 10104 17222 10160
rect 17278 10104 17283 10160
rect 15656 10102 17283 10104
rect 17217 10099 17283 10102
rect 17718 10100 17724 10164
rect 17788 10162 17835 10164
rect 17788 10160 17880 10162
rect 17830 10104 17880 10160
rect 17788 10102 17880 10104
rect 17788 10100 17835 10102
rect 19374 10100 19380 10164
rect 19444 10162 19450 10164
rect 19793 10162 19859 10165
rect 19444 10160 19859 10162
rect 19444 10104 19798 10160
rect 19854 10104 19859 10160
rect 19444 10102 19859 10104
rect 19444 10100 19450 10102
rect 17769 10099 17835 10100
rect 19793 10099 19859 10102
rect 21541 10162 21607 10165
rect 26877 10162 26943 10165
rect 21541 10160 26943 10162
rect 21541 10104 21546 10160
rect 21602 10104 26882 10160
rect 26938 10104 26943 10160
rect 21541 10102 26943 10104
rect 21541 10099 21607 10102
rect 26877 10099 26943 10102
rect 14273 10026 14339 10029
rect 23197 10026 23263 10029
rect 14273 10024 23263 10026
rect 14273 9968 14278 10024
rect 14334 9968 23202 10024
rect 23258 9968 23263 10024
rect 14273 9966 23263 9968
rect 14273 9963 14339 9966
rect 23197 9963 23263 9966
rect 12433 9890 12499 9893
rect 14641 9890 14707 9893
rect 12433 9888 14707 9890
rect 12433 9832 12438 9888
rect 12494 9832 14646 9888
rect 14702 9832 14707 9888
rect 12433 9830 14707 9832
rect 12433 9827 12499 9830
rect 14641 9827 14707 9830
rect 15745 9890 15811 9893
rect 19241 9890 19307 9893
rect 15745 9888 19307 9890
rect 15745 9832 15750 9888
rect 15806 9832 19246 9888
rect 19302 9832 19307 9888
rect 15745 9830 19307 9832
rect 15745 9827 15811 9830
rect 19241 9827 19307 9830
rect 4246 9824 4562 9825
rect 4246 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4562 9824
rect 4246 9759 4562 9760
rect 11951 9824 12267 9825
rect 11951 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12267 9824
rect 11951 9759 12267 9760
rect 19656 9824 19972 9825
rect 19656 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19972 9824
rect 19656 9759 19972 9760
rect 27361 9824 27677 9825
rect 27361 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27677 9824
rect 27361 9759 27677 9760
rect 13261 9754 13327 9757
rect 14917 9754 14983 9757
rect 13261 9752 14983 9754
rect 13261 9696 13266 9752
rect 13322 9696 14922 9752
rect 14978 9696 14983 9752
rect 13261 9694 14983 9696
rect 13261 9691 13327 9694
rect 14917 9691 14983 9694
rect 15285 9754 15351 9757
rect 21357 9754 21423 9757
rect 15285 9752 19442 9754
rect 15285 9696 15290 9752
rect 15346 9696 19442 9752
rect 15285 9694 19442 9696
rect 15285 9691 15351 9694
rect 14917 9620 14983 9621
rect 14917 9618 14964 9620
rect 14872 9616 14964 9618
rect 14872 9560 14922 9616
rect 14872 9558 14964 9560
rect 14917 9556 14964 9558
rect 15028 9556 15034 9620
rect 15510 9556 15516 9620
rect 15580 9618 15586 9620
rect 16113 9618 16179 9621
rect 16665 9620 16731 9621
rect 17585 9620 17651 9621
rect 15580 9616 16179 9618
rect 15580 9560 16118 9616
rect 16174 9560 16179 9616
rect 15580 9558 16179 9560
rect 15580 9556 15586 9558
rect 14917 9555 14983 9556
rect 16113 9555 16179 9558
rect 16614 9556 16620 9620
rect 16684 9618 16731 9620
rect 16684 9616 16776 9618
rect 16726 9560 16776 9616
rect 16684 9558 16776 9560
rect 16684 9556 16731 9558
rect 17534 9556 17540 9620
rect 17604 9618 17651 9620
rect 18689 9618 18755 9621
rect 18822 9618 18828 9620
rect 17604 9616 17696 9618
rect 17646 9560 17696 9616
rect 17604 9558 17696 9560
rect 18689 9616 18828 9618
rect 18689 9560 18694 9616
rect 18750 9560 18828 9616
rect 18689 9558 18828 9560
rect 17604 9556 17651 9558
rect 16665 9555 16731 9556
rect 17585 9555 17651 9556
rect 18689 9555 18755 9558
rect 18822 9556 18828 9558
rect 18892 9556 18898 9620
rect 19382 9618 19442 9694
rect 20118 9752 21423 9754
rect 20118 9696 21362 9752
rect 21418 9696 21423 9752
rect 20118 9694 21423 9696
rect 20118 9618 20178 9694
rect 21357 9691 21423 9694
rect 19382 9558 20178 9618
rect 20529 9618 20595 9621
rect 22369 9618 22435 9621
rect 20529 9616 22435 9618
rect 20529 9560 20534 9616
rect 20590 9560 22374 9616
rect 22430 9560 22435 9616
rect 20529 9558 22435 9560
rect 20529 9555 20595 9558
rect 22369 9555 22435 9558
rect 25681 9618 25747 9621
rect 31600 9618 32000 9648
rect 25681 9616 32000 9618
rect 25681 9560 25686 9616
rect 25742 9560 32000 9616
rect 25681 9558 32000 9560
rect 25681 9555 25747 9558
rect 31600 9528 32000 9558
rect 14273 9482 14339 9485
rect 15193 9482 15259 9485
rect 14273 9480 15259 9482
rect 14273 9424 14278 9480
rect 14334 9424 15198 9480
rect 15254 9424 15259 9480
rect 14273 9422 15259 9424
rect 14273 9419 14339 9422
rect 15193 9419 15259 9422
rect 15745 9482 15811 9485
rect 16982 9482 16988 9484
rect 15745 9480 16988 9482
rect 15745 9424 15750 9480
rect 15806 9424 16988 9480
rect 15745 9422 16988 9424
rect 15745 9419 15811 9422
rect 16982 9420 16988 9422
rect 17052 9420 17058 9484
rect 17166 9420 17172 9484
rect 17236 9482 17242 9484
rect 26325 9482 26391 9485
rect 17236 9480 26391 9482
rect 17236 9424 26330 9480
rect 26386 9424 26391 9480
rect 17236 9422 26391 9424
rect 17236 9420 17242 9422
rect 26325 9419 26391 9422
rect 18045 9346 18111 9349
rect 16254 9344 18111 9346
rect 16254 9288 18050 9344
rect 18106 9288 18111 9344
rect 16254 9286 18111 9288
rect 8098 9280 8414 9281
rect 8098 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8414 9280
rect 8098 9215 8414 9216
rect 15803 9280 16119 9281
rect 15803 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16119 9280
rect 15803 9215 16119 9216
rect 7741 9074 7807 9077
rect 16254 9074 16314 9286
rect 18045 9283 18111 9286
rect 23508 9280 23824 9281
rect 23508 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23824 9280
rect 23508 9215 23824 9216
rect 31213 9280 31529 9281
rect 31213 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31529 9280
rect 31213 9215 31529 9216
rect 16389 9210 16455 9213
rect 20437 9210 20503 9213
rect 16389 9208 20503 9210
rect 16389 9152 16394 9208
rect 16450 9152 20442 9208
rect 20498 9152 20503 9208
rect 16389 9150 20503 9152
rect 16389 9147 16455 9150
rect 20437 9147 20503 9150
rect 24117 9210 24183 9213
rect 30925 9210 30991 9213
rect 24117 9208 30991 9210
rect 24117 9152 24122 9208
rect 24178 9152 30930 9208
rect 30986 9152 30991 9208
rect 24117 9150 30991 9152
rect 24117 9147 24183 9150
rect 30925 9147 30991 9150
rect 17033 9076 17099 9077
rect 7741 9072 16314 9074
rect 7741 9016 7746 9072
rect 7802 9016 16314 9072
rect 7741 9014 16314 9016
rect 7741 9011 7807 9014
rect 16982 9012 16988 9076
rect 17052 9074 17099 9076
rect 17585 9074 17651 9077
rect 18505 9076 18571 9077
rect 18454 9074 18460 9076
rect 17052 9072 17144 9074
rect 17094 9016 17144 9072
rect 17052 9014 17144 9016
rect 17585 9072 18460 9074
rect 18524 9074 18571 9076
rect 19885 9074 19951 9077
rect 24485 9074 24551 9077
rect 18524 9072 18616 9074
rect 17585 9016 17590 9072
rect 17646 9016 18460 9072
rect 18566 9016 18616 9072
rect 17585 9014 18460 9016
rect 17052 9012 17099 9014
rect 17033 9011 17099 9012
rect 17585 9011 17651 9014
rect 18454 9012 18460 9014
rect 18524 9014 18616 9016
rect 19885 9072 24551 9074
rect 19885 9016 19890 9072
rect 19946 9016 24490 9072
rect 24546 9016 24551 9072
rect 19885 9014 24551 9016
rect 18524 9012 18571 9014
rect 18505 9011 18571 9012
rect 19885 9011 19951 9014
rect 24485 9011 24551 9014
rect 13445 8938 13511 8941
rect 24761 8938 24827 8941
rect 13445 8936 24827 8938
rect 13445 8880 13450 8936
rect 13506 8880 24766 8936
rect 24822 8880 24827 8936
rect 13445 8878 24827 8880
rect 13445 8875 13511 8878
rect 24761 8875 24827 8878
rect 16665 8802 16731 8805
rect 17677 8804 17743 8805
rect 17534 8802 17540 8804
rect 16665 8800 17540 8802
rect 16665 8744 16670 8800
rect 16726 8744 17540 8800
rect 16665 8742 17540 8744
rect 16665 8739 16731 8742
rect 17534 8740 17540 8742
rect 17604 8740 17610 8804
rect 17677 8800 17724 8804
rect 17788 8802 17794 8804
rect 20437 8802 20503 8805
rect 24853 8802 24919 8805
rect 17677 8744 17682 8800
rect 17677 8740 17724 8744
rect 17788 8742 17834 8802
rect 20437 8800 24919 8802
rect 20437 8744 20442 8800
rect 20498 8744 24858 8800
rect 24914 8744 24919 8800
rect 20437 8742 24919 8744
rect 17788 8740 17794 8742
rect 17677 8739 17743 8740
rect 20437 8739 20503 8742
rect 24853 8739 24919 8742
rect 4246 8736 4562 8737
rect 4246 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4562 8736
rect 4246 8671 4562 8672
rect 11951 8736 12267 8737
rect 11951 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12267 8736
rect 11951 8671 12267 8672
rect 19656 8736 19972 8737
rect 19656 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19972 8736
rect 19656 8671 19972 8672
rect 27361 8736 27677 8737
rect 27361 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27677 8736
rect 27361 8671 27677 8672
rect 12709 8666 12775 8669
rect 14549 8666 14615 8669
rect 12709 8664 14615 8666
rect 12709 8608 12714 8664
rect 12770 8608 14554 8664
rect 14610 8608 14615 8664
rect 12709 8606 14615 8608
rect 12709 8603 12775 8606
rect 14549 8603 14615 8606
rect 14958 8604 14964 8668
rect 15028 8666 15034 8668
rect 16573 8666 16639 8669
rect 15028 8664 16639 8666
rect 15028 8608 16578 8664
rect 16634 8608 16639 8664
rect 15028 8606 16639 8608
rect 15028 8604 15034 8606
rect 16573 8603 16639 8606
rect 7373 8530 7439 8533
rect 19149 8530 19215 8533
rect 7373 8528 19215 8530
rect 7373 8472 7378 8528
rect 7434 8472 19154 8528
rect 19210 8472 19215 8528
rect 7373 8470 19215 8472
rect 7373 8467 7439 8470
rect 19149 8467 19215 8470
rect 12709 8394 12775 8397
rect 13670 8394 13676 8396
rect 12709 8392 13676 8394
rect 12709 8336 12714 8392
rect 12770 8336 13676 8392
rect 12709 8334 13676 8336
rect 12709 8331 12775 8334
rect 13670 8332 13676 8334
rect 13740 8332 13746 8396
rect 15469 8394 15535 8397
rect 17166 8394 17172 8396
rect 15469 8392 17172 8394
rect 15469 8336 15474 8392
rect 15530 8336 17172 8392
rect 15469 8334 17172 8336
rect 15469 8331 15535 8334
rect 17166 8332 17172 8334
rect 17236 8332 17242 8396
rect 17309 8394 17375 8397
rect 18505 8394 18571 8397
rect 17309 8392 18571 8394
rect 17309 8336 17314 8392
rect 17370 8336 18510 8392
rect 18566 8336 18571 8392
rect 17309 8334 18571 8336
rect 17309 8331 17375 8334
rect 18505 8331 18571 8334
rect 16430 8196 16436 8260
rect 16500 8258 16506 8260
rect 20437 8258 20503 8261
rect 16500 8256 20503 8258
rect 16500 8200 20442 8256
rect 20498 8200 20503 8256
rect 16500 8198 20503 8200
rect 16500 8196 16506 8198
rect 20437 8195 20503 8198
rect 20621 8258 20687 8261
rect 23105 8258 23171 8261
rect 20621 8256 23171 8258
rect 20621 8200 20626 8256
rect 20682 8200 23110 8256
rect 23166 8200 23171 8256
rect 20621 8198 23171 8200
rect 20621 8195 20687 8198
rect 23105 8195 23171 8198
rect 8098 8192 8414 8193
rect 8098 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8414 8192
rect 8098 8127 8414 8128
rect 15803 8192 16119 8193
rect 15803 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16119 8192
rect 15803 8127 16119 8128
rect 23508 8192 23824 8193
rect 23508 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23824 8192
rect 23508 8127 23824 8128
rect 31213 8192 31529 8193
rect 31213 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31529 8192
rect 31213 8127 31529 8128
rect 13445 8122 13511 8125
rect 14549 8122 14615 8125
rect 13445 8120 14615 8122
rect 13445 8064 13450 8120
rect 13506 8064 14554 8120
rect 14610 8064 14615 8120
rect 13445 8062 14615 8064
rect 13445 8059 13511 8062
rect 14549 8059 14615 8062
rect 16941 8122 17007 8125
rect 19374 8122 19380 8124
rect 16941 8120 19380 8122
rect 16941 8064 16946 8120
rect 17002 8064 19380 8120
rect 16941 8062 19380 8064
rect 16941 8059 17007 8062
rect 19374 8060 19380 8062
rect 19444 8060 19450 8124
rect 14273 7986 14339 7989
rect 18229 7986 18295 7989
rect 14273 7984 18295 7986
rect 14273 7928 14278 7984
rect 14334 7928 18234 7984
rect 18290 7928 18295 7984
rect 14273 7926 18295 7928
rect 14273 7923 14339 7926
rect 18229 7923 18295 7926
rect 19701 7986 19767 7989
rect 30925 7986 30991 7989
rect 19701 7984 30991 7986
rect 19701 7928 19706 7984
rect 19762 7928 30930 7984
rect 30986 7928 30991 7984
rect 19701 7926 30991 7928
rect 19701 7923 19767 7926
rect 30925 7923 30991 7926
rect 14917 7850 14983 7853
rect 16573 7850 16639 7853
rect 14917 7848 16639 7850
rect 14917 7792 14922 7848
rect 14978 7792 16578 7848
rect 16634 7792 16639 7848
rect 14917 7790 16639 7792
rect 14917 7787 14983 7790
rect 16573 7787 16639 7790
rect 18965 7850 19031 7853
rect 26693 7850 26759 7853
rect 18965 7848 26759 7850
rect 18965 7792 18970 7848
rect 19026 7792 26698 7848
rect 26754 7792 26759 7848
rect 18965 7790 26759 7792
rect 18965 7787 19031 7790
rect 26693 7787 26759 7790
rect 4246 7648 4562 7649
rect 4246 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4562 7648
rect 4246 7583 4562 7584
rect 11951 7648 12267 7649
rect 11951 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12267 7648
rect 11951 7583 12267 7584
rect 19656 7648 19972 7649
rect 19656 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19972 7648
rect 19656 7583 19972 7584
rect 27361 7648 27677 7649
rect 27361 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27677 7648
rect 27361 7583 27677 7584
rect 8098 7104 8414 7105
rect 8098 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8414 7104
rect 8098 7039 8414 7040
rect 15803 7104 16119 7105
rect 15803 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16119 7104
rect 15803 7039 16119 7040
rect 23508 7104 23824 7105
rect 23508 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23824 7104
rect 23508 7039 23824 7040
rect 31213 7104 31529 7105
rect 31213 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31529 7104
rect 31213 7039 31529 7040
rect 12801 7034 12867 7037
rect 15101 7034 15167 7037
rect 12801 7032 15167 7034
rect 12801 6976 12806 7032
rect 12862 6976 15106 7032
rect 15162 6976 15167 7032
rect 12801 6974 15167 6976
rect 12801 6971 12867 6974
rect 15101 6971 15167 6974
rect 13721 6898 13787 6901
rect 14038 6898 14044 6900
rect 13721 6896 14044 6898
rect 13721 6840 13726 6896
rect 13782 6840 14044 6896
rect 13721 6838 14044 6840
rect 13721 6835 13787 6838
rect 14038 6836 14044 6838
rect 14108 6836 14114 6900
rect 19701 6898 19767 6901
rect 31017 6898 31083 6901
rect 19701 6896 31083 6898
rect 19701 6840 19706 6896
rect 19762 6840 31022 6896
rect 31078 6840 31083 6896
rect 19701 6838 31083 6840
rect 19701 6835 19767 6838
rect 31017 6835 31083 6838
rect 12249 6762 12315 6765
rect 14222 6762 14228 6764
rect 12249 6760 14228 6762
rect 12249 6704 12254 6760
rect 12310 6704 14228 6760
rect 12249 6702 14228 6704
rect 12249 6699 12315 6702
rect 14222 6700 14228 6702
rect 14292 6700 14298 6764
rect 17585 6762 17651 6765
rect 17585 6760 20178 6762
rect 17585 6704 17590 6760
rect 17646 6704 20178 6760
rect 17585 6702 20178 6704
rect 17585 6699 17651 6702
rect 20118 6626 20178 6702
rect 22829 6626 22895 6629
rect 20118 6624 22895 6626
rect 20118 6568 22834 6624
rect 22890 6568 22895 6624
rect 20118 6566 22895 6568
rect 22829 6563 22895 6566
rect 4246 6560 4562 6561
rect 4246 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4562 6560
rect 4246 6495 4562 6496
rect 11951 6560 12267 6561
rect 11951 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12267 6560
rect 11951 6495 12267 6496
rect 19656 6560 19972 6561
rect 19656 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19972 6560
rect 19656 6495 19972 6496
rect 27361 6560 27677 6561
rect 27361 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27677 6560
rect 27361 6495 27677 6496
rect 13997 6490 14063 6493
rect 17953 6490 18019 6493
rect 13997 6488 18019 6490
rect 13997 6432 14002 6488
rect 14058 6432 17958 6488
rect 18014 6432 18019 6488
rect 13997 6430 18019 6432
rect 13997 6427 14063 6430
rect 17953 6427 18019 6430
rect 13077 6354 13143 6357
rect 15142 6354 15148 6356
rect 13077 6352 15148 6354
rect 13077 6296 13082 6352
rect 13138 6296 15148 6352
rect 13077 6294 15148 6296
rect 13077 6291 13143 6294
rect 15142 6292 15148 6294
rect 15212 6292 15218 6356
rect 4613 6218 4679 6221
rect 12525 6218 12591 6221
rect 4613 6216 12591 6218
rect 4613 6160 4618 6216
rect 4674 6160 12530 6216
rect 12586 6160 12591 6216
rect 4613 6158 12591 6160
rect 4613 6155 4679 6158
rect 12525 6155 12591 6158
rect 14457 6218 14523 6221
rect 14774 6218 14780 6220
rect 14457 6216 14780 6218
rect 14457 6160 14462 6216
rect 14518 6160 14780 6216
rect 14457 6158 14780 6160
rect 14457 6155 14523 6158
rect 14774 6156 14780 6158
rect 14844 6156 14850 6220
rect 17861 6218 17927 6221
rect 18454 6218 18460 6220
rect 17861 6216 18460 6218
rect 17861 6160 17866 6216
rect 17922 6160 18460 6216
rect 17861 6158 18460 6160
rect 17861 6155 17927 6158
rect 18454 6156 18460 6158
rect 18524 6218 18530 6220
rect 18873 6218 18939 6221
rect 18524 6216 18939 6218
rect 18524 6160 18878 6216
rect 18934 6160 18939 6216
rect 18524 6158 18939 6160
rect 18524 6156 18530 6158
rect 18873 6155 18939 6158
rect 8098 6016 8414 6017
rect 8098 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8414 6016
rect 8098 5951 8414 5952
rect 15803 6016 16119 6017
rect 15803 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16119 6016
rect 15803 5951 16119 5952
rect 23508 6016 23824 6017
rect 23508 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23824 6016
rect 23508 5951 23824 5952
rect 31213 6016 31529 6017
rect 31213 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31529 6016
rect 31213 5951 31529 5952
rect 11605 5946 11671 5949
rect 14365 5946 14431 5949
rect 11605 5944 14431 5946
rect 11605 5888 11610 5944
rect 11666 5888 14370 5944
rect 14426 5888 14431 5944
rect 11605 5886 14431 5888
rect 11605 5883 11671 5886
rect 14365 5883 14431 5886
rect 19885 5946 19951 5949
rect 22921 5946 22987 5949
rect 19885 5944 22987 5946
rect 19885 5888 19890 5944
rect 19946 5888 22926 5944
rect 22982 5888 22987 5944
rect 19885 5886 22987 5888
rect 19885 5883 19951 5886
rect 22921 5883 22987 5886
rect 19885 5810 19951 5813
rect 19885 5808 22110 5810
rect 19885 5752 19890 5808
rect 19946 5752 22110 5808
rect 19885 5750 22110 5752
rect 19885 5747 19951 5750
rect 19333 5674 19399 5677
rect 19609 5674 19675 5677
rect 19333 5672 19675 5674
rect 19333 5616 19338 5672
rect 19394 5616 19614 5672
rect 19670 5616 19675 5672
rect 19333 5614 19675 5616
rect 22050 5674 22110 5750
rect 29361 5674 29427 5677
rect 22050 5672 29427 5674
rect 22050 5616 29366 5672
rect 29422 5616 29427 5672
rect 22050 5614 29427 5616
rect 19333 5611 19399 5614
rect 19609 5611 19675 5614
rect 29361 5611 29427 5614
rect 4246 5472 4562 5473
rect 4246 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4562 5472
rect 4246 5407 4562 5408
rect 11951 5472 12267 5473
rect 11951 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12267 5472
rect 11951 5407 12267 5408
rect 19656 5472 19972 5473
rect 19656 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19972 5472
rect 19656 5407 19972 5408
rect 27361 5472 27677 5473
rect 27361 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27677 5472
rect 27361 5407 27677 5408
rect 9213 5402 9279 5405
rect 10409 5402 10475 5405
rect 9213 5400 10475 5402
rect 9213 5344 9218 5400
rect 9274 5344 10414 5400
rect 10470 5344 10475 5400
rect 9213 5342 10475 5344
rect 9213 5339 9279 5342
rect 10409 5339 10475 5342
rect 15929 5402 15995 5405
rect 16246 5402 16252 5404
rect 15929 5400 16252 5402
rect 15929 5344 15934 5400
rect 15990 5344 16252 5400
rect 15929 5342 16252 5344
rect 15929 5339 15995 5342
rect 16246 5340 16252 5342
rect 16316 5340 16322 5404
rect 15285 5266 15351 5269
rect 20713 5266 20779 5269
rect 15285 5264 20779 5266
rect 15285 5208 15290 5264
rect 15346 5208 20718 5264
rect 20774 5208 20779 5264
rect 15285 5206 20779 5208
rect 15285 5203 15351 5206
rect 20713 5203 20779 5206
rect 13629 5130 13695 5133
rect 22737 5130 22803 5133
rect 13629 5128 22803 5130
rect 13629 5072 13634 5128
rect 13690 5072 22742 5128
rect 22798 5072 22803 5128
rect 13629 5070 22803 5072
rect 13629 5067 13695 5070
rect 22737 5067 22803 5070
rect 8098 4928 8414 4929
rect 8098 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8414 4928
rect 8098 4863 8414 4864
rect 15803 4928 16119 4929
rect 15803 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16119 4928
rect 15803 4863 16119 4864
rect 23508 4928 23824 4929
rect 23508 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23824 4928
rect 23508 4863 23824 4864
rect 31213 4928 31529 4929
rect 31213 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31529 4928
rect 31213 4863 31529 4864
rect 7189 4722 7255 4725
rect 18965 4722 19031 4725
rect 7189 4720 19031 4722
rect 7189 4664 7194 4720
rect 7250 4664 18970 4720
rect 19026 4664 19031 4720
rect 7189 4662 19031 4664
rect 7189 4659 7255 4662
rect 18965 4659 19031 4662
rect 4889 4586 4955 4589
rect 18045 4586 18111 4589
rect 4889 4584 18111 4586
rect 4889 4528 4894 4584
rect 4950 4528 18050 4584
rect 18106 4528 18111 4584
rect 4889 4526 18111 4528
rect 4889 4523 4955 4526
rect 18045 4523 18111 4526
rect 19057 4586 19123 4589
rect 21633 4586 21699 4589
rect 23013 4586 23079 4589
rect 19057 4584 23079 4586
rect 19057 4528 19062 4584
rect 19118 4528 21638 4584
rect 21694 4528 23018 4584
rect 23074 4528 23079 4584
rect 19057 4526 23079 4528
rect 19057 4523 19123 4526
rect 21633 4523 21699 4526
rect 23013 4523 23079 4526
rect 13261 4450 13327 4453
rect 15510 4450 15516 4452
rect 13261 4448 15516 4450
rect 13261 4392 13266 4448
rect 13322 4392 15516 4448
rect 13261 4390 15516 4392
rect 13261 4387 13327 4390
rect 15510 4388 15516 4390
rect 15580 4450 15586 4452
rect 15837 4450 15903 4453
rect 15580 4448 15903 4450
rect 15580 4392 15842 4448
rect 15898 4392 15903 4448
rect 15580 4390 15903 4392
rect 15580 4388 15586 4390
rect 15837 4387 15903 4390
rect 17902 4388 17908 4452
rect 17972 4450 17978 4452
rect 18873 4450 18939 4453
rect 17972 4448 18939 4450
rect 17972 4392 18878 4448
rect 18934 4392 18939 4448
rect 17972 4390 18939 4392
rect 17972 4388 17978 4390
rect 18873 4387 18939 4390
rect 4246 4384 4562 4385
rect 4246 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4562 4384
rect 4246 4319 4562 4320
rect 11951 4384 12267 4385
rect 11951 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12267 4384
rect 11951 4319 12267 4320
rect 19656 4384 19972 4385
rect 19656 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19972 4384
rect 19656 4319 19972 4320
rect 27361 4384 27677 4385
rect 27361 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27677 4384
rect 27361 4319 27677 4320
rect 15561 4314 15627 4317
rect 16941 4314 17007 4317
rect 15561 4312 17007 4314
rect 15561 4256 15566 4312
rect 15622 4256 16946 4312
rect 17002 4256 17007 4312
rect 15561 4254 17007 4256
rect 15561 4251 15627 4254
rect 16941 4251 17007 4254
rect 14641 4178 14707 4181
rect 15561 4178 15627 4181
rect 14641 4176 15627 4178
rect 14641 4120 14646 4176
rect 14702 4120 15566 4176
rect 15622 4120 15627 4176
rect 14641 4118 15627 4120
rect 14641 4115 14707 4118
rect 15561 4115 15627 4118
rect 13670 3980 13676 4044
rect 13740 4042 13746 4044
rect 16573 4042 16639 4045
rect 13740 4040 16639 4042
rect 13740 3984 16578 4040
rect 16634 3984 16639 4040
rect 13740 3982 16639 3984
rect 13740 3980 13746 3982
rect 16573 3979 16639 3982
rect 22921 4042 22987 4045
rect 26601 4042 26667 4045
rect 22921 4040 26667 4042
rect 22921 3984 22926 4040
rect 22982 3984 26606 4040
rect 26662 3984 26667 4040
rect 22921 3982 26667 3984
rect 22921 3979 22987 3982
rect 26601 3979 26667 3982
rect 8098 3840 8414 3841
rect 8098 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8414 3840
rect 8098 3775 8414 3776
rect 15803 3840 16119 3841
rect 15803 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16119 3840
rect 15803 3775 16119 3776
rect 23508 3840 23824 3841
rect 23508 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23824 3840
rect 23508 3775 23824 3776
rect 31213 3840 31529 3841
rect 31213 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31529 3840
rect 31213 3775 31529 3776
rect 11973 3770 12039 3773
rect 14273 3770 14339 3773
rect 11973 3768 14339 3770
rect 11973 3712 11978 3768
rect 12034 3712 14278 3768
rect 14334 3712 14339 3768
rect 11973 3710 14339 3712
rect 11973 3707 12039 3710
rect 14273 3707 14339 3710
rect 12525 3634 12591 3637
rect 17217 3634 17283 3637
rect 12525 3632 17283 3634
rect 12525 3576 12530 3632
rect 12586 3576 17222 3632
rect 17278 3576 17283 3632
rect 12525 3574 17283 3576
rect 12525 3571 12591 3574
rect 17217 3571 17283 3574
rect 19057 3498 19123 3501
rect 20713 3498 20779 3501
rect 19057 3496 20779 3498
rect 19057 3440 19062 3496
rect 19118 3440 20718 3496
rect 20774 3440 20779 3496
rect 19057 3438 20779 3440
rect 19057 3435 19123 3438
rect 20713 3435 20779 3438
rect 4246 3296 4562 3297
rect 4246 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4562 3296
rect 4246 3231 4562 3232
rect 11951 3296 12267 3297
rect 11951 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12267 3296
rect 11951 3231 12267 3232
rect 19656 3296 19972 3297
rect 19656 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19972 3296
rect 19656 3231 19972 3232
rect 27361 3296 27677 3297
rect 27361 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27677 3296
rect 27361 3231 27677 3232
rect 5257 2954 5323 2957
rect 14958 2954 14964 2956
rect 5257 2952 14964 2954
rect 5257 2896 5262 2952
rect 5318 2896 14964 2952
rect 5257 2894 14964 2896
rect 5257 2891 5323 2894
rect 14958 2892 14964 2894
rect 15028 2892 15034 2956
rect 31600 2816 32000 2848
rect 31600 2760 31666 2816
rect 31722 2760 32000 2816
rect 8098 2752 8414 2753
rect 8098 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8414 2752
rect 8098 2687 8414 2688
rect 15803 2752 16119 2753
rect 15803 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16119 2752
rect 15803 2687 16119 2688
rect 23508 2752 23824 2753
rect 23508 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23824 2752
rect 23508 2687 23824 2688
rect 31213 2752 31529 2753
rect 31213 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31529 2752
rect 31600 2728 32000 2760
rect 31213 2687 31529 2688
rect 4246 2208 4562 2209
rect 4246 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4562 2208
rect 4246 2143 4562 2144
rect 11951 2208 12267 2209
rect 11951 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12267 2208
rect 11951 2143 12267 2144
rect 19656 2208 19972 2209
rect 19656 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19972 2208
rect 19656 2143 19972 2144
rect 27361 2208 27677 2209
rect 27361 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27677 2208
rect 27361 2143 27677 2144
rect 31017 2138 31083 2141
rect 31600 2138 32000 2168
rect 31017 2136 32000 2138
rect 31017 2080 31022 2136
rect 31078 2080 32000 2136
rect 31017 2078 32000 2080
rect 31017 2075 31083 2078
rect 31600 2048 32000 2078
rect 8098 1664 8414 1665
rect 8098 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8414 1664
rect 8098 1599 8414 1600
rect 15803 1664 16119 1665
rect 15803 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16119 1664
rect 15803 1599 16119 1600
rect 23508 1664 23824 1665
rect 23508 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23824 1664
rect 23508 1599 23824 1600
rect 31213 1664 31529 1665
rect 31213 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31529 1664
rect 31213 1599 31529 1600
rect 31017 1458 31083 1461
rect 31600 1458 32000 1488
rect 31017 1456 32000 1458
rect 31017 1400 31022 1456
rect 31078 1400 32000 1456
rect 31017 1398 32000 1400
rect 31017 1395 31083 1398
rect 31600 1368 32000 1398
rect 4246 1120 4562 1121
rect 4246 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4562 1120
rect 4246 1055 4562 1056
rect 11951 1120 12267 1121
rect 11951 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12267 1120
rect 11951 1055 12267 1056
rect 19656 1120 19972 1121
rect 19656 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19972 1120
rect 19656 1055 19972 1056
rect 27361 1120 27677 1121
rect 27361 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27677 1120
rect 27361 1055 27677 1056
rect 31017 778 31083 781
rect 31600 778 32000 808
rect 31017 776 32000 778
rect 31017 720 31022 776
rect 31078 720 32000 776
rect 31017 718 32000 720
rect 31017 715 31083 718
rect 31600 688 32000 718
rect 8098 576 8414 577
rect 8098 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8414 576
rect 8098 511 8414 512
rect 15803 576 16119 577
rect 15803 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16119 576
rect 15803 511 16119 512
rect 23508 576 23824 577
rect 23508 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23824 576
rect 23508 511 23824 512
rect 31213 576 31529 577
rect 31213 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31529 576
rect 31213 511 31529 512
<< via3 >>
rect 8104 19068 8168 19072
rect 8104 19012 8108 19068
rect 8108 19012 8164 19068
rect 8164 19012 8168 19068
rect 8104 19008 8168 19012
rect 8184 19068 8248 19072
rect 8184 19012 8188 19068
rect 8188 19012 8244 19068
rect 8244 19012 8248 19068
rect 8184 19008 8248 19012
rect 8264 19068 8328 19072
rect 8264 19012 8268 19068
rect 8268 19012 8324 19068
rect 8324 19012 8328 19068
rect 8264 19008 8328 19012
rect 8344 19068 8408 19072
rect 8344 19012 8348 19068
rect 8348 19012 8404 19068
rect 8404 19012 8408 19068
rect 8344 19008 8408 19012
rect 15809 19068 15873 19072
rect 15809 19012 15813 19068
rect 15813 19012 15869 19068
rect 15869 19012 15873 19068
rect 15809 19008 15873 19012
rect 15889 19068 15953 19072
rect 15889 19012 15893 19068
rect 15893 19012 15949 19068
rect 15949 19012 15953 19068
rect 15889 19008 15953 19012
rect 15969 19068 16033 19072
rect 15969 19012 15973 19068
rect 15973 19012 16029 19068
rect 16029 19012 16033 19068
rect 15969 19008 16033 19012
rect 16049 19068 16113 19072
rect 16049 19012 16053 19068
rect 16053 19012 16109 19068
rect 16109 19012 16113 19068
rect 16049 19008 16113 19012
rect 23514 19068 23578 19072
rect 23514 19012 23518 19068
rect 23518 19012 23574 19068
rect 23574 19012 23578 19068
rect 23514 19008 23578 19012
rect 23594 19068 23658 19072
rect 23594 19012 23598 19068
rect 23598 19012 23654 19068
rect 23654 19012 23658 19068
rect 23594 19008 23658 19012
rect 23674 19068 23738 19072
rect 23674 19012 23678 19068
rect 23678 19012 23734 19068
rect 23734 19012 23738 19068
rect 23674 19008 23738 19012
rect 23754 19068 23818 19072
rect 23754 19012 23758 19068
rect 23758 19012 23814 19068
rect 23814 19012 23818 19068
rect 23754 19008 23818 19012
rect 31219 19068 31283 19072
rect 31219 19012 31223 19068
rect 31223 19012 31279 19068
rect 31279 19012 31283 19068
rect 31219 19008 31283 19012
rect 31299 19068 31363 19072
rect 31299 19012 31303 19068
rect 31303 19012 31359 19068
rect 31359 19012 31363 19068
rect 31299 19008 31363 19012
rect 31379 19068 31443 19072
rect 31379 19012 31383 19068
rect 31383 19012 31439 19068
rect 31439 19012 31443 19068
rect 31379 19008 31443 19012
rect 31459 19068 31523 19072
rect 31459 19012 31463 19068
rect 31463 19012 31519 19068
rect 31519 19012 31523 19068
rect 31459 19008 31523 19012
rect 4252 18524 4316 18528
rect 4252 18468 4256 18524
rect 4256 18468 4312 18524
rect 4312 18468 4316 18524
rect 4252 18464 4316 18468
rect 4332 18524 4396 18528
rect 4332 18468 4336 18524
rect 4336 18468 4392 18524
rect 4392 18468 4396 18524
rect 4332 18464 4396 18468
rect 4412 18524 4476 18528
rect 4412 18468 4416 18524
rect 4416 18468 4472 18524
rect 4472 18468 4476 18524
rect 4412 18464 4476 18468
rect 4492 18524 4556 18528
rect 4492 18468 4496 18524
rect 4496 18468 4552 18524
rect 4552 18468 4556 18524
rect 4492 18464 4556 18468
rect 11957 18524 12021 18528
rect 11957 18468 11961 18524
rect 11961 18468 12017 18524
rect 12017 18468 12021 18524
rect 11957 18464 12021 18468
rect 12037 18524 12101 18528
rect 12037 18468 12041 18524
rect 12041 18468 12097 18524
rect 12097 18468 12101 18524
rect 12037 18464 12101 18468
rect 12117 18524 12181 18528
rect 12117 18468 12121 18524
rect 12121 18468 12177 18524
rect 12177 18468 12181 18524
rect 12117 18464 12181 18468
rect 12197 18524 12261 18528
rect 12197 18468 12201 18524
rect 12201 18468 12257 18524
rect 12257 18468 12261 18524
rect 12197 18464 12261 18468
rect 19662 18524 19726 18528
rect 19662 18468 19666 18524
rect 19666 18468 19722 18524
rect 19722 18468 19726 18524
rect 19662 18464 19726 18468
rect 19742 18524 19806 18528
rect 19742 18468 19746 18524
rect 19746 18468 19802 18524
rect 19802 18468 19806 18524
rect 19742 18464 19806 18468
rect 19822 18524 19886 18528
rect 19822 18468 19826 18524
rect 19826 18468 19882 18524
rect 19882 18468 19886 18524
rect 19822 18464 19886 18468
rect 19902 18524 19966 18528
rect 19902 18468 19906 18524
rect 19906 18468 19962 18524
rect 19962 18468 19966 18524
rect 19902 18464 19966 18468
rect 27367 18524 27431 18528
rect 27367 18468 27371 18524
rect 27371 18468 27427 18524
rect 27427 18468 27431 18524
rect 27367 18464 27431 18468
rect 27447 18524 27511 18528
rect 27447 18468 27451 18524
rect 27451 18468 27507 18524
rect 27507 18468 27511 18524
rect 27447 18464 27511 18468
rect 27527 18524 27591 18528
rect 27527 18468 27531 18524
rect 27531 18468 27587 18524
rect 27587 18468 27591 18524
rect 27527 18464 27591 18468
rect 27607 18524 27671 18528
rect 27607 18468 27611 18524
rect 27611 18468 27667 18524
rect 27667 18468 27671 18524
rect 27607 18464 27671 18468
rect 14964 18048 15028 18052
rect 14964 17992 15014 18048
rect 15014 17992 15028 18048
rect 14964 17988 15028 17992
rect 8104 17980 8168 17984
rect 8104 17924 8108 17980
rect 8108 17924 8164 17980
rect 8164 17924 8168 17980
rect 8104 17920 8168 17924
rect 8184 17980 8248 17984
rect 8184 17924 8188 17980
rect 8188 17924 8244 17980
rect 8244 17924 8248 17980
rect 8184 17920 8248 17924
rect 8264 17980 8328 17984
rect 8264 17924 8268 17980
rect 8268 17924 8324 17980
rect 8324 17924 8328 17980
rect 8264 17920 8328 17924
rect 8344 17980 8408 17984
rect 8344 17924 8348 17980
rect 8348 17924 8404 17980
rect 8404 17924 8408 17980
rect 8344 17920 8408 17924
rect 15809 17980 15873 17984
rect 15809 17924 15813 17980
rect 15813 17924 15869 17980
rect 15869 17924 15873 17980
rect 15809 17920 15873 17924
rect 15889 17980 15953 17984
rect 15889 17924 15893 17980
rect 15893 17924 15949 17980
rect 15949 17924 15953 17980
rect 15889 17920 15953 17924
rect 15969 17980 16033 17984
rect 15969 17924 15973 17980
rect 15973 17924 16029 17980
rect 16029 17924 16033 17980
rect 15969 17920 16033 17924
rect 16049 17980 16113 17984
rect 16049 17924 16053 17980
rect 16053 17924 16109 17980
rect 16109 17924 16113 17980
rect 16049 17920 16113 17924
rect 23514 17980 23578 17984
rect 23514 17924 23518 17980
rect 23518 17924 23574 17980
rect 23574 17924 23578 17980
rect 23514 17920 23578 17924
rect 23594 17980 23658 17984
rect 23594 17924 23598 17980
rect 23598 17924 23654 17980
rect 23654 17924 23658 17980
rect 23594 17920 23658 17924
rect 23674 17980 23738 17984
rect 23674 17924 23678 17980
rect 23678 17924 23734 17980
rect 23734 17924 23738 17980
rect 23674 17920 23738 17924
rect 23754 17980 23818 17984
rect 23754 17924 23758 17980
rect 23758 17924 23814 17980
rect 23814 17924 23818 17980
rect 23754 17920 23818 17924
rect 31219 17980 31283 17984
rect 31219 17924 31223 17980
rect 31223 17924 31279 17980
rect 31279 17924 31283 17980
rect 31219 17920 31283 17924
rect 31299 17980 31363 17984
rect 31299 17924 31303 17980
rect 31303 17924 31359 17980
rect 31359 17924 31363 17980
rect 31299 17920 31363 17924
rect 31379 17980 31443 17984
rect 31379 17924 31383 17980
rect 31383 17924 31439 17980
rect 31439 17924 31443 17980
rect 31379 17920 31443 17924
rect 31459 17980 31523 17984
rect 31459 17924 31463 17980
rect 31463 17924 31519 17980
rect 31519 17924 31523 17980
rect 31459 17920 31523 17924
rect 4252 17436 4316 17440
rect 4252 17380 4256 17436
rect 4256 17380 4312 17436
rect 4312 17380 4316 17436
rect 4252 17376 4316 17380
rect 4332 17436 4396 17440
rect 4332 17380 4336 17436
rect 4336 17380 4392 17436
rect 4392 17380 4396 17436
rect 4332 17376 4396 17380
rect 4412 17436 4476 17440
rect 4412 17380 4416 17436
rect 4416 17380 4472 17436
rect 4472 17380 4476 17436
rect 4412 17376 4476 17380
rect 4492 17436 4556 17440
rect 4492 17380 4496 17436
rect 4496 17380 4552 17436
rect 4552 17380 4556 17436
rect 4492 17376 4556 17380
rect 11957 17436 12021 17440
rect 11957 17380 11961 17436
rect 11961 17380 12017 17436
rect 12017 17380 12021 17436
rect 11957 17376 12021 17380
rect 12037 17436 12101 17440
rect 12037 17380 12041 17436
rect 12041 17380 12097 17436
rect 12097 17380 12101 17436
rect 12037 17376 12101 17380
rect 12117 17436 12181 17440
rect 12117 17380 12121 17436
rect 12121 17380 12177 17436
rect 12177 17380 12181 17436
rect 12117 17376 12181 17380
rect 12197 17436 12261 17440
rect 12197 17380 12201 17436
rect 12201 17380 12257 17436
rect 12257 17380 12261 17436
rect 12197 17376 12261 17380
rect 19662 17436 19726 17440
rect 19662 17380 19666 17436
rect 19666 17380 19722 17436
rect 19722 17380 19726 17436
rect 19662 17376 19726 17380
rect 19742 17436 19806 17440
rect 19742 17380 19746 17436
rect 19746 17380 19802 17436
rect 19802 17380 19806 17436
rect 19742 17376 19806 17380
rect 19822 17436 19886 17440
rect 19822 17380 19826 17436
rect 19826 17380 19882 17436
rect 19882 17380 19886 17436
rect 19822 17376 19886 17380
rect 19902 17436 19966 17440
rect 19902 17380 19906 17436
rect 19906 17380 19962 17436
rect 19962 17380 19966 17436
rect 19902 17376 19966 17380
rect 27367 17436 27431 17440
rect 27367 17380 27371 17436
rect 27371 17380 27427 17436
rect 27427 17380 27431 17436
rect 27367 17376 27431 17380
rect 27447 17436 27511 17440
rect 27447 17380 27451 17436
rect 27451 17380 27507 17436
rect 27507 17380 27511 17436
rect 27447 17376 27511 17380
rect 27527 17436 27591 17440
rect 27527 17380 27531 17436
rect 27531 17380 27587 17436
rect 27587 17380 27591 17436
rect 27527 17376 27591 17380
rect 27607 17436 27671 17440
rect 27607 17380 27611 17436
rect 27611 17380 27667 17436
rect 27667 17380 27671 17436
rect 27607 17376 27671 17380
rect 8104 16892 8168 16896
rect 8104 16836 8108 16892
rect 8108 16836 8164 16892
rect 8164 16836 8168 16892
rect 8104 16832 8168 16836
rect 8184 16892 8248 16896
rect 8184 16836 8188 16892
rect 8188 16836 8244 16892
rect 8244 16836 8248 16892
rect 8184 16832 8248 16836
rect 8264 16892 8328 16896
rect 8264 16836 8268 16892
rect 8268 16836 8324 16892
rect 8324 16836 8328 16892
rect 8264 16832 8328 16836
rect 8344 16892 8408 16896
rect 8344 16836 8348 16892
rect 8348 16836 8404 16892
rect 8404 16836 8408 16892
rect 8344 16832 8408 16836
rect 15809 16892 15873 16896
rect 15809 16836 15813 16892
rect 15813 16836 15869 16892
rect 15869 16836 15873 16892
rect 15809 16832 15873 16836
rect 15889 16892 15953 16896
rect 15889 16836 15893 16892
rect 15893 16836 15949 16892
rect 15949 16836 15953 16892
rect 15889 16832 15953 16836
rect 15969 16892 16033 16896
rect 15969 16836 15973 16892
rect 15973 16836 16029 16892
rect 16029 16836 16033 16892
rect 15969 16832 16033 16836
rect 16049 16892 16113 16896
rect 16049 16836 16053 16892
rect 16053 16836 16109 16892
rect 16109 16836 16113 16892
rect 16049 16832 16113 16836
rect 23514 16892 23578 16896
rect 23514 16836 23518 16892
rect 23518 16836 23574 16892
rect 23574 16836 23578 16892
rect 23514 16832 23578 16836
rect 23594 16892 23658 16896
rect 23594 16836 23598 16892
rect 23598 16836 23654 16892
rect 23654 16836 23658 16892
rect 23594 16832 23658 16836
rect 23674 16892 23738 16896
rect 23674 16836 23678 16892
rect 23678 16836 23734 16892
rect 23734 16836 23738 16892
rect 23674 16832 23738 16836
rect 23754 16892 23818 16896
rect 23754 16836 23758 16892
rect 23758 16836 23814 16892
rect 23814 16836 23818 16892
rect 23754 16832 23818 16836
rect 31219 16892 31283 16896
rect 31219 16836 31223 16892
rect 31223 16836 31279 16892
rect 31279 16836 31283 16892
rect 31219 16832 31283 16836
rect 31299 16892 31363 16896
rect 31299 16836 31303 16892
rect 31303 16836 31359 16892
rect 31359 16836 31363 16892
rect 31299 16832 31363 16836
rect 31379 16892 31443 16896
rect 31379 16836 31383 16892
rect 31383 16836 31439 16892
rect 31439 16836 31443 16892
rect 31379 16832 31443 16836
rect 31459 16892 31523 16896
rect 31459 16836 31463 16892
rect 31463 16836 31519 16892
rect 31519 16836 31523 16892
rect 31459 16832 31523 16836
rect 18828 16628 18892 16692
rect 4252 16348 4316 16352
rect 4252 16292 4256 16348
rect 4256 16292 4312 16348
rect 4312 16292 4316 16348
rect 4252 16288 4316 16292
rect 4332 16348 4396 16352
rect 4332 16292 4336 16348
rect 4336 16292 4392 16348
rect 4392 16292 4396 16348
rect 4332 16288 4396 16292
rect 4412 16348 4476 16352
rect 4412 16292 4416 16348
rect 4416 16292 4472 16348
rect 4472 16292 4476 16348
rect 4412 16288 4476 16292
rect 4492 16348 4556 16352
rect 4492 16292 4496 16348
rect 4496 16292 4552 16348
rect 4552 16292 4556 16348
rect 4492 16288 4556 16292
rect 11957 16348 12021 16352
rect 11957 16292 11961 16348
rect 11961 16292 12017 16348
rect 12017 16292 12021 16348
rect 11957 16288 12021 16292
rect 12037 16348 12101 16352
rect 12037 16292 12041 16348
rect 12041 16292 12097 16348
rect 12097 16292 12101 16348
rect 12037 16288 12101 16292
rect 12117 16348 12181 16352
rect 12117 16292 12121 16348
rect 12121 16292 12177 16348
rect 12177 16292 12181 16348
rect 12117 16288 12181 16292
rect 12197 16348 12261 16352
rect 12197 16292 12201 16348
rect 12201 16292 12257 16348
rect 12257 16292 12261 16348
rect 12197 16288 12261 16292
rect 19662 16348 19726 16352
rect 19662 16292 19666 16348
rect 19666 16292 19722 16348
rect 19722 16292 19726 16348
rect 19662 16288 19726 16292
rect 19742 16348 19806 16352
rect 19742 16292 19746 16348
rect 19746 16292 19802 16348
rect 19802 16292 19806 16348
rect 19742 16288 19806 16292
rect 19822 16348 19886 16352
rect 19822 16292 19826 16348
rect 19826 16292 19882 16348
rect 19882 16292 19886 16348
rect 19822 16288 19886 16292
rect 19902 16348 19966 16352
rect 19902 16292 19906 16348
rect 19906 16292 19962 16348
rect 19962 16292 19966 16348
rect 19902 16288 19966 16292
rect 27367 16348 27431 16352
rect 27367 16292 27371 16348
rect 27371 16292 27427 16348
rect 27427 16292 27431 16348
rect 27367 16288 27431 16292
rect 27447 16348 27511 16352
rect 27447 16292 27451 16348
rect 27451 16292 27507 16348
rect 27507 16292 27511 16348
rect 27447 16288 27511 16292
rect 27527 16348 27591 16352
rect 27527 16292 27531 16348
rect 27531 16292 27587 16348
rect 27587 16292 27591 16348
rect 27527 16288 27591 16292
rect 27607 16348 27671 16352
rect 27607 16292 27611 16348
rect 27611 16292 27667 16348
rect 27667 16292 27671 16348
rect 27607 16288 27671 16292
rect 16620 15948 16684 16012
rect 8104 15804 8168 15808
rect 8104 15748 8108 15804
rect 8108 15748 8164 15804
rect 8164 15748 8168 15804
rect 8104 15744 8168 15748
rect 8184 15804 8248 15808
rect 8184 15748 8188 15804
rect 8188 15748 8244 15804
rect 8244 15748 8248 15804
rect 8184 15744 8248 15748
rect 8264 15804 8328 15808
rect 8264 15748 8268 15804
rect 8268 15748 8324 15804
rect 8324 15748 8328 15804
rect 8264 15744 8328 15748
rect 8344 15804 8408 15808
rect 8344 15748 8348 15804
rect 8348 15748 8404 15804
rect 8404 15748 8408 15804
rect 8344 15744 8408 15748
rect 15809 15804 15873 15808
rect 15809 15748 15813 15804
rect 15813 15748 15869 15804
rect 15869 15748 15873 15804
rect 15809 15744 15873 15748
rect 15889 15804 15953 15808
rect 15889 15748 15893 15804
rect 15893 15748 15949 15804
rect 15949 15748 15953 15804
rect 15889 15744 15953 15748
rect 15969 15804 16033 15808
rect 15969 15748 15973 15804
rect 15973 15748 16029 15804
rect 16029 15748 16033 15804
rect 15969 15744 16033 15748
rect 16049 15804 16113 15808
rect 16049 15748 16053 15804
rect 16053 15748 16109 15804
rect 16109 15748 16113 15804
rect 16049 15744 16113 15748
rect 23514 15804 23578 15808
rect 23514 15748 23518 15804
rect 23518 15748 23574 15804
rect 23574 15748 23578 15804
rect 23514 15744 23578 15748
rect 23594 15804 23658 15808
rect 23594 15748 23598 15804
rect 23598 15748 23654 15804
rect 23654 15748 23658 15804
rect 23594 15744 23658 15748
rect 23674 15804 23738 15808
rect 23674 15748 23678 15804
rect 23678 15748 23734 15804
rect 23734 15748 23738 15804
rect 23674 15744 23738 15748
rect 23754 15804 23818 15808
rect 23754 15748 23758 15804
rect 23758 15748 23814 15804
rect 23814 15748 23818 15804
rect 23754 15744 23818 15748
rect 31219 15804 31283 15808
rect 31219 15748 31223 15804
rect 31223 15748 31279 15804
rect 31279 15748 31283 15804
rect 31219 15744 31283 15748
rect 31299 15804 31363 15808
rect 31299 15748 31303 15804
rect 31303 15748 31359 15804
rect 31359 15748 31363 15804
rect 31299 15744 31363 15748
rect 31379 15804 31443 15808
rect 31379 15748 31383 15804
rect 31383 15748 31439 15804
rect 31439 15748 31443 15804
rect 31379 15744 31443 15748
rect 31459 15804 31523 15808
rect 31459 15748 31463 15804
rect 31463 15748 31519 15804
rect 31519 15748 31523 15804
rect 31459 15744 31523 15748
rect 4252 15260 4316 15264
rect 4252 15204 4256 15260
rect 4256 15204 4312 15260
rect 4312 15204 4316 15260
rect 4252 15200 4316 15204
rect 4332 15260 4396 15264
rect 4332 15204 4336 15260
rect 4336 15204 4392 15260
rect 4392 15204 4396 15260
rect 4332 15200 4396 15204
rect 4412 15260 4476 15264
rect 4412 15204 4416 15260
rect 4416 15204 4472 15260
rect 4472 15204 4476 15260
rect 4412 15200 4476 15204
rect 4492 15260 4556 15264
rect 4492 15204 4496 15260
rect 4496 15204 4552 15260
rect 4552 15204 4556 15260
rect 4492 15200 4556 15204
rect 11957 15260 12021 15264
rect 11957 15204 11961 15260
rect 11961 15204 12017 15260
rect 12017 15204 12021 15260
rect 11957 15200 12021 15204
rect 12037 15260 12101 15264
rect 12037 15204 12041 15260
rect 12041 15204 12097 15260
rect 12097 15204 12101 15260
rect 12037 15200 12101 15204
rect 12117 15260 12181 15264
rect 12117 15204 12121 15260
rect 12121 15204 12177 15260
rect 12177 15204 12181 15260
rect 12117 15200 12181 15204
rect 12197 15260 12261 15264
rect 12197 15204 12201 15260
rect 12201 15204 12257 15260
rect 12257 15204 12261 15260
rect 12197 15200 12261 15204
rect 19662 15260 19726 15264
rect 19662 15204 19666 15260
rect 19666 15204 19722 15260
rect 19722 15204 19726 15260
rect 19662 15200 19726 15204
rect 19742 15260 19806 15264
rect 19742 15204 19746 15260
rect 19746 15204 19802 15260
rect 19802 15204 19806 15260
rect 19742 15200 19806 15204
rect 19822 15260 19886 15264
rect 19822 15204 19826 15260
rect 19826 15204 19882 15260
rect 19882 15204 19886 15260
rect 19822 15200 19886 15204
rect 19902 15260 19966 15264
rect 19902 15204 19906 15260
rect 19906 15204 19962 15260
rect 19962 15204 19966 15260
rect 19902 15200 19966 15204
rect 27367 15260 27431 15264
rect 27367 15204 27371 15260
rect 27371 15204 27427 15260
rect 27427 15204 27431 15260
rect 27367 15200 27431 15204
rect 27447 15260 27511 15264
rect 27447 15204 27451 15260
rect 27451 15204 27507 15260
rect 27507 15204 27511 15260
rect 27447 15200 27511 15204
rect 27527 15260 27591 15264
rect 27527 15204 27531 15260
rect 27531 15204 27587 15260
rect 27587 15204 27591 15260
rect 27527 15200 27591 15204
rect 27607 15260 27671 15264
rect 27607 15204 27611 15260
rect 27611 15204 27667 15260
rect 27667 15204 27671 15260
rect 27607 15200 27671 15204
rect 8104 14716 8168 14720
rect 8104 14660 8108 14716
rect 8108 14660 8164 14716
rect 8164 14660 8168 14716
rect 8104 14656 8168 14660
rect 8184 14716 8248 14720
rect 8184 14660 8188 14716
rect 8188 14660 8244 14716
rect 8244 14660 8248 14716
rect 8184 14656 8248 14660
rect 8264 14716 8328 14720
rect 8264 14660 8268 14716
rect 8268 14660 8324 14716
rect 8324 14660 8328 14716
rect 8264 14656 8328 14660
rect 8344 14716 8408 14720
rect 8344 14660 8348 14716
rect 8348 14660 8404 14716
rect 8404 14660 8408 14716
rect 8344 14656 8408 14660
rect 15809 14716 15873 14720
rect 15809 14660 15813 14716
rect 15813 14660 15869 14716
rect 15869 14660 15873 14716
rect 15809 14656 15873 14660
rect 15889 14716 15953 14720
rect 15889 14660 15893 14716
rect 15893 14660 15949 14716
rect 15949 14660 15953 14716
rect 15889 14656 15953 14660
rect 15969 14716 16033 14720
rect 15969 14660 15973 14716
rect 15973 14660 16029 14716
rect 16029 14660 16033 14716
rect 15969 14656 16033 14660
rect 16049 14716 16113 14720
rect 16049 14660 16053 14716
rect 16053 14660 16109 14716
rect 16109 14660 16113 14716
rect 16049 14656 16113 14660
rect 23514 14716 23578 14720
rect 23514 14660 23518 14716
rect 23518 14660 23574 14716
rect 23574 14660 23578 14716
rect 23514 14656 23578 14660
rect 23594 14716 23658 14720
rect 23594 14660 23598 14716
rect 23598 14660 23654 14716
rect 23654 14660 23658 14716
rect 23594 14656 23658 14660
rect 23674 14716 23738 14720
rect 23674 14660 23678 14716
rect 23678 14660 23734 14716
rect 23734 14660 23738 14716
rect 23674 14656 23738 14660
rect 23754 14716 23818 14720
rect 23754 14660 23758 14716
rect 23758 14660 23814 14716
rect 23814 14660 23818 14716
rect 23754 14656 23818 14660
rect 31219 14716 31283 14720
rect 31219 14660 31223 14716
rect 31223 14660 31279 14716
rect 31279 14660 31283 14716
rect 31219 14656 31283 14660
rect 31299 14716 31363 14720
rect 31299 14660 31303 14716
rect 31303 14660 31359 14716
rect 31359 14660 31363 14716
rect 31299 14656 31363 14660
rect 31379 14716 31443 14720
rect 31379 14660 31383 14716
rect 31383 14660 31439 14716
rect 31439 14660 31443 14716
rect 31379 14656 31443 14660
rect 31459 14716 31523 14720
rect 31459 14660 31463 14716
rect 31463 14660 31519 14716
rect 31519 14660 31523 14716
rect 31459 14656 31523 14660
rect 16988 14588 17052 14652
rect 4252 14172 4316 14176
rect 4252 14116 4256 14172
rect 4256 14116 4312 14172
rect 4312 14116 4316 14172
rect 4252 14112 4316 14116
rect 4332 14172 4396 14176
rect 4332 14116 4336 14172
rect 4336 14116 4392 14172
rect 4392 14116 4396 14172
rect 4332 14112 4396 14116
rect 4412 14172 4476 14176
rect 4412 14116 4416 14172
rect 4416 14116 4472 14172
rect 4472 14116 4476 14172
rect 4412 14112 4476 14116
rect 4492 14172 4556 14176
rect 4492 14116 4496 14172
rect 4496 14116 4552 14172
rect 4552 14116 4556 14172
rect 4492 14112 4556 14116
rect 11957 14172 12021 14176
rect 11957 14116 11961 14172
rect 11961 14116 12017 14172
rect 12017 14116 12021 14172
rect 11957 14112 12021 14116
rect 12037 14172 12101 14176
rect 12037 14116 12041 14172
rect 12041 14116 12097 14172
rect 12097 14116 12101 14172
rect 12037 14112 12101 14116
rect 12117 14172 12181 14176
rect 12117 14116 12121 14172
rect 12121 14116 12177 14172
rect 12177 14116 12181 14172
rect 12117 14112 12181 14116
rect 12197 14172 12261 14176
rect 12197 14116 12201 14172
rect 12201 14116 12257 14172
rect 12257 14116 12261 14172
rect 12197 14112 12261 14116
rect 19662 14172 19726 14176
rect 19662 14116 19666 14172
rect 19666 14116 19722 14172
rect 19722 14116 19726 14172
rect 19662 14112 19726 14116
rect 19742 14172 19806 14176
rect 19742 14116 19746 14172
rect 19746 14116 19802 14172
rect 19802 14116 19806 14172
rect 19742 14112 19806 14116
rect 19822 14172 19886 14176
rect 19822 14116 19826 14172
rect 19826 14116 19882 14172
rect 19882 14116 19886 14172
rect 19822 14112 19886 14116
rect 19902 14172 19966 14176
rect 19902 14116 19906 14172
rect 19906 14116 19962 14172
rect 19962 14116 19966 14172
rect 19902 14112 19966 14116
rect 27367 14172 27431 14176
rect 27367 14116 27371 14172
rect 27371 14116 27427 14172
rect 27427 14116 27431 14172
rect 27367 14112 27431 14116
rect 27447 14172 27511 14176
rect 27447 14116 27451 14172
rect 27451 14116 27507 14172
rect 27507 14116 27511 14172
rect 27447 14112 27511 14116
rect 27527 14172 27591 14176
rect 27527 14116 27531 14172
rect 27531 14116 27587 14172
rect 27587 14116 27591 14172
rect 27527 14112 27591 14116
rect 27607 14172 27671 14176
rect 27607 14116 27611 14172
rect 27611 14116 27667 14172
rect 27667 14116 27671 14172
rect 27607 14112 27671 14116
rect 8104 13628 8168 13632
rect 8104 13572 8108 13628
rect 8108 13572 8164 13628
rect 8164 13572 8168 13628
rect 8104 13568 8168 13572
rect 8184 13628 8248 13632
rect 8184 13572 8188 13628
rect 8188 13572 8244 13628
rect 8244 13572 8248 13628
rect 8184 13568 8248 13572
rect 8264 13628 8328 13632
rect 8264 13572 8268 13628
rect 8268 13572 8324 13628
rect 8324 13572 8328 13628
rect 8264 13568 8328 13572
rect 8344 13628 8408 13632
rect 8344 13572 8348 13628
rect 8348 13572 8404 13628
rect 8404 13572 8408 13628
rect 8344 13568 8408 13572
rect 16804 13832 16868 13836
rect 16804 13776 16818 13832
rect 16818 13776 16868 13832
rect 16804 13772 16868 13776
rect 15809 13628 15873 13632
rect 15809 13572 15813 13628
rect 15813 13572 15869 13628
rect 15869 13572 15873 13628
rect 15809 13568 15873 13572
rect 15889 13628 15953 13632
rect 15889 13572 15893 13628
rect 15893 13572 15949 13628
rect 15949 13572 15953 13628
rect 15889 13568 15953 13572
rect 15969 13628 16033 13632
rect 15969 13572 15973 13628
rect 15973 13572 16029 13628
rect 16029 13572 16033 13628
rect 15969 13568 16033 13572
rect 16049 13628 16113 13632
rect 16049 13572 16053 13628
rect 16053 13572 16109 13628
rect 16109 13572 16113 13628
rect 16049 13568 16113 13572
rect 23514 13628 23578 13632
rect 23514 13572 23518 13628
rect 23518 13572 23574 13628
rect 23574 13572 23578 13628
rect 23514 13568 23578 13572
rect 23594 13628 23658 13632
rect 23594 13572 23598 13628
rect 23598 13572 23654 13628
rect 23654 13572 23658 13628
rect 23594 13568 23658 13572
rect 23674 13628 23738 13632
rect 23674 13572 23678 13628
rect 23678 13572 23734 13628
rect 23734 13572 23738 13628
rect 23674 13568 23738 13572
rect 23754 13628 23818 13632
rect 23754 13572 23758 13628
rect 23758 13572 23814 13628
rect 23814 13572 23818 13628
rect 23754 13568 23818 13572
rect 31219 13628 31283 13632
rect 31219 13572 31223 13628
rect 31223 13572 31279 13628
rect 31279 13572 31283 13628
rect 31219 13568 31283 13572
rect 31299 13628 31363 13632
rect 31299 13572 31303 13628
rect 31303 13572 31359 13628
rect 31359 13572 31363 13628
rect 31299 13568 31363 13572
rect 31379 13628 31443 13632
rect 31379 13572 31383 13628
rect 31383 13572 31439 13628
rect 31439 13572 31443 13628
rect 31379 13568 31443 13572
rect 31459 13628 31523 13632
rect 31459 13572 31463 13628
rect 31463 13572 31519 13628
rect 31519 13572 31523 13628
rect 31459 13568 31523 13572
rect 4252 13084 4316 13088
rect 4252 13028 4256 13084
rect 4256 13028 4312 13084
rect 4312 13028 4316 13084
rect 4252 13024 4316 13028
rect 4332 13084 4396 13088
rect 4332 13028 4336 13084
rect 4336 13028 4392 13084
rect 4392 13028 4396 13084
rect 4332 13024 4396 13028
rect 4412 13084 4476 13088
rect 4412 13028 4416 13084
rect 4416 13028 4472 13084
rect 4472 13028 4476 13084
rect 4412 13024 4476 13028
rect 4492 13084 4556 13088
rect 4492 13028 4496 13084
rect 4496 13028 4552 13084
rect 4552 13028 4556 13084
rect 4492 13024 4556 13028
rect 11957 13084 12021 13088
rect 11957 13028 11961 13084
rect 11961 13028 12017 13084
rect 12017 13028 12021 13084
rect 11957 13024 12021 13028
rect 12037 13084 12101 13088
rect 12037 13028 12041 13084
rect 12041 13028 12097 13084
rect 12097 13028 12101 13084
rect 12037 13024 12101 13028
rect 12117 13084 12181 13088
rect 12117 13028 12121 13084
rect 12121 13028 12177 13084
rect 12177 13028 12181 13084
rect 12117 13024 12181 13028
rect 12197 13084 12261 13088
rect 12197 13028 12201 13084
rect 12201 13028 12257 13084
rect 12257 13028 12261 13084
rect 12197 13024 12261 13028
rect 19662 13084 19726 13088
rect 19662 13028 19666 13084
rect 19666 13028 19722 13084
rect 19722 13028 19726 13084
rect 19662 13024 19726 13028
rect 19742 13084 19806 13088
rect 19742 13028 19746 13084
rect 19746 13028 19802 13084
rect 19802 13028 19806 13084
rect 19742 13024 19806 13028
rect 19822 13084 19886 13088
rect 19822 13028 19826 13084
rect 19826 13028 19882 13084
rect 19882 13028 19886 13084
rect 19822 13024 19886 13028
rect 19902 13084 19966 13088
rect 19902 13028 19906 13084
rect 19906 13028 19962 13084
rect 19962 13028 19966 13084
rect 19902 13024 19966 13028
rect 27367 13084 27431 13088
rect 27367 13028 27371 13084
rect 27371 13028 27427 13084
rect 27427 13028 27431 13084
rect 27367 13024 27431 13028
rect 27447 13084 27511 13088
rect 27447 13028 27451 13084
rect 27451 13028 27507 13084
rect 27507 13028 27511 13084
rect 27447 13024 27511 13028
rect 27527 13084 27591 13088
rect 27527 13028 27531 13084
rect 27531 13028 27587 13084
rect 27587 13028 27591 13084
rect 27527 13024 27591 13028
rect 27607 13084 27671 13088
rect 27607 13028 27611 13084
rect 27611 13028 27667 13084
rect 27667 13028 27671 13084
rect 27607 13024 27671 13028
rect 14412 12820 14476 12884
rect 19196 12956 19260 13020
rect 14044 12548 14108 12612
rect 8104 12540 8168 12544
rect 8104 12484 8108 12540
rect 8108 12484 8164 12540
rect 8164 12484 8168 12540
rect 8104 12480 8168 12484
rect 8184 12540 8248 12544
rect 8184 12484 8188 12540
rect 8188 12484 8244 12540
rect 8244 12484 8248 12540
rect 8184 12480 8248 12484
rect 8264 12540 8328 12544
rect 8264 12484 8268 12540
rect 8268 12484 8324 12540
rect 8324 12484 8328 12540
rect 8264 12480 8328 12484
rect 8344 12540 8408 12544
rect 8344 12484 8348 12540
rect 8348 12484 8404 12540
rect 8404 12484 8408 12540
rect 8344 12480 8408 12484
rect 15809 12540 15873 12544
rect 15809 12484 15813 12540
rect 15813 12484 15869 12540
rect 15869 12484 15873 12540
rect 15809 12480 15873 12484
rect 15889 12540 15953 12544
rect 15889 12484 15893 12540
rect 15893 12484 15949 12540
rect 15949 12484 15953 12540
rect 15889 12480 15953 12484
rect 15969 12540 16033 12544
rect 15969 12484 15973 12540
rect 15973 12484 16029 12540
rect 16029 12484 16033 12540
rect 15969 12480 16033 12484
rect 16049 12540 16113 12544
rect 16049 12484 16053 12540
rect 16053 12484 16109 12540
rect 16109 12484 16113 12540
rect 16049 12480 16113 12484
rect 23514 12540 23578 12544
rect 23514 12484 23518 12540
rect 23518 12484 23574 12540
rect 23574 12484 23578 12540
rect 23514 12480 23578 12484
rect 23594 12540 23658 12544
rect 23594 12484 23598 12540
rect 23598 12484 23654 12540
rect 23654 12484 23658 12540
rect 23594 12480 23658 12484
rect 23674 12540 23738 12544
rect 23674 12484 23678 12540
rect 23678 12484 23734 12540
rect 23734 12484 23738 12540
rect 23674 12480 23738 12484
rect 23754 12540 23818 12544
rect 23754 12484 23758 12540
rect 23758 12484 23814 12540
rect 23814 12484 23818 12540
rect 23754 12480 23818 12484
rect 31219 12540 31283 12544
rect 31219 12484 31223 12540
rect 31223 12484 31279 12540
rect 31279 12484 31283 12540
rect 31219 12480 31283 12484
rect 31299 12540 31363 12544
rect 31299 12484 31303 12540
rect 31303 12484 31359 12540
rect 31359 12484 31363 12540
rect 31299 12480 31363 12484
rect 31379 12540 31443 12544
rect 31379 12484 31383 12540
rect 31383 12484 31439 12540
rect 31439 12484 31443 12540
rect 31379 12480 31443 12484
rect 31459 12540 31523 12544
rect 31459 12484 31463 12540
rect 31463 12484 31519 12540
rect 31519 12484 31523 12540
rect 31459 12480 31523 12484
rect 4252 11996 4316 12000
rect 4252 11940 4256 11996
rect 4256 11940 4312 11996
rect 4312 11940 4316 11996
rect 4252 11936 4316 11940
rect 4332 11996 4396 12000
rect 4332 11940 4336 11996
rect 4336 11940 4392 11996
rect 4392 11940 4396 11996
rect 4332 11936 4396 11940
rect 4412 11996 4476 12000
rect 4412 11940 4416 11996
rect 4416 11940 4472 11996
rect 4472 11940 4476 11996
rect 4412 11936 4476 11940
rect 4492 11996 4556 12000
rect 4492 11940 4496 11996
rect 4496 11940 4552 11996
rect 4552 11940 4556 11996
rect 4492 11936 4556 11940
rect 11957 11996 12021 12000
rect 11957 11940 11961 11996
rect 11961 11940 12017 11996
rect 12017 11940 12021 11996
rect 11957 11936 12021 11940
rect 12037 11996 12101 12000
rect 12037 11940 12041 11996
rect 12041 11940 12097 11996
rect 12097 11940 12101 11996
rect 12037 11936 12101 11940
rect 12117 11996 12181 12000
rect 12117 11940 12121 11996
rect 12121 11940 12177 11996
rect 12177 11940 12181 11996
rect 12117 11936 12181 11940
rect 12197 11996 12261 12000
rect 12197 11940 12201 11996
rect 12201 11940 12257 11996
rect 12257 11940 12261 11996
rect 12197 11936 12261 11940
rect 19662 11996 19726 12000
rect 19662 11940 19666 11996
rect 19666 11940 19722 11996
rect 19722 11940 19726 11996
rect 19662 11936 19726 11940
rect 19742 11996 19806 12000
rect 19742 11940 19746 11996
rect 19746 11940 19802 11996
rect 19802 11940 19806 11996
rect 19742 11936 19806 11940
rect 19822 11996 19886 12000
rect 19822 11940 19826 11996
rect 19826 11940 19882 11996
rect 19882 11940 19886 11996
rect 19822 11936 19886 11940
rect 19902 11996 19966 12000
rect 19902 11940 19906 11996
rect 19906 11940 19962 11996
rect 19962 11940 19966 11996
rect 19902 11936 19966 11940
rect 27367 11996 27431 12000
rect 27367 11940 27371 11996
rect 27371 11940 27427 11996
rect 27427 11940 27431 11996
rect 27367 11936 27431 11940
rect 27447 11996 27511 12000
rect 27447 11940 27451 11996
rect 27451 11940 27507 11996
rect 27507 11940 27511 11996
rect 27447 11936 27511 11940
rect 27527 11996 27591 12000
rect 27527 11940 27531 11996
rect 27531 11940 27587 11996
rect 27587 11940 27591 11996
rect 27527 11936 27591 11940
rect 27607 11996 27671 12000
rect 27607 11940 27611 11996
rect 27611 11940 27667 11996
rect 27667 11940 27671 11996
rect 27607 11936 27671 11940
rect 17908 11732 17972 11796
rect 8104 11452 8168 11456
rect 8104 11396 8108 11452
rect 8108 11396 8164 11452
rect 8164 11396 8168 11452
rect 8104 11392 8168 11396
rect 8184 11452 8248 11456
rect 8184 11396 8188 11452
rect 8188 11396 8244 11452
rect 8244 11396 8248 11452
rect 8184 11392 8248 11396
rect 8264 11452 8328 11456
rect 8264 11396 8268 11452
rect 8268 11396 8324 11452
rect 8324 11396 8328 11452
rect 8264 11392 8328 11396
rect 8344 11452 8408 11456
rect 8344 11396 8348 11452
rect 8348 11396 8404 11452
rect 8404 11396 8408 11452
rect 8344 11392 8408 11396
rect 16804 11520 16868 11524
rect 16804 11464 16818 11520
rect 16818 11464 16868 11520
rect 16804 11460 16868 11464
rect 15809 11452 15873 11456
rect 15809 11396 15813 11452
rect 15813 11396 15869 11452
rect 15869 11396 15873 11452
rect 15809 11392 15873 11396
rect 15889 11452 15953 11456
rect 15889 11396 15893 11452
rect 15893 11396 15949 11452
rect 15949 11396 15953 11452
rect 15889 11392 15953 11396
rect 15969 11452 16033 11456
rect 15969 11396 15973 11452
rect 15973 11396 16029 11452
rect 16029 11396 16033 11452
rect 15969 11392 16033 11396
rect 16049 11452 16113 11456
rect 16049 11396 16053 11452
rect 16053 11396 16109 11452
rect 16109 11396 16113 11452
rect 16049 11392 16113 11396
rect 23514 11452 23578 11456
rect 23514 11396 23518 11452
rect 23518 11396 23574 11452
rect 23574 11396 23578 11452
rect 23514 11392 23578 11396
rect 23594 11452 23658 11456
rect 23594 11396 23598 11452
rect 23598 11396 23654 11452
rect 23654 11396 23658 11452
rect 23594 11392 23658 11396
rect 23674 11452 23738 11456
rect 23674 11396 23678 11452
rect 23678 11396 23734 11452
rect 23734 11396 23738 11452
rect 23674 11392 23738 11396
rect 23754 11452 23818 11456
rect 23754 11396 23758 11452
rect 23758 11396 23814 11452
rect 23814 11396 23818 11452
rect 23754 11392 23818 11396
rect 31219 11452 31283 11456
rect 31219 11396 31223 11452
rect 31223 11396 31279 11452
rect 31279 11396 31283 11452
rect 31219 11392 31283 11396
rect 31299 11452 31363 11456
rect 31299 11396 31303 11452
rect 31303 11396 31359 11452
rect 31359 11396 31363 11452
rect 31299 11392 31363 11396
rect 31379 11452 31443 11456
rect 31379 11396 31383 11452
rect 31383 11396 31439 11452
rect 31439 11396 31443 11452
rect 31379 11392 31443 11396
rect 31459 11452 31523 11456
rect 31459 11396 31463 11452
rect 31463 11396 31519 11452
rect 31519 11396 31523 11452
rect 31459 11392 31523 11396
rect 15148 11324 15212 11388
rect 4252 10908 4316 10912
rect 4252 10852 4256 10908
rect 4256 10852 4312 10908
rect 4312 10852 4316 10908
rect 4252 10848 4316 10852
rect 4332 10908 4396 10912
rect 4332 10852 4336 10908
rect 4336 10852 4392 10908
rect 4392 10852 4396 10908
rect 4332 10848 4396 10852
rect 4412 10908 4476 10912
rect 4412 10852 4416 10908
rect 4416 10852 4472 10908
rect 4472 10852 4476 10908
rect 4412 10848 4476 10852
rect 4492 10908 4556 10912
rect 4492 10852 4496 10908
rect 4496 10852 4552 10908
rect 4552 10852 4556 10908
rect 4492 10848 4556 10852
rect 11957 10908 12021 10912
rect 11957 10852 11961 10908
rect 11961 10852 12017 10908
rect 12017 10852 12021 10908
rect 11957 10848 12021 10852
rect 12037 10908 12101 10912
rect 12037 10852 12041 10908
rect 12041 10852 12097 10908
rect 12097 10852 12101 10908
rect 12037 10848 12101 10852
rect 12117 10908 12181 10912
rect 12117 10852 12121 10908
rect 12121 10852 12177 10908
rect 12177 10852 12181 10908
rect 12117 10848 12181 10852
rect 12197 10908 12261 10912
rect 12197 10852 12201 10908
rect 12201 10852 12257 10908
rect 12257 10852 12261 10908
rect 12197 10848 12261 10852
rect 16252 10916 16316 10980
rect 19662 10908 19726 10912
rect 19662 10852 19666 10908
rect 19666 10852 19722 10908
rect 19722 10852 19726 10908
rect 19662 10848 19726 10852
rect 19742 10908 19806 10912
rect 19742 10852 19746 10908
rect 19746 10852 19802 10908
rect 19802 10852 19806 10908
rect 19742 10848 19806 10852
rect 19822 10908 19886 10912
rect 19822 10852 19826 10908
rect 19826 10852 19882 10908
rect 19882 10852 19886 10908
rect 19822 10848 19886 10852
rect 19902 10908 19966 10912
rect 19902 10852 19906 10908
rect 19906 10852 19962 10908
rect 19962 10852 19966 10908
rect 19902 10848 19966 10852
rect 27367 10908 27431 10912
rect 27367 10852 27371 10908
rect 27371 10852 27427 10908
rect 27427 10852 27431 10908
rect 27367 10848 27431 10852
rect 27447 10908 27511 10912
rect 27447 10852 27451 10908
rect 27451 10852 27507 10908
rect 27507 10852 27511 10908
rect 27447 10848 27511 10852
rect 27527 10908 27591 10912
rect 27527 10852 27531 10908
rect 27531 10852 27587 10908
rect 27587 10852 27591 10908
rect 27527 10848 27591 10852
rect 27607 10908 27671 10912
rect 27607 10852 27611 10908
rect 27611 10852 27667 10908
rect 27667 10852 27671 10908
rect 27607 10848 27671 10852
rect 16436 10508 16500 10572
rect 19196 10508 19260 10572
rect 8104 10364 8168 10368
rect 8104 10308 8108 10364
rect 8108 10308 8164 10364
rect 8164 10308 8168 10364
rect 8104 10304 8168 10308
rect 8184 10364 8248 10368
rect 8184 10308 8188 10364
rect 8188 10308 8244 10364
rect 8244 10308 8248 10364
rect 8184 10304 8248 10308
rect 8264 10364 8328 10368
rect 8264 10308 8268 10364
rect 8268 10308 8324 10364
rect 8324 10308 8328 10364
rect 8264 10304 8328 10308
rect 8344 10364 8408 10368
rect 8344 10308 8348 10364
rect 8348 10308 8404 10364
rect 8404 10308 8408 10364
rect 8344 10304 8408 10308
rect 15809 10364 15873 10368
rect 15809 10308 15813 10364
rect 15813 10308 15869 10364
rect 15869 10308 15873 10364
rect 15809 10304 15873 10308
rect 15889 10364 15953 10368
rect 15889 10308 15893 10364
rect 15893 10308 15949 10364
rect 15949 10308 15953 10364
rect 15889 10304 15953 10308
rect 15969 10364 16033 10368
rect 15969 10308 15973 10364
rect 15973 10308 16029 10364
rect 16029 10308 16033 10364
rect 15969 10304 16033 10308
rect 16049 10364 16113 10368
rect 16049 10308 16053 10364
rect 16053 10308 16109 10364
rect 16109 10308 16113 10364
rect 16049 10304 16113 10308
rect 23514 10364 23578 10368
rect 23514 10308 23518 10364
rect 23518 10308 23574 10364
rect 23574 10308 23578 10364
rect 23514 10304 23578 10308
rect 23594 10364 23658 10368
rect 23594 10308 23598 10364
rect 23598 10308 23654 10364
rect 23654 10308 23658 10364
rect 23594 10304 23658 10308
rect 23674 10364 23738 10368
rect 23674 10308 23678 10364
rect 23678 10308 23734 10364
rect 23734 10308 23738 10364
rect 23674 10304 23738 10308
rect 23754 10364 23818 10368
rect 23754 10308 23758 10364
rect 23758 10308 23814 10364
rect 23814 10308 23818 10364
rect 23754 10304 23818 10308
rect 31219 10364 31283 10368
rect 31219 10308 31223 10364
rect 31223 10308 31279 10364
rect 31279 10308 31283 10364
rect 31219 10304 31283 10308
rect 31299 10364 31363 10368
rect 31299 10308 31303 10364
rect 31303 10308 31359 10364
rect 31359 10308 31363 10364
rect 31299 10304 31363 10308
rect 31379 10364 31443 10368
rect 31379 10308 31383 10364
rect 31383 10308 31439 10364
rect 31439 10308 31443 10364
rect 31379 10304 31443 10308
rect 31459 10364 31523 10368
rect 31459 10308 31463 10364
rect 31463 10308 31519 10364
rect 31519 10308 31523 10364
rect 31459 10304 31523 10308
rect 14780 10100 14844 10164
rect 17724 10160 17788 10164
rect 17724 10104 17774 10160
rect 17774 10104 17788 10160
rect 17724 10100 17788 10104
rect 19380 10100 19444 10164
rect 4252 9820 4316 9824
rect 4252 9764 4256 9820
rect 4256 9764 4312 9820
rect 4312 9764 4316 9820
rect 4252 9760 4316 9764
rect 4332 9820 4396 9824
rect 4332 9764 4336 9820
rect 4336 9764 4392 9820
rect 4392 9764 4396 9820
rect 4332 9760 4396 9764
rect 4412 9820 4476 9824
rect 4412 9764 4416 9820
rect 4416 9764 4472 9820
rect 4472 9764 4476 9820
rect 4412 9760 4476 9764
rect 4492 9820 4556 9824
rect 4492 9764 4496 9820
rect 4496 9764 4552 9820
rect 4552 9764 4556 9820
rect 4492 9760 4556 9764
rect 11957 9820 12021 9824
rect 11957 9764 11961 9820
rect 11961 9764 12017 9820
rect 12017 9764 12021 9820
rect 11957 9760 12021 9764
rect 12037 9820 12101 9824
rect 12037 9764 12041 9820
rect 12041 9764 12097 9820
rect 12097 9764 12101 9820
rect 12037 9760 12101 9764
rect 12117 9820 12181 9824
rect 12117 9764 12121 9820
rect 12121 9764 12177 9820
rect 12177 9764 12181 9820
rect 12117 9760 12181 9764
rect 12197 9820 12261 9824
rect 12197 9764 12201 9820
rect 12201 9764 12257 9820
rect 12257 9764 12261 9820
rect 12197 9760 12261 9764
rect 19662 9820 19726 9824
rect 19662 9764 19666 9820
rect 19666 9764 19722 9820
rect 19722 9764 19726 9820
rect 19662 9760 19726 9764
rect 19742 9820 19806 9824
rect 19742 9764 19746 9820
rect 19746 9764 19802 9820
rect 19802 9764 19806 9820
rect 19742 9760 19806 9764
rect 19822 9820 19886 9824
rect 19822 9764 19826 9820
rect 19826 9764 19882 9820
rect 19882 9764 19886 9820
rect 19822 9760 19886 9764
rect 19902 9820 19966 9824
rect 19902 9764 19906 9820
rect 19906 9764 19962 9820
rect 19962 9764 19966 9820
rect 19902 9760 19966 9764
rect 27367 9820 27431 9824
rect 27367 9764 27371 9820
rect 27371 9764 27427 9820
rect 27427 9764 27431 9820
rect 27367 9760 27431 9764
rect 27447 9820 27511 9824
rect 27447 9764 27451 9820
rect 27451 9764 27507 9820
rect 27507 9764 27511 9820
rect 27447 9760 27511 9764
rect 27527 9820 27591 9824
rect 27527 9764 27531 9820
rect 27531 9764 27587 9820
rect 27587 9764 27591 9820
rect 27527 9760 27591 9764
rect 27607 9820 27671 9824
rect 27607 9764 27611 9820
rect 27611 9764 27667 9820
rect 27667 9764 27671 9820
rect 27607 9760 27671 9764
rect 14964 9616 15028 9620
rect 14964 9560 14978 9616
rect 14978 9560 15028 9616
rect 14964 9556 15028 9560
rect 15516 9556 15580 9620
rect 16620 9616 16684 9620
rect 16620 9560 16670 9616
rect 16670 9560 16684 9616
rect 16620 9556 16684 9560
rect 17540 9616 17604 9620
rect 17540 9560 17590 9616
rect 17590 9560 17604 9616
rect 17540 9556 17604 9560
rect 18828 9556 18892 9620
rect 16988 9420 17052 9484
rect 17172 9420 17236 9484
rect 8104 9276 8168 9280
rect 8104 9220 8108 9276
rect 8108 9220 8164 9276
rect 8164 9220 8168 9276
rect 8104 9216 8168 9220
rect 8184 9276 8248 9280
rect 8184 9220 8188 9276
rect 8188 9220 8244 9276
rect 8244 9220 8248 9276
rect 8184 9216 8248 9220
rect 8264 9276 8328 9280
rect 8264 9220 8268 9276
rect 8268 9220 8324 9276
rect 8324 9220 8328 9276
rect 8264 9216 8328 9220
rect 8344 9276 8408 9280
rect 8344 9220 8348 9276
rect 8348 9220 8404 9276
rect 8404 9220 8408 9276
rect 8344 9216 8408 9220
rect 15809 9276 15873 9280
rect 15809 9220 15813 9276
rect 15813 9220 15869 9276
rect 15869 9220 15873 9276
rect 15809 9216 15873 9220
rect 15889 9276 15953 9280
rect 15889 9220 15893 9276
rect 15893 9220 15949 9276
rect 15949 9220 15953 9276
rect 15889 9216 15953 9220
rect 15969 9276 16033 9280
rect 15969 9220 15973 9276
rect 15973 9220 16029 9276
rect 16029 9220 16033 9276
rect 15969 9216 16033 9220
rect 16049 9276 16113 9280
rect 16049 9220 16053 9276
rect 16053 9220 16109 9276
rect 16109 9220 16113 9276
rect 16049 9216 16113 9220
rect 23514 9276 23578 9280
rect 23514 9220 23518 9276
rect 23518 9220 23574 9276
rect 23574 9220 23578 9276
rect 23514 9216 23578 9220
rect 23594 9276 23658 9280
rect 23594 9220 23598 9276
rect 23598 9220 23654 9276
rect 23654 9220 23658 9276
rect 23594 9216 23658 9220
rect 23674 9276 23738 9280
rect 23674 9220 23678 9276
rect 23678 9220 23734 9276
rect 23734 9220 23738 9276
rect 23674 9216 23738 9220
rect 23754 9276 23818 9280
rect 23754 9220 23758 9276
rect 23758 9220 23814 9276
rect 23814 9220 23818 9276
rect 23754 9216 23818 9220
rect 31219 9276 31283 9280
rect 31219 9220 31223 9276
rect 31223 9220 31279 9276
rect 31279 9220 31283 9276
rect 31219 9216 31283 9220
rect 31299 9276 31363 9280
rect 31299 9220 31303 9276
rect 31303 9220 31359 9276
rect 31359 9220 31363 9276
rect 31299 9216 31363 9220
rect 31379 9276 31443 9280
rect 31379 9220 31383 9276
rect 31383 9220 31439 9276
rect 31439 9220 31443 9276
rect 31379 9216 31443 9220
rect 31459 9276 31523 9280
rect 31459 9220 31463 9276
rect 31463 9220 31519 9276
rect 31519 9220 31523 9276
rect 31459 9216 31523 9220
rect 16988 9072 17052 9076
rect 16988 9016 17038 9072
rect 17038 9016 17052 9072
rect 16988 9012 17052 9016
rect 18460 9072 18524 9076
rect 18460 9016 18510 9072
rect 18510 9016 18524 9072
rect 18460 9012 18524 9016
rect 17540 8740 17604 8804
rect 17724 8800 17788 8804
rect 17724 8744 17738 8800
rect 17738 8744 17788 8800
rect 17724 8740 17788 8744
rect 4252 8732 4316 8736
rect 4252 8676 4256 8732
rect 4256 8676 4312 8732
rect 4312 8676 4316 8732
rect 4252 8672 4316 8676
rect 4332 8732 4396 8736
rect 4332 8676 4336 8732
rect 4336 8676 4392 8732
rect 4392 8676 4396 8732
rect 4332 8672 4396 8676
rect 4412 8732 4476 8736
rect 4412 8676 4416 8732
rect 4416 8676 4472 8732
rect 4472 8676 4476 8732
rect 4412 8672 4476 8676
rect 4492 8732 4556 8736
rect 4492 8676 4496 8732
rect 4496 8676 4552 8732
rect 4552 8676 4556 8732
rect 4492 8672 4556 8676
rect 11957 8732 12021 8736
rect 11957 8676 11961 8732
rect 11961 8676 12017 8732
rect 12017 8676 12021 8732
rect 11957 8672 12021 8676
rect 12037 8732 12101 8736
rect 12037 8676 12041 8732
rect 12041 8676 12097 8732
rect 12097 8676 12101 8732
rect 12037 8672 12101 8676
rect 12117 8732 12181 8736
rect 12117 8676 12121 8732
rect 12121 8676 12177 8732
rect 12177 8676 12181 8732
rect 12117 8672 12181 8676
rect 12197 8732 12261 8736
rect 12197 8676 12201 8732
rect 12201 8676 12257 8732
rect 12257 8676 12261 8732
rect 12197 8672 12261 8676
rect 19662 8732 19726 8736
rect 19662 8676 19666 8732
rect 19666 8676 19722 8732
rect 19722 8676 19726 8732
rect 19662 8672 19726 8676
rect 19742 8732 19806 8736
rect 19742 8676 19746 8732
rect 19746 8676 19802 8732
rect 19802 8676 19806 8732
rect 19742 8672 19806 8676
rect 19822 8732 19886 8736
rect 19822 8676 19826 8732
rect 19826 8676 19882 8732
rect 19882 8676 19886 8732
rect 19822 8672 19886 8676
rect 19902 8732 19966 8736
rect 19902 8676 19906 8732
rect 19906 8676 19962 8732
rect 19962 8676 19966 8732
rect 19902 8672 19966 8676
rect 27367 8732 27431 8736
rect 27367 8676 27371 8732
rect 27371 8676 27427 8732
rect 27427 8676 27431 8732
rect 27367 8672 27431 8676
rect 27447 8732 27511 8736
rect 27447 8676 27451 8732
rect 27451 8676 27507 8732
rect 27507 8676 27511 8732
rect 27447 8672 27511 8676
rect 27527 8732 27591 8736
rect 27527 8676 27531 8732
rect 27531 8676 27587 8732
rect 27587 8676 27591 8732
rect 27527 8672 27591 8676
rect 27607 8732 27671 8736
rect 27607 8676 27611 8732
rect 27611 8676 27667 8732
rect 27667 8676 27671 8732
rect 27607 8672 27671 8676
rect 14964 8604 15028 8668
rect 13676 8332 13740 8396
rect 17172 8332 17236 8396
rect 16436 8196 16500 8260
rect 8104 8188 8168 8192
rect 8104 8132 8108 8188
rect 8108 8132 8164 8188
rect 8164 8132 8168 8188
rect 8104 8128 8168 8132
rect 8184 8188 8248 8192
rect 8184 8132 8188 8188
rect 8188 8132 8244 8188
rect 8244 8132 8248 8188
rect 8184 8128 8248 8132
rect 8264 8188 8328 8192
rect 8264 8132 8268 8188
rect 8268 8132 8324 8188
rect 8324 8132 8328 8188
rect 8264 8128 8328 8132
rect 8344 8188 8408 8192
rect 8344 8132 8348 8188
rect 8348 8132 8404 8188
rect 8404 8132 8408 8188
rect 8344 8128 8408 8132
rect 15809 8188 15873 8192
rect 15809 8132 15813 8188
rect 15813 8132 15869 8188
rect 15869 8132 15873 8188
rect 15809 8128 15873 8132
rect 15889 8188 15953 8192
rect 15889 8132 15893 8188
rect 15893 8132 15949 8188
rect 15949 8132 15953 8188
rect 15889 8128 15953 8132
rect 15969 8188 16033 8192
rect 15969 8132 15973 8188
rect 15973 8132 16029 8188
rect 16029 8132 16033 8188
rect 15969 8128 16033 8132
rect 16049 8188 16113 8192
rect 16049 8132 16053 8188
rect 16053 8132 16109 8188
rect 16109 8132 16113 8188
rect 16049 8128 16113 8132
rect 23514 8188 23578 8192
rect 23514 8132 23518 8188
rect 23518 8132 23574 8188
rect 23574 8132 23578 8188
rect 23514 8128 23578 8132
rect 23594 8188 23658 8192
rect 23594 8132 23598 8188
rect 23598 8132 23654 8188
rect 23654 8132 23658 8188
rect 23594 8128 23658 8132
rect 23674 8188 23738 8192
rect 23674 8132 23678 8188
rect 23678 8132 23734 8188
rect 23734 8132 23738 8188
rect 23674 8128 23738 8132
rect 23754 8188 23818 8192
rect 23754 8132 23758 8188
rect 23758 8132 23814 8188
rect 23814 8132 23818 8188
rect 23754 8128 23818 8132
rect 31219 8188 31283 8192
rect 31219 8132 31223 8188
rect 31223 8132 31279 8188
rect 31279 8132 31283 8188
rect 31219 8128 31283 8132
rect 31299 8188 31363 8192
rect 31299 8132 31303 8188
rect 31303 8132 31359 8188
rect 31359 8132 31363 8188
rect 31299 8128 31363 8132
rect 31379 8188 31443 8192
rect 31379 8132 31383 8188
rect 31383 8132 31439 8188
rect 31439 8132 31443 8188
rect 31379 8128 31443 8132
rect 31459 8188 31523 8192
rect 31459 8132 31463 8188
rect 31463 8132 31519 8188
rect 31519 8132 31523 8188
rect 31459 8128 31523 8132
rect 19380 8060 19444 8124
rect 4252 7644 4316 7648
rect 4252 7588 4256 7644
rect 4256 7588 4312 7644
rect 4312 7588 4316 7644
rect 4252 7584 4316 7588
rect 4332 7644 4396 7648
rect 4332 7588 4336 7644
rect 4336 7588 4392 7644
rect 4392 7588 4396 7644
rect 4332 7584 4396 7588
rect 4412 7644 4476 7648
rect 4412 7588 4416 7644
rect 4416 7588 4472 7644
rect 4472 7588 4476 7644
rect 4412 7584 4476 7588
rect 4492 7644 4556 7648
rect 4492 7588 4496 7644
rect 4496 7588 4552 7644
rect 4552 7588 4556 7644
rect 4492 7584 4556 7588
rect 11957 7644 12021 7648
rect 11957 7588 11961 7644
rect 11961 7588 12017 7644
rect 12017 7588 12021 7644
rect 11957 7584 12021 7588
rect 12037 7644 12101 7648
rect 12037 7588 12041 7644
rect 12041 7588 12097 7644
rect 12097 7588 12101 7644
rect 12037 7584 12101 7588
rect 12117 7644 12181 7648
rect 12117 7588 12121 7644
rect 12121 7588 12177 7644
rect 12177 7588 12181 7644
rect 12117 7584 12181 7588
rect 12197 7644 12261 7648
rect 12197 7588 12201 7644
rect 12201 7588 12257 7644
rect 12257 7588 12261 7644
rect 12197 7584 12261 7588
rect 19662 7644 19726 7648
rect 19662 7588 19666 7644
rect 19666 7588 19722 7644
rect 19722 7588 19726 7644
rect 19662 7584 19726 7588
rect 19742 7644 19806 7648
rect 19742 7588 19746 7644
rect 19746 7588 19802 7644
rect 19802 7588 19806 7644
rect 19742 7584 19806 7588
rect 19822 7644 19886 7648
rect 19822 7588 19826 7644
rect 19826 7588 19882 7644
rect 19882 7588 19886 7644
rect 19822 7584 19886 7588
rect 19902 7644 19966 7648
rect 19902 7588 19906 7644
rect 19906 7588 19962 7644
rect 19962 7588 19966 7644
rect 19902 7584 19966 7588
rect 27367 7644 27431 7648
rect 27367 7588 27371 7644
rect 27371 7588 27427 7644
rect 27427 7588 27431 7644
rect 27367 7584 27431 7588
rect 27447 7644 27511 7648
rect 27447 7588 27451 7644
rect 27451 7588 27507 7644
rect 27507 7588 27511 7644
rect 27447 7584 27511 7588
rect 27527 7644 27591 7648
rect 27527 7588 27531 7644
rect 27531 7588 27587 7644
rect 27587 7588 27591 7644
rect 27527 7584 27591 7588
rect 27607 7644 27671 7648
rect 27607 7588 27611 7644
rect 27611 7588 27667 7644
rect 27667 7588 27671 7644
rect 27607 7584 27671 7588
rect 8104 7100 8168 7104
rect 8104 7044 8108 7100
rect 8108 7044 8164 7100
rect 8164 7044 8168 7100
rect 8104 7040 8168 7044
rect 8184 7100 8248 7104
rect 8184 7044 8188 7100
rect 8188 7044 8244 7100
rect 8244 7044 8248 7100
rect 8184 7040 8248 7044
rect 8264 7100 8328 7104
rect 8264 7044 8268 7100
rect 8268 7044 8324 7100
rect 8324 7044 8328 7100
rect 8264 7040 8328 7044
rect 8344 7100 8408 7104
rect 8344 7044 8348 7100
rect 8348 7044 8404 7100
rect 8404 7044 8408 7100
rect 8344 7040 8408 7044
rect 15809 7100 15873 7104
rect 15809 7044 15813 7100
rect 15813 7044 15869 7100
rect 15869 7044 15873 7100
rect 15809 7040 15873 7044
rect 15889 7100 15953 7104
rect 15889 7044 15893 7100
rect 15893 7044 15949 7100
rect 15949 7044 15953 7100
rect 15889 7040 15953 7044
rect 15969 7100 16033 7104
rect 15969 7044 15973 7100
rect 15973 7044 16029 7100
rect 16029 7044 16033 7100
rect 15969 7040 16033 7044
rect 16049 7100 16113 7104
rect 16049 7044 16053 7100
rect 16053 7044 16109 7100
rect 16109 7044 16113 7100
rect 16049 7040 16113 7044
rect 23514 7100 23578 7104
rect 23514 7044 23518 7100
rect 23518 7044 23574 7100
rect 23574 7044 23578 7100
rect 23514 7040 23578 7044
rect 23594 7100 23658 7104
rect 23594 7044 23598 7100
rect 23598 7044 23654 7100
rect 23654 7044 23658 7100
rect 23594 7040 23658 7044
rect 23674 7100 23738 7104
rect 23674 7044 23678 7100
rect 23678 7044 23734 7100
rect 23734 7044 23738 7100
rect 23674 7040 23738 7044
rect 23754 7100 23818 7104
rect 23754 7044 23758 7100
rect 23758 7044 23814 7100
rect 23814 7044 23818 7100
rect 23754 7040 23818 7044
rect 31219 7100 31283 7104
rect 31219 7044 31223 7100
rect 31223 7044 31279 7100
rect 31279 7044 31283 7100
rect 31219 7040 31283 7044
rect 31299 7100 31363 7104
rect 31299 7044 31303 7100
rect 31303 7044 31359 7100
rect 31359 7044 31363 7100
rect 31299 7040 31363 7044
rect 31379 7100 31443 7104
rect 31379 7044 31383 7100
rect 31383 7044 31439 7100
rect 31439 7044 31443 7100
rect 31379 7040 31443 7044
rect 31459 7100 31523 7104
rect 31459 7044 31463 7100
rect 31463 7044 31519 7100
rect 31519 7044 31523 7100
rect 31459 7040 31523 7044
rect 14044 6836 14108 6900
rect 14228 6700 14292 6764
rect 4252 6556 4316 6560
rect 4252 6500 4256 6556
rect 4256 6500 4312 6556
rect 4312 6500 4316 6556
rect 4252 6496 4316 6500
rect 4332 6556 4396 6560
rect 4332 6500 4336 6556
rect 4336 6500 4392 6556
rect 4392 6500 4396 6556
rect 4332 6496 4396 6500
rect 4412 6556 4476 6560
rect 4412 6500 4416 6556
rect 4416 6500 4472 6556
rect 4472 6500 4476 6556
rect 4412 6496 4476 6500
rect 4492 6556 4556 6560
rect 4492 6500 4496 6556
rect 4496 6500 4552 6556
rect 4552 6500 4556 6556
rect 4492 6496 4556 6500
rect 11957 6556 12021 6560
rect 11957 6500 11961 6556
rect 11961 6500 12017 6556
rect 12017 6500 12021 6556
rect 11957 6496 12021 6500
rect 12037 6556 12101 6560
rect 12037 6500 12041 6556
rect 12041 6500 12097 6556
rect 12097 6500 12101 6556
rect 12037 6496 12101 6500
rect 12117 6556 12181 6560
rect 12117 6500 12121 6556
rect 12121 6500 12177 6556
rect 12177 6500 12181 6556
rect 12117 6496 12181 6500
rect 12197 6556 12261 6560
rect 12197 6500 12201 6556
rect 12201 6500 12257 6556
rect 12257 6500 12261 6556
rect 12197 6496 12261 6500
rect 19662 6556 19726 6560
rect 19662 6500 19666 6556
rect 19666 6500 19722 6556
rect 19722 6500 19726 6556
rect 19662 6496 19726 6500
rect 19742 6556 19806 6560
rect 19742 6500 19746 6556
rect 19746 6500 19802 6556
rect 19802 6500 19806 6556
rect 19742 6496 19806 6500
rect 19822 6556 19886 6560
rect 19822 6500 19826 6556
rect 19826 6500 19882 6556
rect 19882 6500 19886 6556
rect 19822 6496 19886 6500
rect 19902 6556 19966 6560
rect 19902 6500 19906 6556
rect 19906 6500 19962 6556
rect 19962 6500 19966 6556
rect 19902 6496 19966 6500
rect 27367 6556 27431 6560
rect 27367 6500 27371 6556
rect 27371 6500 27427 6556
rect 27427 6500 27431 6556
rect 27367 6496 27431 6500
rect 27447 6556 27511 6560
rect 27447 6500 27451 6556
rect 27451 6500 27507 6556
rect 27507 6500 27511 6556
rect 27447 6496 27511 6500
rect 27527 6556 27591 6560
rect 27527 6500 27531 6556
rect 27531 6500 27587 6556
rect 27587 6500 27591 6556
rect 27527 6496 27591 6500
rect 27607 6556 27671 6560
rect 27607 6500 27611 6556
rect 27611 6500 27667 6556
rect 27667 6500 27671 6556
rect 27607 6496 27671 6500
rect 15148 6292 15212 6356
rect 14780 6156 14844 6220
rect 18460 6156 18524 6220
rect 8104 6012 8168 6016
rect 8104 5956 8108 6012
rect 8108 5956 8164 6012
rect 8164 5956 8168 6012
rect 8104 5952 8168 5956
rect 8184 6012 8248 6016
rect 8184 5956 8188 6012
rect 8188 5956 8244 6012
rect 8244 5956 8248 6012
rect 8184 5952 8248 5956
rect 8264 6012 8328 6016
rect 8264 5956 8268 6012
rect 8268 5956 8324 6012
rect 8324 5956 8328 6012
rect 8264 5952 8328 5956
rect 8344 6012 8408 6016
rect 8344 5956 8348 6012
rect 8348 5956 8404 6012
rect 8404 5956 8408 6012
rect 8344 5952 8408 5956
rect 15809 6012 15873 6016
rect 15809 5956 15813 6012
rect 15813 5956 15869 6012
rect 15869 5956 15873 6012
rect 15809 5952 15873 5956
rect 15889 6012 15953 6016
rect 15889 5956 15893 6012
rect 15893 5956 15949 6012
rect 15949 5956 15953 6012
rect 15889 5952 15953 5956
rect 15969 6012 16033 6016
rect 15969 5956 15973 6012
rect 15973 5956 16029 6012
rect 16029 5956 16033 6012
rect 15969 5952 16033 5956
rect 16049 6012 16113 6016
rect 16049 5956 16053 6012
rect 16053 5956 16109 6012
rect 16109 5956 16113 6012
rect 16049 5952 16113 5956
rect 23514 6012 23578 6016
rect 23514 5956 23518 6012
rect 23518 5956 23574 6012
rect 23574 5956 23578 6012
rect 23514 5952 23578 5956
rect 23594 6012 23658 6016
rect 23594 5956 23598 6012
rect 23598 5956 23654 6012
rect 23654 5956 23658 6012
rect 23594 5952 23658 5956
rect 23674 6012 23738 6016
rect 23674 5956 23678 6012
rect 23678 5956 23734 6012
rect 23734 5956 23738 6012
rect 23674 5952 23738 5956
rect 23754 6012 23818 6016
rect 23754 5956 23758 6012
rect 23758 5956 23814 6012
rect 23814 5956 23818 6012
rect 23754 5952 23818 5956
rect 31219 6012 31283 6016
rect 31219 5956 31223 6012
rect 31223 5956 31279 6012
rect 31279 5956 31283 6012
rect 31219 5952 31283 5956
rect 31299 6012 31363 6016
rect 31299 5956 31303 6012
rect 31303 5956 31359 6012
rect 31359 5956 31363 6012
rect 31299 5952 31363 5956
rect 31379 6012 31443 6016
rect 31379 5956 31383 6012
rect 31383 5956 31439 6012
rect 31439 5956 31443 6012
rect 31379 5952 31443 5956
rect 31459 6012 31523 6016
rect 31459 5956 31463 6012
rect 31463 5956 31519 6012
rect 31519 5956 31523 6012
rect 31459 5952 31523 5956
rect 4252 5468 4316 5472
rect 4252 5412 4256 5468
rect 4256 5412 4312 5468
rect 4312 5412 4316 5468
rect 4252 5408 4316 5412
rect 4332 5468 4396 5472
rect 4332 5412 4336 5468
rect 4336 5412 4392 5468
rect 4392 5412 4396 5468
rect 4332 5408 4396 5412
rect 4412 5468 4476 5472
rect 4412 5412 4416 5468
rect 4416 5412 4472 5468
rect 4472 5412 4476 5468
rect 4412 5408 4476 5412
rect 4492 5468 4556 5472
rect 4492 5412 4496 5468
rect 4496 5412 4552 5468
rect 4552 5412 4556 5468
rect 4492 5408 4556 5412
rect 11957 5468 12021 5472
rect 11957 5412 11961 5468
rect 11961 5412 12017 5468
rect 12017 5412 12021 5468
rect 11957 5408 12021 5412
rect 12037 5468 12101 5472
rect 12037 5412 12041 5468
rect 12041 5412 12097 5468
rect 12097 5412 12101 5468
rect 12037 5408 12101 5412
rect 12117 5468 12181 5472
rect 12117 5412 12121 5468
rect 12121 5412 12177 5468
rect 12177 5412 12181 5468
rect 12117 5408 12181 5412
rect 12197 5468 12261 5472
rect 12197 5412 12201 5468
rect 12201 5412 12257 5468
rect 12257 5412 12261 5468
rect 12197 5408 12261 5412
rect 19662 5468 19726 5472
rect 19662 5412 19666 5468
rect 19666 5412 19722 5468
rect 19722 5412 19726 5468
rect 19662 5408 19726 5412
rect 19742 5468 19806 5472
rect 19742 5412 19746 5468
rect 19746 5412 19802 5468
rect 19802 5412 19806 5468
rect 19742 5408 19806 5412
rect 19822 5468 19886 5472
rect 19822 5412 19826 5468
rect 19826 5412 19882 5468
rect 19882 5412 19886 5468
rect 19822 5408 19886 5412
rect 19902 5468 19966 5472
rect 19902 5412 19906 5468
rect 19906 5412 19962 5468
rect 19962 5412 19966 5468
rect 19902 5408 19966 5412
rect 27367 5468 27431 5472
rect 27367 5412 27371 5468
rect 27371 5412 27427 5468
rect 27427 5412 27431 5468
rect 27367 5408 27431 5412
rect 27447 5468 27511 5472
rect 27447 5412 27451 5468
rect 27451 5412 27507 5468
rect 27507 5412 27511 5468
rect 27447 5408 27511 5412
rect 27527 5468 27591 5472
rect 27527 5412 27531 5468
rect 27531 5412 27587 5468
rect 27587 5412 27591 5468
rect 27527 5408 27591 5412
rect 27607 5468 27671 5472
rect 27607 5412 27611 5468
rect 27611 5412 27667 5468
rect 27667 5412 27671 5468
rect 27607 5408 27671 5412
rect 16252 5340 16316 5404
rect 8104 4924 8168 4928
rect 8104 4868 8108 4924
rect 8108 4868 8164 4924
rect 8164 4868 8168 4924
rect 8104 4864 8168 4868
rect 8184 4924 8248 4928
rect 8184 4868 8188 4924
rect 8188 4868 8244 4924
rect 8244 4868 8248 4924
rect 8184 4864 8248 4868
rect 8264 4924 8328 4928
rect 8264 4868 8268 4924
rect 8268 4868 8324 4924
rect 8324 4868 8328 4924
rect 8264 4864 8328 4868
rect 8344 4924 8408 4928
rect 8344 4868 8348 4924
rect 8348 4868 8404 4924
rect 8404 4868 8408 4924
rect 8344 4864 8408 4868
rect 15809 4924 15873 4928
rect 15809 4868 15813 4924
rect 15813 4868 15869 4924
rect 15869 4868 15873 4924
rect 15809 4864 15873 4868
rect 15889 4924 15953 4928
rect 15889 4868 15893 4924
rect 15893 4868 15949 4924
rect 15949 4868 15953 4924
rect 15889 4864 15953 4868
rect 15969 4924 16033 4928
rect 15969 4868 15973 4924
rect 15973 4868 16029 4924
rect 16029 4868 16033 4924
rect 15969 4864 16033 4868
rect 16049 4924 16113 4928
rect 16049 4868 16053 4924
rect 16053 4868 16109 4924
rect 16109 4868 16113 4924
rect 16049 4864 16113 4868
rect 23514 4924 23578 4928
rect 23514 4868 23518 4924
rect 23518 4868 23574 4924
rect 23574 4868 23578 4924
rect 23514 4864 23578 4868
rect 23594 4924 23658 4928
rect 23594 4868 23598 4924
rect 23598 4868 23654 4924
rect 23654 4868 23658 4924
rect 23594 4864 23658 4868
rect 23674 4924 23738 4928
rect 23674 4868 23678 4924
rect 23678 4868 23734 4924
rect 23734 4868 23738 4924
rect 23674 4864 23738 4868
rect 23754 4924 23818 4928
rect 23754 4868 23758 4924
rect 23758 4868 23814 4924
rect 23814 4868 23818 4924
rect 23754 4864 23818 4868
rect 31219 4924 31283 4928
rect 31219 4868 31223 4924
rect 31223 4868 31279 4924
rect 31279 4868 31283 4924
rect 31219 4864 31283 4868
rect 31299 4924 31363 4928
rect 31299 4868 31303 4924
rect 31303 4868 31359 4924
rect 31359 4868 31363 4924
rect 31299 4864 31363 4868
rect 31379 4924 31443 4928
rect 31379 4868 31383 4924
rect 31383 4868 31439 4924
rect 31439 4868 31443 4924
rect 31379 4864 31443 4868
rect 31459 4924 31523 4928
rect 31459 4868 31463 4924
rect 31463 4868 31519 4924
rect 31519 4868 31523 4924
rect 31459 4864 31523 4868
rect 15516 4388 15580 4452
rect 17908 4388 17972 4452
rect 4252 4380 4316 4384
rect 4252 4324 4256 4380
rect 4256 4324 4312 4380
rect 4312 4324 4316 4380
rect 4252 4320 4316 4324
rect 4332 4380 4396 4384
rect 4332 4324 4336 4380
rect 4336 4324 4392 4380
rect 4392 4324 4396 4380
rect 4332 4320 4396 4324
rect 4412 4380 4476 4384
rect 4412 4324 4416 4380
rect 4416 4324 4472 4380
rect 4472 4324 4476 4380
rect 4412 4320 4476 4324
rect 4492 4380 4556 4384
rect 4492 4324 4496 4380
rect 4496 4324 4552 4380
rect 4552 4324 4556 4380
rect 4492 4320 4556 4324
rect 11957 4380 12021 4384
rect 11957 4324 11961 4380
rect 11961 4324 12017 4380
rect 12017 4324 12021 4380
rect 11957 4320 12021 4324
rect 12037 4380 12101 4384
rect 12037 4324 12041 4380
rect 12041 4324 12097 4380
rect 12097 4324 12101 4380
rect 12037 4320 12101 4324
rect 12117 4380 12181 4384
rect 12117 4324 12121 4380
rect 12121 4324 12177 4380
rect 12177 4324 12181 4380
rect 12117 4320 12181 4324
rect 12197 4380 12261 4384
rect 12197 4324 12201 4380
rect 12201 4324 12257 4380
rect 12257 4324 12261 4380
rect 12197 4320 12261 4324
rect 19662 4380 19726 4384
rect 19662 4324 19666 4380
rect 19666 4324 19722 4380
rect 19722 4324 19726 4380
rect 19662 4320 19726 4324
rect 19742 4380 19806 4384
rect 19742 4324 19746 4380
rect 19746 4324 19802 4380
rect 19802 4324 19806 4380
rect 19742 4320 19806 4324
rect 19822 4380 19886 4384
rect 19822 4324 19826 4380
rect 19826 4324 19882 4380
rect 19882 4324 19886 4380
rect 19822 4320 19886 4324
rect 19902 4380 19966 4384
rect 19902 4324 19906 4380
rect 19906 4324 19962 4380
rect 19962 4324 19966 4380
rect 19902 4320 19966 4324
rect 27367 4380 27431 4384
rect 27367 4324 27371 4380
rect 27371 4324 27427 4380
rect 27427 4324 27431 4380
rect 27367 4320 27431 4324
rect 27447 4380 27511 4384
rect 27447 4324 27451 4380
rect 27451 4324 27507 4380
rect 27507 4324 27511 4380
rect 27447 4320 27511 4324
rect 27527 4380 27591 4384
rect 27527 4324 27531 4380
rect 27531 4324 27587 4380
rect 27587 4324 27591 4380
rect 27527 4320 27591 4324
rect 27607 4380 27671 4384
rect 27607 4324 27611 4380
rect 27611 4324 27667 4380
rect 27667 4324 27671 4380
rect 27607 4320 27671 4324
rect 13676 3980 13740 4044
rect 8104 3836 8168 3840
rect 8104 3780 8108 3836
rect 8108 3780 8164 3836
rect 8164 3780 8168 3836
rect 8104 3776 8168 3780
rect 8184 3836 8248 3840
rect 8184 3780 8188 3836
rect 8188 3780 8244 3836
rect 8244 3780 8248 3836
rect 8184 3776 8248 3780
rect 8264 3836 8328 3840
rect 8264 3780 8268 3836
rect 8268 3780 8324 3836
rect 8324 3780 8328 3836
rect 8264 3776 8328 3780
rect 8344 3836 8408 3840
rect 8344 3780 8348 3836
rect 8348 3780 8404 3836
rect 8404 3780 8408 3836
rect 8344 3776 8408 3780
rect 15809 3836 15873 3840
rect 15809 3780 15813 3836
rect 15813 3780 15869 3836
rect 15869 3780 15873 3836
rect 15809 3776 15873 3780
rect 15889 3836 15953 3840
rect 15889 3780 15893 3836
rect 15893 3780 15949 3836
rect 15949 3780 15953 3836
rect 15889 3776 15953 3780
rect 15969 3836 16033 3840
rect 15969 3780 15973 3836
rect 15973 3780 16029 3836
rect 16029 3780 16033 3836
rect 15969 3776 16033 3780
rect 16049 3836 16113 3840
rect 16049 3780 16053 3836
rect 16053 3780 16109 3836
rect 16109 3780 16113 3836
rect 16049 3776 16113 3780
rect 23514 3836 23578 3840
rect 23514 3780 23518 3836
rect 23518 3780 23574 3836
rect 23574 3780 23578 3836
rect 23514 3776 23578 3780
rect 23594 3836 23658 3840
rect 23594 3780 23598 3836
rect 23598 3780 23654 3836
rect 23654 3780 23658 3836
rect 23594 3776 23658 3780
rect 23674 3836 23738 3840
rect 23674 3780 23678 3836
rect 23678 3780 23734 3836
rect 23734 3780 23738 3836
rect 23674 3776 23738 3780
rect 23754 3836 23818 3840
rect 23754 3780 23758 3836
rect 23758 3780 23814 3836
rect 23814 3780 23818 3836
rect 23754 3776 23818 3780
rect 31219 3836 31283 3840
rect 31219 3780 31223 3836
rect 31223 3780 31279 3836
rect 31279 3780 31283 3836
rect 31219 3776 31283 3780
rect 31299 3836 31363 3840
rect 31299 3780 31303 3836
rect 31303 3780 31359 3836
rect 31359 3780 31363 3836
rect 31299 3776 31363 3780
rect 31379 3836 31443 3840
rect 31379 3780 31383 3836
rect 31383 3780 31439 3836
rect 31439 3780 31443 3836
rect 31379 3776 31443 3780
rect 31459 3836 31523 3840
rect 31459 3780 31463 3836
rect 31463 3780 31519 3836
rect 31519 3780 31523 3836
rect 31459 3776 31523 3780
rect 4252 3292 4316 3296
rect 4252 3236 4256 3292
rect 4256 3236 4312 3292
rect 4312 3236 4316 3292
rect 4252 3232 4316 3236
rect 4332 3292 4396 3296
rect 4332 3236 4336 3292
rect 4336 3236 4392 3292
rect 4392 3236 4396 3292
rect 4332 3232 4396 3236
rect 4412 3292 4476 3296
rect 4412 3236 4416 3292
rect 4416 3236 4472 3292
rect 4472 3236 4476 3292
rect 4412 3232 4476 3236
rect 4492 3292 4556 3296
rect 4492 3236 4496 3292
rect 4496 3236 4552 3292
rect 4552 3236 4556 3292
rect 4492 3232 4556 3236
rect 11957 3292 12021 3296
rect 11957 3236 11961 3292
rect 11961 3236 12017 3292
rect 12017 3236 12021 3292
rect 11957 3232 12021 3236
rect 12037 3292 12101 3296
rect 12037 3236 12041 3292
rect 12041 3236 12097 3292
rect 12097 3236 12101 3292
rect 12037 3232 12101 3236
rect 12117 3292 12181 3296
rect 12117 3236 12121 3292
rect 12121 3236 12177 3292
rect 12177 3236 12181 3292
rect 12117 3232 12181 3236
rect 12197 3292 12261 3296
rect 12197 3236 12201 3292
rect 12201 3236 12257 3292
rect 12257 3236 12261 3292
rect 12197 3232 12261 3236
rect 19662 3292 19726 3296
rect 19662 3236 19666 3292
rect 19666 3236 19722 3292
rect 19722 3236 19726 3292
rect 19662 3232 19726 3236
rect 19742 3292 19806 3296
rect 19742 3236 19746 3292
rect 19746 3236 19802 3292
rect 19802 3236 19806 3292
rect 19742 3232 19806 3236
rect 19822 3292 19886 3296
rect 19822 3236 19826 3292
rect 19826 3236 19882 3292
rect 19882 3236 19886 3292
rect 19822 3232 19886 3236
rect 19902 3292 19966 3296
rect 19902 3236 19906 3292
rect 19906 3236 19962 3292
rect 19962 3236 19966 3292
rect 19902 3232 19966 3236
rect 27367 3292 27431 3296
rect 27367 3236 27371 3292
rect 27371 3236 27427 3292
rect 27427 3236 27431 3292
rect 27367 3232 27431 3236
rect 27447 3292 27511 3296
rect 27447 3236 27451 3292
rect 27451 3236 27507 3292
rect 27507 3236 27511 3292
rect 27447 3232 27511 3236
rect 27527 3292 27591 3296
rect 27527 3236 27531 3292
rect 27531 3236 27587 3292
rect 27587 3236 27591 3292
rect 27527 3232 27591 3236
rect 27607 3292 27671 3296
rect 27607 3236 27611 3292
rect 27611 3236 27667 3292
rect 27667 3236 27671 3292
rect 27607 3232 27671 3236
rect 14964 2892 15028 2956
rect 8104 2748 8168 2752
rect 8104 2692 8108 2748
rect 8108 2692 8164 2748
rect 8164 2692 8168 2748
rect 8104 2688 8168 2692
rect 8184 2748 8248 2752
rect 8184 2692 8188 2748
rect 8188 2692 8244 2748
rect 8244 2692 8248 2748
rect 8184 2688 8248 2692
rect 8264 2748 8328 2752
rect 8264 2692 8268 2748
rect 8268 2692 8324 2748
rect 8324 2692 8328 2748
rect 8264 2688 8328 2692
rect 8344 2748 8408 2752
rect 8344 2692 8348 2748
rect 8348 2692 8404 2748
rect 8404 2692 8408 2748
rect 8344 2688 8408 2692
rect 15809 2748 15873 2752
rect 15809 2692 15813 2748
rect 15813 2692 15869 2748
rect 15869 2692 15873 2748
rect 15809 2688 15873 2692
rect 15889 2748 15953 2752
rect 15889 2692 15893 2748
rect 15893 2692 15949 2748
rect 15949 2692 15953 2748
rect 15889 2688 15953 2692
rect 15969 2748 16033 2752
rect 15969 2692 15973 2748
rect 15973 2692 16029 2748
rect 16029 2692 16033 2748
rect 15969 2688 16033 2692
rect 16049 2748 16113 2752
rect 16049 2692 16053 2748
rect 16053 2692 16109 2748
rect 16109 2692 16113 2748
rect 16049 2688 16113 2692
rect 23514 2748 23578 2752
rect 23514 2692 23518 2748
rect 23518 2692 23574 2748
rect 23574 2692 23578 2748
rect 23514 2688 23578 2692
rect 23594 2748 23658 2752
rect 23594 2692 23598 2748
rect 23598 2692 23654 2748
rect 23654 2692 23658 2748
rect 23594 2688 23658 2692
rect 23674 2748 23738 2752
rect 23674 2692 23678 2748
rect 23678 2692 23734 2748
rect 23734 2692 23738 2748
rect 23674 2688 23738 2692
rect 23754 2748 23818 2752
rect 23754 2692 23758 2748
rect 23758 2692 23814 2748
rect 23814 2692 23818 2748
rect 23754 2688 23818 2692
rect 31219 2748 31283 2752
rect 31219 2692 31223 2748
rect 31223 2692 31279 2748
rect 31279 2692 31283 2748
rect 31219 2688 31283 2692
rect 31299 2748 31363 2752
rect 31299 2692 31303 2748
rect 31303 2692 31359 2748
rect 31359 2692 31363 2748
rect 31299 2688 31363 2692
rect 31379 2748 31443 2752
rect 31379 2692 31383 2748
rect 31383 2692 31439 2748
rect 31439 2692 31443 2748
rect 31379 2688 31443 2692
rect 31459 2748 31523 2752
rect 31459 2692 31463 2748
rect 31463 2692 31519 2748
rect 31519 2692 31523 2748
rect 31459 2688 31523 2692
rect 4252 2204 4316 2208
rect 4252 2148 4256 2204
rect 4256 2148 4312 2204
rect 4312 2148 4316 2204
rect 4252 2144 4316 2148
rect 4332 2204 4396 2208
rect 4332 2148 4336 2204
rect 4336 2148 4392 2204
rect 4392 2148 4396 2204
rect 4332 2144 4396 2148
rect 4412 2204 4476 2208
rect 4412 2148 4416 2204
rect 4416 2148 4472 2204
rect 4472 2148 4476 2204
rect 4412 2144 4476 2148
rect 4492 2204 4556 2208
rect 4492 2148 4496 2204
rect 4496 2148 4552 2204
rect 4552 2148 4556 2204
rect 4492 2144 4556 2148
rect 11957 2204 12021 2208
rect 11957 2148 11961 2204
rect 11961 2148 12017 2204
rect 12017 2148 12021 2204
rect 11957 2144 12021 2148
rect 12037 2204 12101 2208
rect 12037 2148 12041 2204
rect 12041 2148 12097 2204
rect 12097 2148 12101 2204
rect 12037 2144 12101 2148
rect 12117 2204 12181 2208
rect 12117 2148 12121 2204
rect 12121 2148 12177 2204
rect 12177 2148 12181 2204
rect 12117 2144 12181 2148
rect 12197 2204 12261 2208
rect 12197 2148 12201 2204
rect 12201 2148 12257 2204
rect 12257 2148 12261 2204
rect 12197 2144 12261 2148
rect 19662 2204 19726 2208
rect 19662 2148 19666 2204
rect 19666 2148 19722 2204
rect 19722 2148 19726 2204
rect 19662 2144 19726 2148
rect 19742 2204 19806 2208
rect 19742 2148 19746 2204
rect 19746 2148 19802 2204
rect 19802 2148 19806 2204
rect 19742 2144 19806 2148
rect 19822 2204 19886 2208
rect 19822 2148 19826 2204
rect 19826 2148 19882 2204
rect 19882 2148 19886 2204
rect 19822 2144 19886 2148
rect 19902 2204 19966 2208
rect 19902 2148 19906 2204
rect 19906 2148 19962 2204
rect 19962 2148 19966 2204
rect 19902 2144 19966 2148
rect 27367 2204 27431 2208
rect 27367 2148 27371 2204
rect 27371 2148 27427 2204
rect 27427 2148 27431 2204
rect 27367 2144 27431 2148
rect 27447 2204 27511 2208
rect 27447 2148 27451 2204
rect 27451 2148 27507 2204
rect 27507 2148 27511 2204
rect 27447 2144 27511 2148
rect 27527 2204 27591 2208
rect 27527 2148 27531 2204
rect 27531 2148 27587 2204
rect 27587 2148 27591 2204
rect 27527 2144 27591 2148
rect 27607 2204 27671 2208
rect 27607 2148 27611 2204
rect 27611 2148 27667 2204
rect 27667 2148 27671 2204
rect 27607 2144 27671 2148
rect 8104 1660 8168 1664
rect 8104 1604 8108 1660
rect 8108 1604 8164 1660
rect 8164 1604 8168 1660
rect 8104 1600 8168 1604
rect 8184 1660 8248 1664
rect 8184 1604 8188 1660
rect 8188 1604 8244 1660
rect 8244 1604 8248 1660
rect 8184 1600 8248 1604
rect 8264 1660 8328 1664
rect 8264 1604 8268 1660
rect 8268 1604 8324 1660
rect 8324 1604 8328 1660
rect 8264 1600 8328 1604
rect 8344 1660 8408 1664
rect 8344 1604 8348 1660
rect 8348 1604 8404 1660
rect 8404 1604 8408 1660
rect 8344 1600 8408 1604
rect 15809 1660 15873 1664
rect 15809 1604 15813 1660
rect 15813 1604 15869 1660
rect 15869 1604 15873 1660
rect 15809 1600 15873 1604
rect 15889 1660 15953 1664
rect 15889 1604 15893 1660
rect 15893 1604 15949 1660
rect 15949 1604 15953 1660
rect 15889 1600 15953 1604
rect 15969 1660 16033 1664
rect 15969 1604 15973 1660
rect 15973 1604 16029 1660
rect 16029 1604 16033 1660
rect 15969 1600 16033 1604
rect 16049 1660 16113 1664
rect 16049 1604 16053 1660
rect 16053 1604 16109 1660
rect 16109 1604 16113 1660
rect 16049 1600 16113 1604
rect 23514 1660 23578 1664
rect 23514 1604 23518 1660
rect 23518 1604 23574 1660
rect 23574 1604 23578 1660
rect 23514 1600 23578 1604
rect 23594 1660 23658 1664
rect 23594 1604 23598 1660
rect 23598 1604 23654 1660
rect 23654 1604 23658 1660
rect 23594 1600 23658 1604
rect 23674 1660 23738 1664
rect 23674 1604 23678 1660
rect 23678 1604 23734 1660
rect 23734 1604 23738 1660
rect 23674 1600 23738 1604
rect 23754 1660 23818 1664
rect 23754 1604 23758 1660
rect 23758 1604 23814 1660
rect 23814 1604 23818 1660
rect 23754 1600 23818 1604
rect 31219 1660 31283 1664
rect 31219 1604 31223 1660
rect 31223 1604 31279 1660
rect 31279 1604 31283 1660
rect 31219 1600 31283 1604
rect 31299 1660 31363 1664
rect 31299 1604 31303 1660
rect 31303 1604 31359 1660
rect 31359 1604 31363 1660
rect 31299 1600 31363 1604
rect 31379 1660 31443 1664
rect 31379 1604 31383 1660
rect 31383 1604 31439 1660
rect 31439 1604 31443 1660
rect 31379 1600 31443 1604
rect 31459 1660 31523 1664
rect 31459 1604 31463 1660
rect 31463 1604 31519 1660
rect 31519 1604 31523 1660
rect 31459 1600 31523 1604
rect 4252 1116 4316 1120
rect 4252 1060 4256 1116
rect 4256 1060 4312 1116
rect 4312 1060 4316 1116
rect 4252 1056 4316 1060
rect 4332 1116 4396 1120
rect 4332 1060 4336 1116
rect 4336 1060 4392 1116
rect 4392 1060 4396 1116
rect 4332 1056 4396 1060
rect 4412 1116 4476 1120
rect 4412 1060 4416 1116
rect 4416 1060 4472 1116
rect 4472 1060 4476 1116
rect 4412 1056 4476 1060
rect 4492 1116 4556 1120
rect 4492 1060 4496 1116
rect 4496 1060 4552 1116
rect 4552 1060 4556 1116
rect 4492 1056 4556 1060
rect 11957 1116 12021 1120
rect 11957 1060 11961 1116
rect 11961 1060 12017 1116
rect 12017 1060 12021 1116
rect 11957 1056 12021 1060
rect 12037 1116 12101 1120
rect 12037 1060 12041 1116
rect 12041 1060 12097 1116
rect 12097 1060 12101 1116
rect 12037 1056 12101 1060
rect 12117 1116 12181 1120
rect 12117 1060 12121 1116
rect 12121 1060 12177 1116
rect 12177 1060 12181 1116
rect 12117 1056 12181 1060
rect 12197 1116 12261 1120
rect 12197 1060 12201 1116
rect 12201 1060 12257 1116
rect 12257 1060 12261 1116
rect 12197 1056 12261 1060
rect 19662 1116 19726 1120
rect 19662 1060 19666 1116
rect 19666 1060 19722 1116
rect 19722 1060 19726 1116
rect 19662 1056 19726 1060
rect 19742 1116 19806 1120
rect 19742 1060 19746 1116
rect 19746 1060 19802 1116
rect 19802 1060 19806 1116
rect 19742 1056 19806 1060
rect 19822 1116 19886 1120
rect 19822 1060 19826 1116
rect 19826 1060 19882 1116
rect 19882 1060 19886 1116
rect 19822 1056 19886 1060
rect 19902 1116 19966 1120
rect 19902 1060 19906 1116
rect 19906 1060 19962 1116
rect 19962 1060 19966 1116
rect 19902 1056 19966 1060
rect 27367 1116 27431 1120
rect 27367 1060 27371 1116
rect 27371 1060 27427 1116
rect 27427 1060 27431 1116
rect 27367 1056 27431 1060
rect 27447 1116 27511 1120
rect 27447 1060 27451 1116
rect 27451 1060 27507 1116
rect 27507 1060 27511 1116
rect 27447 1056 27511 1060
rect 27527 1116 27591 1120
rect 27527 1060 27531 1116
rect 27531 1060 27587 1116
rect 27587 1060 27591 1116
rect 27527 1056 27591 1060
rect 27607 1116 27671 1120
rect 27607 1060 27611 1116
rect 27611 1060 27667 1116
rect 27667 1060 27671 1116
rect 27607 1056 27671 1060
rect 8104 572 8168 576
rect 8104 516 8108 572
rect 8108 516 8164 572
rect 8164 516 8168 572
rect 8104 512 8168 516
rect 8184 572 8248 576
rect 8184 516 8188 572
rect 8188 516 8244 572
rect 8244 516 8248 572
rect 8184 512 8248 516
rect 8264 572 8328 576
rect 8264 516 8268 572
rect 8268 516 8324 572
rect 8324 516 8328 572
rect 8264 512 8328 516
rect 8344 572 8408 576
rect 8344 516 8348 572
rect 8348 516 8404 572
rect 8404 516 8408 572
rect 8344 512 8408 516
rect 15809 572 15873 576
rect 15809 516 15813 572
rect 15813 516 15869 572
rect 15869 516 15873 572
rect 15809 512 15873 516
rect 15889 572 15953 576
rect 15889 516 15893 572
rect 15893 516 15949 572
rect 15949 516 15953 572
rect 15889 512 15953 516
rect 15969 572 16033 576
rect 15969 516 15973 572
rect 15973 516 16029 572
rect 16029 516 16033 572
rect 15969 512 16033 516
rect 16049 572 16113 576
rect 16049 516 16053 572
rect 16053 516 16109 572
rect 16109 516 16113 572
rect 16049 512 16113 516
rect 23514 572 23578 576
rect 23514 516 23518 572
rect 23518 516 23574 572
rect 23574 516 23578 572
rect 23514 512 23578 516
rect 23594 572 23658 576
rect 23594 516 23598 572
rect 23598 516 23654 572
rect 23654 516 23658 572
rect 23594 512 23658 516
rect 23674 572 23738 576
rect 23674 516 23678 572
rect 23678 516 23734 572
rect 23734 516 23738 572
rect 23674 512 23738 516
rect 23754 572 23818 576
rect 23754 516 23758 572
rect 23758 516 23814 572
rect 23814 516 23818 572
rect 23754 512 23818 516
rect 31219 572 31283 576
rect 31219 516 31223 572
rect 31223 516 31279 572
rect 31279 516 31283 572
rect 31219 512 31283 516
rect 31299 572 31363 576
rect 31299 516 31303 572
rect 31303 516 31359 572
rect 31359 516 31363 572
rect 31299 512 31363 516
rect 31379 572 31443 576
rect 31379 516 31383 572
rect 31383 516 31439 572
rect 31439 516 31443 572
rect 31379 512 31443 516
rect 31459 572 31523 576
rect 31459 516 31463 572
rect 31463 516 31519 572
rect 31519 516 31523 572
rect 31459 512 31523 516
<< metal4 >>
rect 4244 18528 4564 19088
rect 4244 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4564 18528
rect 4244 17440 4564 18464
rect 4244 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4564 17440
rect 4244 16352 4564 17376
rect 4244 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4564 16352
rect 4244 15264 4564 16288
rect 4244 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4564 15264
rect 4244 14176 4564 15200
rect 4244 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4564 14176
rect 4244 13088 4564 14112
rect 4244 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4564 13088
rect 4244 12000 4564 13024
rect 4244 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4564 12000
rect 4244 10912 4564 11936
rect 4244 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4564 10912
rect 4244 9824 4564 10848
rect 4244 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4564 9824
rect 4244 8736 4564 9760
rect 4244 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4564 8736
rect 4244 7648 4564 8672
rect 4244 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4564 7648
rect 4244 6560 4564 7584
rect 4244 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4564 6560
rect 4244 5472 4564 6496
rect 4244 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4564 5472
rect 4244 4384 4564 5408
rect 4244 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4564 4384
rect 4244 3296 4564 4320
rect 4244 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4564 3296
rect 4244 2208 4564 3232
rect 4244 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4564 2208
rect 4244 1120 4564 2144
rect 4244 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4564 1120
rect 4244 496 4564 1056
rect 8096 19072 8416 19088
rect 8096 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8416 19072
rect 8096 17984 8416 19008
rect 8096 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8416 17984
rect 8096 16896 8416 17920
rect 8096 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8416 16896
rect 8096 15808 8416 16832
rect 8096 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8416 15808
rect 8096 14720 8416 15744
rect 8096 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8416 14720
rect 8096 13632 8416 14656
rect 8096 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8416 13632
rect 8096 12544 8416 13568
rect 8096 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8416 12544
rect 8096 11456 8416 12480
rect 8096 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8416 11456
rect 8096 10368 8416 11392
rect 8096 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8416 10368
rect 8096 9280 8416 10304
rect 8096 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8416 9280
rect 8096 8192 8416 9216
rect 8096 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8416 8192
rect 8096 7104 8416 8128
rect 8096 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8416 7104
rect 8096 6016 8416 7040
rect 8096 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8416 6016
rect 8096 4928 8416 5952
rect 8096 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8416 4928
rect 8096 3840 8416 4864
rect 8096 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8416 3840
rect 8096 2752 8416 3776
rect 8096 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8416 2752
rect 8096 1664 8416 2688
rect 8096 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8416 1664
rect 8096 576 8416 1600
rect 8096 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8416 576
rect 8096 496 8416 512
rect 11949 18528 12269 19088
rect 11949 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12269 18528
rect 11949 17440 12269 18464
rect 15801 19072 16121 19088
rect 15801 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16121 19072
rect 14963 18052 15029 18053
rect 14963 17988 14964 18052
rect 15028 17988 15029 18052
rect 14963 17987 15029 17988
rect 11949 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12269 17440
rect 11949 16352 12269 17376
rect 11949 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12269 16352
rect 11949 15264 12269 16288
rect 11949 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12269 15264
rect 11949 14176 12269 15200
rect 11949 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12269 14176
rect 11949 13088 12269 14112
rect 11949 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12269 13088
rect 11949 12000 12269 13024
rect 14411 12884 14477 12885
rect 14411 12820 14412 12884
rect 14476 12820 14477 12884
rect 14411 12819 14477 12820
rect 14043 12612 14109 12613
rect 14043 12548 14044 12612
rect 14108 12548 14109 12612
rect 14043 12547 14109 12548
rect 11949 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12269 12000
rect 11949 10912 12269 11936
rect 11949 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12269 10912
rect 11949 9824 12269 10848
rect 11949 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12269 9824
rect 11949 8736 12269 9760
rect 11949 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12269 8736
rect 11949 7648 12269 8672
rect 13675 8396 13741 8397
rect 13675 8332 13676 8396
rect 13740 8332 13741 8396
rect 13675 8331 13741 8332
rect 11949 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12269 7648
rect 11949 6560 12269 7584
rect 11949 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12269 6560
rect 11949 5472 12269 6496
rect 11949 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12269 5472
rect 11949 4384 12269 5408
rect 11949 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12269 4384
rect 11949 3296 12269 4320
rect 13678 4045 13738 8331
rect 14046 6901 14106 12547
rect 14414 12450 14474 12819
rect 14230 12390 14474 12450
rect 14043 6900 14109 6901
rect 14043 6836 14044 6900
rect 14108 6836 14109 6900
rect 14043 6835 14109 6836
rect 14230 6765 14290 12390
rect 14779 10164 14845 10165
rect 14779 10100 14780 10164
rect 14844 10100 14845 10164
rect 14779 10099 14845 10100
rect 14227 6764 14293 6765
rect 14227 6700 14228 6764
rect 14292 6700 14293 6764
rect 14227 6699 14293 6700
rect 14782 6221 14842 10099
rect 14966 9621 15026 17987
rect 15801 17984 16121 19008
rect 15801 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16121 17984
rect 15801 16896 16121 17920
rect 15801 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16121 16896
rect 15801 15808 16121 16832
rect 19654 18528 19974 19088
rect 19654 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19974 18528
rect 19654 17440 19974 18464
rect 19654 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19974 17440
rect 18827 16692 18893 16693
rect 18827 16628 18828 16692
rect 18892 16628 18893 16692
rect 18827 16627 18893 16628
rect 16619 16012 16685 16013
rect 16619 15948 16620 16012
rect 16684 15948 16685 16012
rect 16619 15947 16685 15948
rect 15801 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16121 15808
rect 15801 14720 16121 15744
rect 15801 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16121 14720
rect 15801 13632 16121 14656
rect 15801 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16121 13632
rect 15801 12544 16121 13568
rect 15801 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16121 12544
rect 15801 11456 16121 12480
rect 15801 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16121 11456
rect 15147 11388 15213 11389
rect 15147 11324 15148 11388
rect 15212 11324 15213 11388
rect 15147 11323 15213 11324
rect 14963 9620 15029 9621
rect 14963 9556 14964 9620
rect 15028 9556 15029 9620
rect 14963 9555 15029 9556
rect 14963 8668 15029 8669
rect 14963 8604 14964 8668
rect 15028 8604 15029 8668
rect 14963 8603 15029 8604
rect 14779 6220 14845 6221
rect 14779 6156 14780 6220
rect 14844 6156 14845 6220
rect 14779 6155 14845 6156
rect 13675 4044 13741 4045
rect 13675 3980 13676 4044
rect 13740 3980 13741 4044
rect 13675 3979 13741 3980
rect 11949 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12269 3296
rect 11949 2208 12269 3232
rect 14966 2957 15026 8603
rect 15150 6357 15210 11323
rect 15801 10368 16121 11392
rect 16251 10980 16317 10981
rect 16251 10916 16252 10980
rect 16316 10916 16317 10980
rect 16251 10915 16317 10916
rect 15801 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16121 10368
rect 15515 9620 15581 9621
rect 15515 9556 15516 9620
rect 15580 9556 15581 9620
rect 15515 9555 15581 9556
rect 15147 6356 15213 6357
rect 15147 6292 15148 6356
rect 15212 6292 15213 6356
rect 15147 6291 15213 6292
rect 15518 4453 15578 9555
rect 15801 9280 16121 10304
rect 15801 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16121 9280
rect 15801 8192 16121 9216
rect 15801 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16121 8192
rect 15801 7104 16121 8128
rect 15801 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16121 7104
rect 15801 6016 16121 7040
rect 15801 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16121 6016
rect 15801 4928 16121 5952
rect 16254 5405 16314 10915
rect 16435 10572 16501 10573
rect 16435 10508 16436 10572
rect 16500 10508 16501 10572
rect 16435 10507 16501 10508
rect 16438 8261 16498 10507
rect 16622 9621 16682 15947
rect 16987 14652 17053 14653
rect 16987 14588 16988 14652
rect 17052 14588 17053 14652
rect 16987 14587 17053 14588
rect 16803 13836 16869 13837
rect 16803 13772 16804 13836
rect 16868 13772 16869 13836
rect 16803 13771 16869 13772
rect 16806 11525 16866 13771
rect 16803 11524 16869 11525
rect 16803 11460 16804 11524
rect 16868 11460 16869 11524
rect 16803 11459 16869 11460
rect 16619 9620 16685 9621
rect 16619 9556 16620 9620
rect 16684 9556 16685 9620
rect 16619 9555 16685 9556
rect 16990 9485 17050 14587
rect 17907 11796 17973 11797
rect 17907 11732 17908 11796
rect 17972 11732 17973 11796
rect 17907 11731 17973 11732
rect 17723 10164 17789 10165
rect 17723 10100 17724 10164
rect 17788 10100 17789 10164
rect 17723 10099 17789 10100
rect 17539 9620 17605 9621
rect 17539 9556 17540 9620
rect 17604 9556 17605 9620
rect 17539 9555 17605 9556
rect 16987 9484 17053 9485
rect 16987 9420 16988 9484
rect 17052 9420 17053 9484
rect 16987 9419 17053 9420
rect 17171 9484 17237 9485
rect 17171 9420 17172 9484
rect 17236 9420 17237 9484
rect 17171 9419 17237 9420
rect 16990 9077 17050 9419
rect 16987 9076 17053 9077
rect 16987 9012 16988 9076
rect 17052 9012 17053 9076
rect 16987 9011 17053 9012
rect 17174 8397 17234 9419
rect 17542 8805 17602 9555
rect 17726 8805 17786 10099
rect 17539 8804 17605 8805
rect 17539 8740 17540 8804
rect 17604 8740 17605 8804
rect 17539 8739 17605 8740
rect 17723 8804 17789 8805
rect 17723 8740 17724 8804
rect 17788 8740 17789 8804
rect 17723 8739 17789 8740
rect 17171 8396 17237 8397
rect 17171 8332 17172 8396
rect 17236 8332 17237 8396
rect 17171 8331 17237 8332
rect 16435 8260 16501 8261
rect 16435 8196 16436 8260
rect 16500 8196 16501 8260
rect 16435 8195 16501 8196
rect 16251 5404 16317 5405
rect 16251 5340 16252 5404
rect 16316 5340 16317 5404
rect 16251 5339 16317 5340
rect 15801 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16121 4928
rect 15515 4452 15581 4453
rect 15515 4388 15516 4452
rect 15580 4388 15581 4452
rect 15515 4387 15581 4388
rect 15801 3840 16121 4864
rect 17910 4453 17970 11731
rect 18830 9621 18890 16627
rect 19654 16352 19974 17376
rect 19654 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19974 16352
rect 19654 15264 19974 16288
rect 19654 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19974 15264
rect 19654 14176 19974 15200
rect 19654 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19974 14176
rect 19654 13088 19974 14112
rect 19654 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19974 13088
rect 19195 13020 19261 13021
rect 19195 12956 19196 13020
rect 19260 12956 19261 13020
rect 19195 12955 19261 12956
rect 19198 10573 19258 12955
rect 19654 12000 19974 13024
rect 19654 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19974 12000
rect 19654 10912 19974 11936
rect 19654 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19974 10912
rect 19195 10572 19261 10573
rect 19195 10508 19196 10572
rect 19260 10508 19261 10572
rect 19195 10507 19261 10508
rect 19379 10164 19445 10165
rect 19379 10100 19380 10164
rect 19444 10100 19445 10164
rect 19379 10099 19445 10100
rect 18827 9620 18893 9621
rect 18827 9556 18828 9620
rect 18892 9556 18893 9620
rect 18827 9555 18893 9556
rect 18459 9076 18525 9077
rect 18459 9012 18460 9076
rect 18524 9012 18525 9076
rect 18459 9011 18525 9012
rect 18462 6221 18522 9011
rect 19382 8125 19442 10099
rect 19654 9824 19974 10848
rect 19654 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19974 9824
rect 19654 8736 19974 9760
rect 19654 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19974 8736
rect 19379 8124 19445 8125
rect 19379 8060 19380 8124
rect 19444 8060 19445 8124
rect 19379 8059 19445 8060
rect 19654 7648 19974 8672
rect 19654 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19974 7648
rect 19654 6560 19974 7584
rect 19654 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19974 6560
rect 18459 6220 18525 6221
rect 18459 6156 18460 6220
rect 18524 6156 18525 6220
rect 18459 6155 18525 6156
rect 19654 5472 19974 6496
rect 19654 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19974 5472
rect 17907 4452 17973 4453
rect 17907 4388 17908 4452
rect 17972 4388 17973 4452
rect 17907 4387 17973 4388
rect 15801 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16121 3840
rect 14963 2956 15029 2957
rect 14963 2892 14964 2956
rect 15028 2892 15029 2956
rect 14963 2891 15029 2892
rect 11949 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12269 2208
rect 11949 1120 12269 2144
rect 11949 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12269 1120
rect 11949 496 12269 1056
rect 15801 2752 16121 3776
rect 15801 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16121 2752
rect 15801 1664 16121 2688
rect 15801 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16121 1664
rect 15801 576 16121 1600
rect 15801 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16121 576
rect 15801 496 16121 512
rect 19654 4384 19974 5408
rect 19654 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19974 4384
rect 19654 3296 19974 4320
rect 19654 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19974 3296
rect 19654 2208 19974 3232
rect 19654 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19974 2208
rect 19654 1120 19974 2144
rect 19654 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19974 1120
rect 19654 496 19974 1056
rect 23506 19072 23826 19088
rect 23506 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23826 19072
rect 23506 17984 23826 19008
rect 23506 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23826 17984
rect 23506 16896 23826 17920
rect 23506 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23826 16896
rect 23506 15808 23826 16832
rect 23506 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23826 15808
rect 23506 14720 23826 15744
rect 23506 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23826 14720
rect 23506 13632 23826 14656
rect 23506 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23826 13632
rect 23506 12544 23826 13568
rect 23506 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23826 12544
rect 23506 11456 23826 12480
rect 23506 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23826 11456
rect 23506 10368 23826 11392
rect 23506 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23826 10368
rect 23506 9280 23826 10304
rect 23506 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23826 9280
rect 23506 8192 23826 9216
rect 23506 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23826 8192
rect 23506 7104 23826 8128
rect 23506 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23826 7104
rect 23506 6016 23826 7040
rect 23506 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23826 6016
rect 23506 4928 23826 5952
rect 23506 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23826 4928
rect 23506 3840 23826 4864
rect 23506 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23826 3840
rect 23506 2752 23826 3776
rect 23506 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23826 2752
rect 23506 1664 23826 2688
rect 23506 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23826 1664
rect 23506 576 23826 1600
rect 23506 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23826 576
rect 23506 496 23826 512
rect 27359 18528 27679 19088
rect 27359 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27679 18528
rect 27359 17440 27679 18464
rect 27359 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27679 17440
rect 27359 16352 27679 17376
rect 27359 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27679 16352
rect 27359 15264 27679 16288
rect 27359 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27679 15264
rect 27359 14176 27679 15200
rect 27359 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27679 14176
rect 27359 13088 27679 14112
rect 27359 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27679 13088
rect 27359 12000 27679 13024
rect 27359 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27679 12000
rect 27359 10912 27679 11936
rect 27359 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27679 10912
rect 27359 9824 27679 10848
rect 27359 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27679 9824
rect 27359 8736 27679 9760
rect 27359 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27679 8736
rect 27359 7648 27679 8672
rect 27359 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27679 7648
rect 27359 6560 27679 7584
rect 27359 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27679 6560
rect 27359 5472 27679 6496
rect 27359 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27679 5472
rect 27359 4384 27679 5408
rect 27359 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27679 4384
rect 27359 3296 27679 4320
rect 27359 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27679 3296
rect 27359 2208 27679 3232
rect 27359 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27679 2208
rect 27359 1120 27679 2144
rect 27359 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27679 1120
rect 27359 496 27679 1056
rect 31211 19072 31531 19088
rect 31211 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31531 19072
rect 31211 17984 31531 19008
rect 31211 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31531 17984
rect 31211 16896 31531 17920
rect 31211 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31531 16896
rect 31211 15808 31531 16832
rect 31211 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31531 15808
rect 31211 14720 31531 15744
rect 31211 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31531 14720
rect 31211 13632 31531 14656
rect 31211 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31531 13632
rect 31211 12544 31531 13568
rect 31211 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31531 12544
rect 31211 11456 31531 12480
rect 31211 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31531 11456
rect 31211 10368 31531 11392
rect 31211 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31531 10368
rect 31211 9280 31531 10304
rect 31211 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31531 9280
rect 31211 8192 31531 9216
rect 31211 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31531 8192
rect 31211 7104 31531 8128
rect 31211 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31531 7104
rect 31211 6016 31531 7040
rect 31211 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31531 6016
rect 31211 4928 31531 5952
rect 31211 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31531 4928
rect 31211 3840 31531 4864
rect 31211 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31531 3840
rect 31211 2752 31531 3776
rect 31211 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31531 2752
rect 31211 1664 31531 2688
rect 31211 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31531 1664
rect 31211 576 31531 1600
rect 31211 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31531 576
rect 31211 496 31531 512
use sky130_fd_sc_hd__nor3_1  _211_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17480 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _212_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18032 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _213_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16652 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _214_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18676 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _215_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 21252 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _216_
timestamp 1701704242
transform 1 0 14996 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _217_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15640 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _218_
timestamp 1701704242
transform -1 0 15272 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _219_
timestamp 1701704242
transform 1 0 15548 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _220_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _221_
timestamp 1701704242
transform 1 0 17664 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_4  _222_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16468 0 -1 5984
box -38 -48 1418 592
use sky130_fd_sc_hd__buf_2  _223_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 19780 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _224_
timestamp 1701704242
transform -1 0 16008 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _225_
timestamp 1701704242
transform -1 0 16284 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _226_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 23920 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _227_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 19688 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _228_
timestamp 1701704242
transform 1 0 19228 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _229_
timestamp 1701704242
transform 1 0 17296 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _230_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18492 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _231_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17940 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _232_
timestamp 1701704242
transform -1 0 17112 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _233_
timestamp 1701704242
transform -1 0 16836 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _234_
timestamp 1701704242
transform -1 0 14444 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _235_
timestamp 1701704242
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _236_
timestamp 1701704242
transform 1 0 13984 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _237_
timestamp 1701704242
transform -1 0 15640 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _238_
timestamp 1701704242
transform -1 0 12052 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _239_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8372 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _240_
timestamp 1701704242
transform 1 0 17572 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _241_
timestamp 1701704242
transform 1 0 17296 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _242_
timestamp 1701704242
transform 1 0 18676 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _243_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15456 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _244_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 17664 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _245_
timestamp 1701704242
transform -1 0 17756 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _246_
timestamp 1701704242
transform -1 0 14720 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _247_
timestamp 1701704242
transform 1 0 16652 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _248_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16652 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _249_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17296 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _250_
timestamp 1701704242
transform 1 0 15272 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _251_
timestamp 1701704242
transform -1 0 17756 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _252_
timestamp 1701704242
transform 1 0 13708 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _253_
timestamp 1701704242
transform 1 0 16192 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _254_
timestamp 1701704242
transform 1 0 17204 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _255_
timestamp 1701704242
transform 1 0 13432 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _256_
timestamp 1701704242
transform -1 0 19780 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _257_
timestamp 1701704242
transform -1 0 14352 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _258_
timestamp 1701704242
transform -1 0 15548 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _259_
timestamp 1701704242
transform 1 0 16192 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _260_
timestamp 1701704242
transform -1 0 17572 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _261_
timestamp 1701704242
transform -1 0 17204 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _262_
timestamp 1701704242
transform 1 0 20332 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _263_
timestamp 1701704242
transform -1 0 23460 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _264_
timestamp 1701704242
transform -1 0 17480 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _265_
timestamp 1701704242
transform 1 0 17112 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _266_
timestamp 1701704242
transform 1 0 20884 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _267_
timestamp 1701704242
transform -1 0 16836 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _268_
timestamp 1701704242
transform 1 0 16284 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _269_
timestamp 1701704242
transform 1 0 18676 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _270_
timestamp 1701704242
transform 1 0 16468 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _271_
timestamp 1701704242
transform 1 0 16100 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _272_
timestamp 1701704242
transform -1 0 19320 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _273_
timestamp 1701704242
transform 1 0 16560 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _274_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16560 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_4  _275_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 19228 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__o32a_4  _276_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 20332 0 1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__and2_2  _277_
timestamp 1701704242
transform 1 0 16652 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _278_
timestamp 1701704242
transform 1 0 18676 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _279_
timestamp 1701704242
transform -1 0 24840 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _280_
timestamp 1701704242
transform -1 0 21896 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _281_
timestamp 1701704242
transform 1 0 19872 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _282_
timestamp 1701704242
transform -1 0 20608 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _283_
timestamp 1701704242
transform 1 0 20516 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _284_
timestamp 1701704242
transform 1 0 13984 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _285_
timestamp 1701704242
transform -1 0 15088 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _286_
timestamp 1701704242
transform -1 0 14536 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _287_
timestamp 1701704242
transform -1 0 14812 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _288_
timestamp 1701704242
transform -1 0 14352 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _289_
timestamp 1701704242
transform 1 0 14352 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _290_
timestamp 1701704242
transform -1 0 19504 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _291_
timestamp 1701704242
transform 1 0 14168 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _292_
timestamp 1701704242
transform 1 0 14720 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _293_
timestamp 1701704242
transform 1 0 14996 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _294_
timestamp 1701704242
transform -1 0 21712 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _295_
timestamp 1701704242
transform 1 0 14352 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _296_
timestamp 1701704242
transform 1 0 14812 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _297_
timestamp 1701704242
transform -1 0 16652 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _298_
timestamp 1701704242
transform 1 0 11776 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _299_
timestamp 1701704242
transform 1 0 11132 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _300_
timestamp 1701704242
transform 1 0 11224 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _301_
timestamp 1701704242
transform -1 0 13156 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _302_
timestamp 1701704242
transform 1 0 14536 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_4  _303_
timestamp 1701704242
transform 1 0 24104 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__a32o_1  _304_
timestamp 1701704242
transform 1 0 14628 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _305_
timestamp 1701704242
transform 1 0 7452 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _306_
timestamp 1701704242
transform 1 0 13524 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _307_
timestamp 1701704242
transform 1 0 16652 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _308_
timestamp 1701704242
transform -1 0 18768 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _309_
timestamp 1701704242
transform -1 0 19044 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _310_
timestamp 1701704242
transform 1 0 17480 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _311_
timestamp 1701704242
transform 1 0 14076 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _312_
timestamp 1701704242
transform 1 0 14352 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _313_
timestamp 1701704242
transform 1 0 14536 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _314_
timestamp 1701704242
transform 1 0 14904 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _315_
timestamp 1701704242
transform 1 0 15364 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _316_
timestamp 1701704242
transform -1 0 22172 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _317_
timestamp 1701704242
transform 1 0 17020 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _318_
timestamp 1701704242
transform -1 0 17848 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _319_
timestamp 1701704242
transform -1 0 25760 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _320_
timestamp 1701704242
transform 1 0 21896 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _321_
timestamp 1701704242
transform -1 0 24748 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _322_
timestamp 1701704242
transform 1 0 23828 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _323_
timestamp 1701704242
transform 1 0 17204 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_4  _324_
timestamp 1701704242
transform 1 0 17388 0 -1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__a32o_1  _325_
timestamp 1701704242
transform -1 0 18124 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _326_
timestamp 1701704242
transform -1 0 18216 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _327_
timestamp 1701704242
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _328_
timestamp 1701704242
transform 1 0 15916 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _329_
timestamp 1701704242
transform -1 0 20240 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _330_
timestamp 1701704242
transform 1 0 12512 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _331_
timestamp 1701704242
transform 1 0 14352 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _332_
timestamp 1701704242
transform -1 0 20424 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _333_
timestamp 1701704242
transform 1 0 13708 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _334_
timestamp 1701704242
transform 1 0 14076 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _335_
timestamp 1701704242
transform -1 0 14904 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _336_
timestamp 1701704242
transform 1 0 12512 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _337_
timestamp 1701704242
transform -1 0 15548 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _338_
timestamp 1701704242
transform 1 0 11408 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _339_
timestamp 1701704242
transform -1 0 13248 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _340_
timestamp 1701704242
transform 1 0 23276 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _341_
timestamp 1701704242
transform -1 0 25116 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _342_
timestamp 1701704242
transform -1 0 24288 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _343_
timestamp 1701704242
transform 1 0 23184 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _344_
timestamp 1701704242
transform 1 0 15088 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_4  _345_
timestamp 1701704242
transform 1 0 17940 0 -1 10336
box -38 -48 1694 592
use sky130_fd_sc_hd__a22o_1  _346_
timestamp 1701704242
transform -1 0 5704 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _347_
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _348_
timestamp 1701704242
transform 1 0 22540 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _349_
timestamp 1701704242
transform 1 0 15916 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _350_
timestamp 1701704242
transform 1 0 12972 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _351_
timestamp 1701704242
transform -1 0 20424 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _352_
timestamp 1701704242
transform 1 0 19412 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _353_
timestamp 1701704242
transform 1 0 11684 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _354_
timestamp 1701704242
transform 1 0 12696 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _355_
timestamp 1701704242
transform -1 0 19228 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _356_
timestamp 1701704242
transform -1 0 13984 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _357_
timestamp 1701704242
transform -1 0 19136 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _358_
timestamp 1701704242
transform 1 0 12144 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _359_
timestamp 1701704242
transform 1 0 17848 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _360_
timestamp 1701704242
transform -1 0 18676 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _361_
timestamp 1701704242
transform -1 0 23736 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _362_
timestamp 1701704242
transform -1 0 23276 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _363_
timestamp 1701704242
transform 1 0 22264 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _364_
timestamp 1701704242
transform 1 0 22724 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _365_
timestamp 1701704242
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_4  _366_
timestamp 1701704242
transform 1 0 18676 0 1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__a22o_1  _367_
timestamp 1701704242
transform 1 0 17664 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _368_
timestamp 1701704242
transform 1 0 23920 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _369_
timestamp 1701704242
transform -1 0 13708 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _370_
timestamp 1701704242
transform 1 0 22724 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _371_
timestamp 1701704242
transform 1 0 13248 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _372_
timestamp 1701704242
transform 1 0 12972 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _373_
timestamp 1701704242
transform -1 0 14352 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _374_
timestamp 1701704242
transform -1 0 19780 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _375_
timestamp 1701704242
transform -1 0 20240 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _376_
timestamp 1701704242
transform -1 0 20700 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _377_
timestamp 1701704242
transform -1 0 19780 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _378_
timestamp 1701704242
transform -1 0 15272 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _379_
timestamp 1701704242
transform -1 0 23000 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _380_
timestamp 1701704242
transform 1 0 12696 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _381_
timestamp 1701704242
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _382_
timestamp 1701704242
transform 1 0 12512 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _383_
timestamp 1701704242
transform 1 0 11684 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _384_
timestamp 1701704242
transform -1 0 17020 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _385_
timestamp 1701704242
transform -1 0 13064 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _386_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12972 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_4  _387_
timestamp 1701704242
transform 1 0 23920 0 -1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__a22o_1  _388_
timestamp 1701704242
transform 1 0 4968 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _389_
timestamp 1701704242
transform 1 0 5612 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _390_
timestamp 1701704242
transform -1 0 15548 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _391_
timestamp 1701704242
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _392_
timestamp 1701704242
transform 1 0 18124 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _393_
timestamp 1701704242
transform -1 0 20332 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _394_
timestamp 1701704242
transform 1 0 19688 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _395_
timestamp 1701704242
transform 1 0 12880 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _396_
timestamp 1701704242
transform 1 0 12788 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _397_
timestamp 1701704242
transform 1 0 13340 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _398_
timestamp 1701704242
transform -1 0 14352 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _399_
timestamp 1701704242
transform 1 0 14260 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _400_
timestamp 1701704242
transform -1 0 21988 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _401_
timestamp 1701704242
transform 1 0 19872 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _402_
timestamp 1701704242
transform 1 0 20332 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _403_
timestamp 1701704242
transform -1 0 25300 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _404_
timestamp 1701704242
transform 1 0 23828 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _405_
timestamp 1701704242
transform 1 0 23276 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _406_
timestamp 1701704242
transform 1 0 23920 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _407_
timestamp 1701704242
transform 1 0 19136 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_4  _408_
timestamp 1701704242
transform 1 0 19228 0 -1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__a22o_1  _409_
timestamp 1701704242
transform 1 0 8464 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _410_
timestamp 1701704242
transform 1 0 6164 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _411_
timestamp 1701704242
transform -1 0 23736 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _412_
timestamp 1701704242
transform 1 0 23828 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _413_
timestamp 1701704242
transform 1 0 14904 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _414_
timestamp 1701704242
transform -1 0 20884 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _415_
timestamp 1701704242
transform 1 0 20240 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _416_
timestamp 1701704242
transform 1 0 12972 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _417_
timestamp 1701704242
transform 1 0 12972 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _418_
timestamp 1701704242
transform 1 0 13616 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _419_
timestamp 1701704242
transform -1 0 14352 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _420_
timestamp 1701704242
transform -1 0 19964 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _421_
timestamp 1701704242
transform 1 0 11500 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _422_
timestamp 1701704242
transform -1 0 19780 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _423_
timestamp 1701704242
transform -1 0 19688 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _424_
timestamp 1701704242
transform 1 0 15548 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _425_
timestamp 1701704242
transform -1 0 20884 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _426_
timestamp 1701704242
transform 1 0 18676 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _427_
timestamp 1701704242
transform 1 0 19136 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _428_
timestamp 1701704242
transform 1 0 19228 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_4  _429_
timestamp 1701704242
transform 1 0 20148 0 1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__dfxtp_1  _430_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 26128 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _431_
timestamp 1701704242
transform -1 0 27232 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _432_
timestamp 1701704242
transform -1 0 24472 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _433_
timestamp 1701704242
transform -1 0 28336 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _434_
timestamp 1701704242
transform -1 0 27600 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _435_
timestamp 1701704242
transform -1 0 28336 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _436_
timestamp 1701704242
transform -1 0 29900 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _437_
timestamp 1701704242
transform -1 0 31004 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _438_
timestamp 1701704242
transform -1 0 31004 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _439_
timestamp 1701704242
transform 1 0 29532 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _440_
timestamp 1701704242
transform -1 0 27968 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _441_
timestamp 1701704242
transform 1 0 29348 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _442_
timestamp 1701704242
transform 1 0 28980 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _443_
timestamp 1701704242
transform 1 0 29532 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _444_
timestamp 1701704242
transform -1 0 27968 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _445_
timestamp 1701704242
transform -1 0 30820 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _446_
timestamp 1701704242
transform 1 0 29624 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _447_
timestamp 1701704242
transform -1 0 28520 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _448_
timestamp 1701704242
transform -1 0 28152 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _449_
timestamp 1701704242
transform -1 0 27600 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _450_
timestamp 1701704242
transform -1 0 26772 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp 1701704242
transform -1 0 26128 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _452_
timestamp 1701704242
transform -1 0 26312 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _453_
timestamp 1701704242
transform -1 0 25300 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _454_
timestamp 1701704242
transform -1 0 24288 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _455_
timestamp 1701704242
transform -1 0 20884 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _456_
timestamp 1701704242
transform 1 0 23000 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _457_
timestamp 1701704242
transform -1 0 20608 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _458_
timestamp 1701704242
transform 1 0 21252 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _459_
timestamp 1701704242
transform -1 0 22448 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _460_
timestamp 1701704242
transform 1 0 22448 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _461_
timestamp 1701704242
transform 1 0 21620 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _462_
timestamp 1701704242
transform -1 0 20884 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _463_
timestamp 1701704242
transform -1 0 21068 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _464_
timestamp 1701704242
transform -1 0 22724 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _465_
timestamp 1701704242
transform 1 0 22264 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _466_
timestamp 1701704242
transform 1 0 22080 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _467_
timestamp 1701704242
transform -1 0 23276 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _468_
timestamp 1701704242
transform -1 0 26772 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _469_
timestamp 1701704242
transform -1 0 26036 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _470_
timestamp 1701704242
transform -1 0 28428 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _471_
timestamp 1701704242
transform -1 0 26680 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _472_
timestamp 1701704242
transform -1 0 29900 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _473_
timestamp 1701704242
transform 1 0 29348 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _474_
timestamp 1701704242
transform 1 0 29532 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _475_
timestamp 1701704242
transform 1 0 29532 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _476_
timestamp 1701704242
transform -1 0 30084 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _477_
timestamp 1701704242
transform -1 0 27876 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _478_
timestamp 1701704242
transform -1 0 26772 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _479_
timestamp 1701704242
transform -1 0 25300 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _480_
timestamp 1701704242
transform -1 0 27784 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _481_
timestamp 1701704242
transform 1 0 23552 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _482_
timestamp 1701704242
transform -1 0 24196 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _483_
timestamp 1701704242
transform -1 0 25300 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _484_
timestamp 1701704242
transform -1 0 22724 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _485_
timestamp 1701704242
transform 1 0 18952 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _486_
timestamp 1701704242
transform 1 0 16100 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _487_
timestamp 1701704242
transform 1 0 17112 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _488_
timestamp 1701704242
transform 1 0 16376 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _489_
timestamp 1701704242
transform -1 0 17940 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _490_
timestamp 1701704242
transform 1 0 17756 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _491_
timestamp 1701704242
transform 1 0 21712 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _492_
timestamp 1701704242
transform 1 0 22080 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _493_
timestamp 1701704242
transform 1 0 21896 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 1701704242
transform -1 0 17572 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _495_
timestamp 1701704242
transform 1 0 19320 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _496_
timestamp 1701704242
transform 1 0 20700 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _497_
timestamp 1701704242
transform 1 0 14628 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 1701704242
transform 1 0 19504 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 1701704242
transform 1 0 16192 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _500_
timestamp 1701704242
transform 1 0 16560 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _501_
timestamp 1701704242
transform 1 0 11960 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 1701704242
transform 1 0 14904 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 1701704242
transform 1 0 10856 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 1701704242
transform 1 0 11960 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _505_
timestamp 1701704242
transform 1 0 11868 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 1701704242
transform 1 0 14168 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 1701704242
transform 1 0 10396 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _508_
timestamp 1701704242
transform 1 0 9292 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 1701704242
transform 1 0 6992 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _510_
timestamp 1701704242
transform 1 0 9936 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _511_
timestamp 1701704242
transform 1 0 9844 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _512_
timestamp 1701704242
transform 1 0 9844 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _513_
timestamp 1701704242
transform 1 0 10028 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _514_
timestamp 1701704242
transform 1 0 10948 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _515_
timestamp 1701704242
transform 1 0 11500 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _516_
timestamp 1701704242
transform 1 0 13616 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _517_
timestamp 1701704242
transform 1 0 11960 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _518_
timestamp 1701704242
transform 1 0 14720 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _519_
timestamp 1701704242
transform 1 0 13156 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _520_
timestamp 1701704242
transform 1 0 13616 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _521_
timestamp 1701704242
transform 1 0 13616 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _522_
timestamp 1701704242
transform 1 0 14536 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _523_
timestamp 1701704242
transform 1 0 11132 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _524_
timestamp 1701704242
transform 1 0 9936 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _525_
timestamp 1701704242
transform 1 0 9660 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _526_
timestamp 1701704242
transform 1 0 8280 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _527_
timestamp 1701704242
transform 1 0 8004 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _528_
timestamp 1701704242
transform 1 0 6348 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _529_
timestamp 1701704242
transform 1 0 8372 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _530_
timestamp 1701704242
transform 1 0 3680 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _531_
timestamp 1701704242
transform 1 0 6440 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _532_
timestamp 1701704242
transform 1 0 4140 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _533_
timestamp 1701704242
transform 1 0 4968 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _534_
timestamp 1701704242
transform 1 0 2668 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _535_
timestamp 1701704242
transform 1 0 2760 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _536_
timestamp 1701704242
transform 1 0 1656 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _537_
timestamp 1701704242
transform 1 0 1656 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _538_
timestamp 1701704242
transform 1 0 1656 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _539_
timestamp 1701704242
transform 1 0 920 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _540_
timestamp 1701704242
transform 1 0 1288 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _541_
timestamp 1701704242
transform 1 0 1656 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _542_
timestamp 1701704242
transform 1 0 1840 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _543_
timestamp 1701704242
transform 1 0 1104 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _544_
timestamp 1701704242
transform 1 0 4232 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _545_
timestamp 1701704242
transform 1 0 2208 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _546_
timestamp 1701704242
transform 1 0 3312 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _547_
timestamp 1701704242
transform 1 0 3680 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _548_
timestamp 1701704242
transform 1 0 3404 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _549_
timestamp 1701704242
transform 1 0 4232 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _550_
timestamp 1701704242
transform 1 0 4876 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _551_
timestamp 1701704242
transform 1 0 4600 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _552_
timestamp 1701704242
transform 1 0 5796 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _553_
timestamp 1701704242
transform 1 0 6532 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _554_
timestamp 1701704242
transform 1 0 8372 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _555_
timestamp 1701704242
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _556_
timestamp 1701704242
transform 1 0 8372 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _557_
timestamp 1701704242
transform 1 0 7360 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _558_
timestamp 1701704242
transform 1 0 6624 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _559_
timestamp 1701704242
transform 1 0 8832 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _560_
timestamp 1701704242
transform 1 0 8372 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _561_
timestamp 1701704242
transform 1 0 7820 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _562_
timestamp 1701704242
transform 1 0 4416 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _563_
timestamp 1701704242
transform 1 0 4140 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _564_
timestamp 1701704242
transform 1 0 8924 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _565_
timestamp 1701704242
transform 1 0 6716 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _566_
timestamp 1701704242
transform -1 0 8280 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _567_
timestamp 1701704242
transform 1 0 10948 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _568_
timestamp 1701704242
transform 1 0 9568 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _569_
timestamp 1701704242
transform 1 0 10948 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _570_
timestamp 1701704242
transform 1 0 10948 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _571_
timestamp 1701704242
transform 1 0 9200 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _572_
timestamp 1701704242
transform 1 0 10580 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _573_
timestamp 1701704242
transform 1 0 7268 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _574_
timestamp 1701704242
transform 1 0 12144 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _575_
timestamp 1701704242
transform 1 0 5796 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _576_
timestamp 1701704242
transform 1 0 4416 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _577_
timestamp 1701704242
transform 1 0 3220 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _578_
timestamp 1701704242
transform 1 0 3496 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _579_
timestamp 1701704242
transform 1 0 1104 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _580_
timestamp 1701704242
transform 1 0 2116 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _581_
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _582_
timestamp 1701704242
transform 1 0 2024 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _583_
timestamp 1701704242
transform 1 0 3588 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _584_
timestamp 1701704242
transform 1 0 2760 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _585_
timestamp 1701704242
transform 1 0 3864 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _586_
timestamp 1701704242
transform 1 0 5336 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _587_
timestamp 1701704242
transform 1 0 5612 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _588_
timestamp 1701704242
transform 1 0 6532 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _589_
timestamp 1701704242
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _590_
timestamp 1701704242
transform 1 0 8004 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _591_
timestamp 1701704242
transform 1 0 7912 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _592_
timestamp 1701704242
transform 1 0 9568 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _593_
timestamp 1701704242
transform 1 0 9384 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _594_
timestamp 1701704242
transform 1 0 10764 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _595_
timestamp 1701704242
transform 1 0 11592 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _596_
timestamp 1701704242
transform 1 0 11224 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _597_
timestamp 1701704242
transform 1 0 11224 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _598_
timestamp 1701704242
transform 1 0 14536 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _599_
timestamp 1701704242
transform 1 0 13064 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _600_
timestamp 1701704242
transform 1 0 16100 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _601_
timestamp 1701704242
transform 1 0 13524 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _602_
timestamp 1701704242
transform 1 0 16560 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _603_
timestamp 1701704242
transform 1 0 15732 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _604_
timestamp 1701704242
transform 1 0 18676 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _605_
timestamp 1701704242
transform 1 0 18124 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _606_
timestamp 1701704242
transform -1 0 20148 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _607_
timestamp 1701704242
transform 1 0 20148 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _608_
timestamp 1701704242
transform 1 0 20332 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _609_
timestamp 1701704242
transform 1 0 22080 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _610_
timestamp 1701704242
transform -1 0 25208 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _611_
timestamp 1701704242
transform -1 0 23184 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _612_
timestamp 1701704242
transform -1 0 26588 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _613_
timestamp 1701704242
transform -1 0 25300 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _614_
timestamp 1701704242
transform 1 0 21896 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _615_
timestamp 1701704242
transform -1 0 26220 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _616_
timestamp 1701704242
transform -1 0 26036 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _617_
timestamp 1701704242
transform -1 0 28888 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _618_
timestamp 1701704242
transform -1 0 28060 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _619_
timestamp 1701704242
transform -1 0 28060 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _620_
timestamp 1701704242
transform 1 0 29532 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _621_
timestamp 1701704242
transform -1 0 30912 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _638_
timestamp 1701704242
transform -1 0 25576 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16100 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 7360 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1701704242
transform -1 0 7360 0 -1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1701704242
transform -1 0 12144 0 -1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1701704242
transform 1 0 10396 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1701704242
transform 1 0 6440 0 1 12512
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1701704242
transform 1 0 7268 0 -1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1701704242
transform 1 0 12144 0 -1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1701704242
transform -1 0 12696 0 1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1701704242
transform -1 0 21988 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1701704242
transform -1 0 23736 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1701704242
transform -1 0 26312 0 -1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1701704242
transform 1 0 26404 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1701704242
transform -1 0 22264 0 -1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1701704242
transform 1 0 19780 0 -1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1701704242
transform 1 0 26772 0 1 12512
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1701704242
transform 1 0 25300 0 -1 13600
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1701704242
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1701704242
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1701704242
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_88 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8648 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_94
timestamp 1701704242
transform 1 0 9200 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_98 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 9568 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_103 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10028 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1701704242
transform 1 0 10764 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1701704242
transform 1 0 10948 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_121
timestamp 1701704242
transform 1 0 11684 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_129
timestamp 1701704242
transform 1 0 12420 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_134
timestamp 1701704242
transform 1 0 12880 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp 1701704242
transform 1 0 13248 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1701704242
transform 1 0 13524 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1701704242
transform 1 0 14260 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_156
timestamp 1701704242
transform 1 0 14904 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_162
timestamp 1701704242
transform 1 0 15456 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1701704242
transform 1 0 15916 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1701704242
transform 1 0 18492 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_213 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 20148 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_217
timestamp 1701704242
transform 1 0 20516 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1701704242
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_250
timestamp 1701704242
transform 1 0 23552 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_262
timestamp 1701704242
transform 1 0 24656 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_274
timestamp 1701704242
transform 1 0 25760 0 1 544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1701704242
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1701704242
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1701704242
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1701704242
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_321
timestamp 1701704242
transform 1 0 30084 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1701704242
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1701704242
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1701704242
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_69
timestamp 1701704242
transform 1 0 6900 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_156
timestamp 1701704242
transform 1 0 14904 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_164
timestamp 1701704242
transform 1 0 15640 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1701704242
transform 1 0 16100 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_174
timestamp 1701704242
transform 1 0 16560 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_246
timestamp 1701704242
transform 1 0 23184 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_251
timestamp 1701704242
transform 1 0 23644 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_268
timestamp 1701704242
transform 1 0 25208 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_272
timestamp 1701704242
transform 1 0 25576 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1701704242
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1701704242
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1701704242
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1701704242
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_329
timestamp 1701704242
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1701704242
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_15
timestamp 1701704242
transform 1 0 1932 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_21
timestamp 1701704242
transform 1 0 2484 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25
timestamp 1701704242
transform 1 0 2852 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_32
timestamp 1701704242
transform 1 0 3496 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_77
timestamp 1701704242
transform 1 0 7636 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_88
timestamp 1701704242
transform 1 0 8648 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_94
timestamp 1701704242
transform 1 0 9200 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_101
timestamp 1701704242
transform 1 0 9844 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_109
timestamp 1701704242
transform 1 0 10580 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1701704242
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1701704242
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_141
timestamp 1701704242
transform 1 0 13524 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_149
timestamp 1701704242
transform 1 0 14260 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_153
timestamp 1701704242
transform 1 0 14628 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_174
timestamp 1701704242
transform 1 0 16560 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_185
timestamp 1701704242
transform 1 0 17572 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1701704242
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_197
timestamp 1701704242
transform 1 0 18676 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_205
timestamp 1701704242
transform 1 0 19412 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_214
timestamp 1701704242
transform 1 0 20240 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_234
timestamp 1701704242
transform 1 0 22080 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_246
timestamp 1701704242
transform 1 0 23184 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_265
timestamp 1701704242
transform 1 0 24932 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_283
timestamp 1701704242
transform 1 0 26588 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_295
timestamp 1701704242
transform 1 0 27692 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1701704242
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1701704242
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1701704242
transform 1 0 30084 0 1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_15
timestamp 1701704242
transform 1 0 1932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_43
timestamp 1701704242
transform 1 0 4508 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_47
timestamp 1701704242
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 1701704242
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_69
timestamp 1701704242
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_75
timestamp 1701704242
transform 1 0 7452 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_79
timestamp 1701704242
transform 1 0 7820 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_113
timestamp 1701704242
transform 1 0 10948 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_119
timestamp 1701704242
transform 1 0 11500 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_169
timestamp 1701704242
transform 1 0 16100 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_173
timestamp 1701704242
transform 1 0 16468 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_190
timestamp 1701704242
transform 1 0 18032 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_207
timestamp 1701704242
transform 1 0 19596 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_216
timestamp 1701704242
transform 1 0 20424 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_225
timestamp 1701704242
transform 1 0 21252 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_229
timestamp 1701704242
transform 1 0 21620 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_246
timestamp 1701704242
transform 1 0 23184 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_260
timestamp 1701704242
transform 1 0 24472 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_281
timestamp 1701704242
transform 1 0 26404 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_288
timestamp 1701704242
transform 1 0 27048 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_295
timestamp 1701704242
transform 1 0 27692 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_307
timestamp 1701704242
transform 1 0 28796 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_319
timestamp 1701704242
transform 1 0 29900 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_327
timestamp 1701704242
transform 1 0 30636 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_11
timestamp 1701704242
transform 1 0 1564 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_18
timestamp 1701704242
transform 1 0 2208 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_35
timestamp 1701704242
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_97
timestamp 1701704242
transform 1 0 9476 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_114
timestamp 1701704242
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_132
timestamp 1701704242
transform 1 0 12696 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1701704242
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_157
timestamp 1701704242
transform 1 0 14996 0 1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_181
timestamp 1701704242
transform 1 0 17204 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1701704242
transform 1 0 18308 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_229
timestamp 1701704242
transform 1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_248
timestamp 1701704242
transform 1 0 23368 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_281
timestamp 1701704242
transform 1 0 26404 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_291
timestamp 1701704242
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_312
timestamp 1701704242
transform 1 0 29256 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_321
timestamp 1701704242
transform 1 0 30084 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_7
timestamp 1701704242
transform 1 0 1196 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_23
timestamp 1701704242
transform 1 0 2668 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_40
timestamp 1701704242
transform 1 0 4232 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 1701704242
transform 1 0 5336 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_97
timestamp 1701704242
transform 1 0 9476 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1701704242
transform 1 0 10580 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1701704242
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_125
timestamp 1701704242
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_129
timestamp 1701704242
transform 1 0 12420 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_145
timestamp 1701704242
transform 1 0 13892 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_163
timestamp 1701704242
transform 1 0 15548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_169
timestamp 1701704242
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_176
timestamp 1701704242
transform 1 0 16744 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_184
timestamp 1701704242
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_196
timestamp 1701704242
transform 1 0 18584 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_209
timestamp 1701704242
transform 1 0 19780 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_215
timestamp 1701704242
transform 1 0 20332 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1701704242
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_235
timestamp 1701704242
transform 1 0 22172 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_252
timestamp 1701704242
transform 1 0 23736 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_260
timestamp 1701704242
transform 1 0 24472 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_277
timestamp 1701704242
transform 1 0 26036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_281
timestamp 1701704242
transform 1 0 26404 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_288
timestamp 1701704242
transform 1 0 27048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_298
timestamp 1701704242
transform 1 0 27968 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_311
timestamp 1701704242
transform 1 0 29164 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_331
timestamp 1701704242
transform 1 0 31004 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_24
timestamp 1701704242
transform 1 0 2760 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_29
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_49
timestamp 1701704242
transform 1 0 5060 0 1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_71
timestamp 1701704242
transform 1 0 7084 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1701704242
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_97
timestamp 1701704242
transform 1 0 9476 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_114
timestamp 1701704242
transform 1 0 11040 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_118
timestamp 1701704242
transform 1 0 11408 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_124
timestamp 1701704242
transform 1 0 11960 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_136
timestamp 1701704242
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_141
timestamp 1701704242
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_154
timestamp 1701704242
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_166
timestamp 1701704242
transform 1 0 15824 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_193
timestamp 1701704242
transform 1 0 18308 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1701704242
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_209
timestamp 1701704242
transform 1 0 19780 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_219
timestamp 1701704242
transform 1 0 20700 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_227
timestamp 1701704242
transform 1 0 21436 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_233
timestamp 1701704242
transform 1 0 21988 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_249
timestamp 1701704242
transform 1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_279
timestamp 1701704242
transform 1 0 26220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_299
timestamp 1701704242
transform 1 0 28060 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_306
timestamp 1701704242
transform 1 0 28704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_330
timestamp 1701704242
transform 1 0 30912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_15
timestamp 1701704242
transform 1 0 1932 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_48
timestamp 1701704242
transform 1 0 4968 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_89
timestamp 1701704242
transform 1 0 8740 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_93
timestamp 1701704242
transform 1 0 9108 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1701704242
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_113
timestamp 1701704242
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_131
timestamp 1701704242
transform 1 0 12604 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_148
timestamp 1701704242
transform 1 0 14168 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_154
timestamp 1701704242
transform 1 0 14720 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1701704242
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_169
timestamp 1701704242
transform 1 0 16100 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_185
timestamp 1701704242
transform 1 0 17572 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_197
timestamp 1701704242
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_208
timestamp 1701704242
transform 1 0 19688 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_225
timestamp 1701704242
transform 1 0 21252 0 -1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_245
timestamp 1701704242
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_257
timestamp 1701704242
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_269
timestamp 1701704242
transform 1 0 25300 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_277
timestamp 1701704242
transform 1 0 26036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_281
timestamp 1701704242
transform 1 0 26404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_299
timestamp 1701704242
transform 1 0 28060 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_305
timestamp 1701704242
transform 1 0 28612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_312
timestamp 1701704242
transform 1 0 29256 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_330
timestamp 1701704242
transform 1 0 30912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_7
timestamp 1701704242
transform 1 0 1196 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1701704242
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_42
timestamp 1701704242
transform 1 0 4416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1701704242
transform 1 0 8372 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_107
timestamp 1701704242
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_125
timestamp 1701704242
transform 1 0 12052 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_133
timestamp 1701704242
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_141
timestamp 1701704242
transform 1 0 13524 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_152
timestamp 1701704242
transform 1 0 14536 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_156
timestamp 1701704242
transform 1 0 14904 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_173
timestamp 1701704242
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_187
timestamp 1701704242
transform 1 0 17756 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1701704242
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_202
timestamp 1701704242
transform 1 0 19136 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_223
timestamp 1701704242
transform 1 0 21068 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_235
timestamp 1701704242
transform 1 0 22172 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_247
timestamp 1701704242
transform 1 0 23276 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1701704242
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_285
timestamp 1701704242
transform 1 0 26772 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_297
timestamp 1701704242
transform 1 0 27876 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_301
timestamp 1701704242
transform 1 0 28244 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_331
timestamp 1701704242
transform 1 0 31004 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_22
timestamp 1701704242
transform 1 0 2576 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_45
timestamp 1701704242
transform 1 0 4692 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_52
timestamp 1701704242
transform 1 0 5336 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_76
timestamp 1701704242
transform 1 0 7544 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_80
timestamp 1701704242
transform 1 0 7912 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_92
timestamp 1701704242
transform 1 0 9016 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_96
timestamp 1701704242
transform 1 0 9384 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_103
timestamp 1701704242
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_108
timestamp 1701704242
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1701704242
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_142
timestamp 1701704242
transform 1 0 13616 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_150
timestamp 1701704242
transform 1 0 14352 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_159
timestamp 1701704242
transform 1 0 15180 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1701704242
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_169
timestamp 1701704242
transform 1 0 16100 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_195
timestamp 1701704242
transform 1 0 18492 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 1701704242
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_241
timestamp 1701704242
transform 1 0 22724 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_252
timestamp 1701704242
transform 1 0 23736 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_256
timestamp 1701704242
transform 1 0 24104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_265
timestamp 1701704242
transform 1 0 24932 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_272
timestamp 1701704242
transform 1 0 25576 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_284
timestamp 1701704242
transform 1 0 26680 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_307
timestamp 1701704242
transform 1 0 28796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_312
timestamp 1701704242
transform 1 0 29256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 1701704242
transform 1 0 828 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1701704242
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_35
timestamp 1701704242
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_58
timestamp 1701704242
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_63
timestamp 1701704242
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_67
timestamp 1701704242
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_103
timestamp 1701704242
transform 1 0 10028 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_129
timestamp 1701704242
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 1701704242
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_155
timestamp 1701704242
transform 1 0 14812 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_161
timestamp 1701704242
transform 1 0 15364 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_168
timestamp 1701704242
transform 1 0 16008 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_184
timestamp 1701704242
transform 1 0 17480 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1701704242
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_203
timestamp 1701704242
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_221
timestamp 1701704242
transform 1 0 20884 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1701704242
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_304
timestamp 1701704242
transform 1 0 28520 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_309
timestamp 1701704242
transform 1 0 28980 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_15
timestamp 1701704242
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_33
timestamp 1701704242
transform 1 0 3588 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 1701704242
transform 1 0 4692 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1701704242
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_80
timestamp 1701704242
transform 1 0 7912 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_90
timestamp 1701704242
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_98
timestamp 1701704242
transform 1 0 9568 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1701704242
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_129
timestamp 1701704242
transform 1 0 12420 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_135
timestamp 1701704242
transform 1 0 12972 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_145
timestamp 1701704242
transform 1 0 13892 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_163
timestamp 1701704242
transform 1 0 15548 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1701704242
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 1701704242
transform 1 0 16100 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_177
timestamp 1701704242
transform 1 0 16836 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_181
timestamp 1701704242
transform 1 0 17204 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_203
timestamp 1701704242
transform 1 0 19228 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_209
timestamp 1701704242
transform 1 0 19780 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_221
timestamp 1701704242
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_225
timestamp 1701704242
transform 1 0 21252 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_240
timestamp 1701704242
transform 1 0 22632 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_258
timestamp 1701704242
transform 1 0 24288 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_270
timestamp 1701704242
transform 1 0 25392 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_276
timestamp 1701704242
transform 1 0 25944 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_298
timestamp 1701704242
transform 1 0 27968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_302
timestamp 1701704242
transform 1 0 28336 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_309
timestamp 1701704242
transform 1 0 28980 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_313
timestamp 1701704242
transform 1 0 29348 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_323
timestamp 1701704242
transform 1 0 30268 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_330
timestamp 1701704242
transform 1 0 30912 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_3
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_22
timestamp 1701704242
transform 1 0 2576 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_37
timestamp 1701704242
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1701704242
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_85
timestamp 1701704242
transform 1 0 8372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_123
timestamp 1701704242
transform 1 0 11868 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_131
timestamp 1701704242
transform 1 0 12604 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1701704242
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 1701704242
transform 1 0 13524 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_145
timestamp 1701704242
transform 1 0 13892 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_155
timestamp 1701704242
transform 1 0 14812 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_170
timestamp 1701704242
transform 1 0 16192 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_177
timestamp 1701704242
transform 1 0 16836 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_184
timestamp 1701704242
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_192
timestamp 1701704242
transform 1 0 18216 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp 1701704242
transform 1 0 18676 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp 1701704242
transform 1 0 19044 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_218
timestamp 1701704242
transform 1 0 20608 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_240
timestamp 1701704242
transform 1 0 22632 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_253
timestamp 1701704242
transform 1 0 23828 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_261
timestamp 1701704242
transform 1 0 24564 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_294
timestamp 1701704242
transform 1 0 27600 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_300
timestamp 1701704242
transform 1 0 28152 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1701704242
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_315
timestamp 1701704242
transform 1 0 29532 0 1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1701704242
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_15
timestamp 1701704242
transform 1 0 1932 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_50
timestamp 1701704242
transform 1 0 5152 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_77
timestamp 1701704242
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_95
timestamp 1701704242
transform 1 0 9292 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_107
timestamp 1701704242
transform 1 0 10396 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1701704242
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_143
timestamp 1701704242
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_151
timestamp 1701704242
transform 1 0 14444 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_163
timestamp 1701704242
transform 1 0 15548 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1701704242
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_180
timestamp 1701704242
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_188
timestamp 1701704242
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_201
timestamp 1701704242
transform 1 0 19044 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_219
timestamp 1701704242
transform 1 0 20700 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1701704242
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_225
timestamp 1701704242
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_241
timestamp 1701704242
transform 1 0 22724 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_260
timestamp 1701704242
transform 1 0 24472 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_268
timestamp 1701704242
transform 1 0 25208 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_281
timestamp 1701704242
transform 1 0 26404 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_300
timestamp 1701704242
transform 1 0 28152 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_313
timestamp 1701704242
transform 1 0 29348 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_331
timestamp 1701704242
transform 1 0 31004 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_14
timestamp 1701704242
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 1701704242
transform 1 0 2852 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_41
timestamp 1701704242
transform 1 0 4324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_58
timestamp 1701704242
transform 1 0 5888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_79
timestamp 1701704242
transform 1 0 7820 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1701704242
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_101
timestamp 1701704242
transform 1 0 9844 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_123
timestamp 1701704242
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_136
timestamp 1701704242
transform 1 0 13064 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_155
timestamp 1701704242
transform 1 0 14812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_171
timestamp 1701704242
transform 1 0 16284 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_187
timestamp 1701704242
transform 1 0 17756 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1701704242
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_197
timestamp 1701704242
transform 1 0 18676 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_214
timestamp 1701704242
transform 1 0 20240 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_238
timestamp 1701704242
transform 1 0 22448 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_246
timestamp 1701704242
transform 1 0 23184 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_262
timestamp 1701704242
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_280
timestamp 1701704242
transform 1 0 26312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_298
timestamp 1701704242
transform 1 0 27968 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_304
timestamp 1701704242
transform 1 0 28520 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_330
timestamp 1701704242
transform 1 0 30912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_3
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_16
timestamp 1701704242
transform 1 0 2024 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_20
timestamp 1701704242
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1701704242
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_81
timestamp 1701704242
transform 1 0 8004 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_89
timestamp 1701704242
transform 1 0 8740 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_106
timestamp 1701704242
transform 1 0 10304 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1701704242
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_125
timestamp 1701704242
transform 1 0 12052 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_133
timestamp 1701704242
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_142
timestamp 1701704242
transform 1 0 13616 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_159
timestamp 1701704242
transform 1 0 15180 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1701704242
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_177
timestamp 1701704242
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_198
timestamp 1701704242
transform 1 0 18768 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_218
timestamp 1701704242
transform 1 0 20608 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_225
timestamp 1701704242
transform 1 0 21252 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_237
timestamp 1701704242
transform 1 0 22356 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_263
timestamp 1701704242
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_274
timestamp 1701704242
transform 1 0 25760 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_281
timestamp 1701704242
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_298
timestamp 1701704242
transform 1 0 27968 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_314
timestamp 1701704242
transform 1 0 29440 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_331
timestamp 1701704242
transform 1 0 31004 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_22
timestamp 1701704242
transform 1 0 2576 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3220 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_33
timestamp 1701704242
transform 1 0 3588 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_43
timestamp 1701704242
transform 1 0 4508 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_63
timestamp 1701704242
transform 1 0 6348 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_101
timestamp 1701704242
transform 1 0 9844 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_109
timestamp 1701704242
transform 1 0 10580 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1701704242
transform 1 0 13156 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_150
timestamp 1701704242
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_164
timestamp 1701704242
transform 1 0 15640 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1701704242
transform 1 0 17940 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1701704242
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 1701704242
transform 1 0 18676 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp 1701704242
transform 1 0 19044 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_225
timestamp 1701704242
transform 1 0 21252 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_229
timestamp 1701704242
transform 1 0 21620 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_242
timestamp 1701704242
transform 1 0 22816 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1701704242
transform 1 0 23552 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_253
timestamp 1701704242
transform 1 0 23828 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_290
timestamp 1701704242
transform 1 0 27232 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_302
timestamp 1701704242
transform 1 0 28336 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_318
timestamp 1701704242
transform 1 0 29808 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_328
timestamp 1701704242
transform 1 0 30728 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_13
timestamp 1701704242
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_48
timestamp 1701704242
transform 1 0 4968 0 -1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1701704242
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_69
timestamp 1701704242
transform 1 0 6900 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_78
timestamp 1701704242
transform 1 0 7728 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_90
timestamp 1701704242
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_94
timestamp 1701704242
transform 1 0 9200 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1701704242
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_113
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_121
timestamp 1701704242
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_144
timestamp 1701704242
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_164
timestamp 1701704242
transform 1 0 15640 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1701704242
transform 1 0 21068 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_225
timestamp 1701704242
transform 1 0 21252 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_245
timestamp 1701704242
transform 1 0 23092 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_255
timestamp 1701704242
transform 1 0 24012 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_275
timestamp 1701704242
transform 1 0 25852 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1701704242
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_281
timestamp 1701704242
transform 1 0 26404 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_285
timestamp 1701704242
transform 1 0 26772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_302
timestamp 1701704242
transform 1 0 28336 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_9
timestamp 1701704242
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_19
timestamp 1701704242
transform 1 0 2300 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1701704242
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1701704242
transform 1 0 3220 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1701704242
transform 1 0 3956 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_41
timestamp 1701704242
transform 1 0 4324 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_47
timestamp 1701704242
transform 1 0 4876 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_55
timestamp 1701704242
transform 1 0 5612 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_63
timestamp 1701704242
transform 1 0 6348 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1701704242
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_92
timestamp 1701704242
transform 1 0 9016 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_99
timestamp 1701704242
transform 1 0 9660 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_103
timestamp 1701704242
transform 1 0 10028 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_107
timestamp 1701704242
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_112
timestamp 1701704242
transform 1 0 10856 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_124
timestamp 1701704242
transform 1 0 11960 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp 1701704242
transform 1 0 12972 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1701704242
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp 1701704242
transform 1 0 13524 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_180
timestamp 1701704242
transform 1 0 17112 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_187
timestamp 1701704242
transform 1 0 17756 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_201
timestamp 1701704242
transform 1 0 19044 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_207
timestamp 1701704242
transform 1 0 19596 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_216
timestamp 1701704242
transform 1 0 20424 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_224
timestamp 1701704242
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_235
timestamp 1701704242
transform 1 0 22172 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1701704242
transform 1 0 23828 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_304
timestamp 1701704242
transform 1 0 28520 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_309
timestamp 1701704242
transform 1 0 28980 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_319
timestamp 1701704242
transform 1 0 29900 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_7
timestamp 1701704242
transform 1 0 1196 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_24
timestamp 1701704242
transform 1 0 2760 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_46
timestamp 1701704242
transform 1 0 4784 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_65
timestamp 1701704242
transform 1 0 6532 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_69
timestamp 1701704242
transform 1 0 6900 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_93
timestamp 1701704242
transform 1 0 9108 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1701704242
transform 1 0 10948 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_120
timestamp 1701704242
transform 1 0 11592 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_133
timestamp 1701704242
transform 1 0 12788 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_145
timestamp 1701704242
transform 1 0 13892 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_164
timestamp 1701704242
transform 1 0 15640 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_201
timestamp 1701704242
transform 1 0 19044 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_221
timestamp 1701704242
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_260
timestamp 1701704242
transform 1 0 24472 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_268
timestamp 1701704242
transform 1 0 25208 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_274
timestamp 1701704242
transform 1 0 25760 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_281
timestamp 1701704242
transform 1 0 26404 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_285
timestamp 1701704242
transform 1 0 26772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_313
timestamp 1701704242
transform 1 0 29348 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_331
timestamp 1701704242
transform 1 0 31004 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_29
timestamp 1701704242
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_47
timestamp 1701704242
transform 1 0 4876 0 1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_63
timestamp 1701704242
transform 1 0 6348 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1701704242
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 1701704242
transform 1 0 8372 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_91
timestamp 1701704242
transform 1 0 8924 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_101
timestamp 1701704242
transform 1 0 9844 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_118
timestamp 1701704242
transform 1 0 11408 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_148
timestamp 1701704242
transform 1 0 14168 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_152
timestamp 1701704242
transform 1 0 14536 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_161
timestamp 1701704242
transform 1 0 15364 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_173
timestamp 1701704242
transform 1 0 16468 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_180
timestamp 1701704242
transform 1 0 17112 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_188
timestamp 1701704242
transform 1 0 17848 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_233
timestamp 1701704242
transform 1 0 21988 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_253
timestamp 1701704242
transform 1 0 23828 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_294
timestamp 1701704242
transform 1 0 27600 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_300
timestamp 1701704242
transform 1 0 28152 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1701704242
transform 1 0 28796 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_331
timestamp 1701704242
transform 1 0 31004 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_3
timestamp 1701704242
transform 1 0 828 0 -1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_18
timestamp 1701704242
transform 1 0 2208 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_30
timestamp 1701704242
transform 1 0 3312 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_39
timestamp 1701704242
transform 1 0 4140 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1701704242
transform 1 0 5796 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_69
timestamp 1701704242
transform 1 0 6900 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_73
timestamp 1701704242
transform 1 0 7268 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_90
timestamp 1701704242
transform 1 0 8832 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_94
timestamp 1701704242
transform 1 0 9200 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1701704242
transform 1 0 10396 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1701704242
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_113
timestamp 1701704242
transform 1 0 10948 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_121
timestamp 1701704242
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_129
timestamp 1701704242
transform 1 0 12420 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_140
timestamp 1701704242
transform 1 0 13432 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_152
timestamp 1701704242
transform 1 0 14536 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_169
timestamp 1701704242
transform 1 0 16100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_173
timestamp 1701704242
transform 1 0 16468 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_191
timestamp 1701704242
transform 1 0 18124 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_221
timestamp 1701704242
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1701704242
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_237
timestamp 1701704242
transform 1 0 22356 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_252
timestamp 1701704242
transform 1 0 23736 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_272
timestamp 1701704242
transform 1 0 25576 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_281
timestamp 1701704242
transform 1 0 26404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_285
timestamp 1701704242
transform 1 0 26772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_302
timestamp 1701704242
transform 1 0 28336 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_322
timestamp 1701704242
transform 1 0 30176 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_330
timestamp 1701704242
transform 1 0 30912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_3
timestamp 1701704242
transform 1 0 828 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_11
timestamp 1701704242
transform 1 0 1564 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_29
timestamp 1701704242
transform 1 0 3220 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_37
timestamp 1701704242
transform 1 0 3956 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_47
timestamp 1701704242
transform 1 0 4876 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_55
timestamp 1701704242
transform 1 0 5612 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_75
timestamp 1701704242
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1701704242
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1701704242
transform 1 0 8372 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_93
timestamp 1701704242
transform 1 0 9108 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_100
timestamp 1701704242
transform 1 0 9752 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_117
timestamp 1701704242
transform 1 0 11316 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_121
timestamp 1701704242
transform 1 0 11684 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_130
timestamp 1701704242
transform 1 0 12512 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_134
timestamp 1701704242
transform 1 0 12880 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_150
timestamp 1701704242
transform 1 0 14352 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_172
timestamp 1701704242
transform 1 0 16376 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_178
timestamp 1701704242
transform 1 0 16928 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_192
timestamp 1701704242
transform 1 0 18216 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_201
timestamp 1701704242
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_247
timestamp 1701704242
transform 1 0 23276 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1701704242
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_253
timestamp 1701704242
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_258
timestamp 1701704242
transform 1 0 24288 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_268
timestamp 1701704242
transform 1 0 25208 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_296
timestamp 1701704242
transform 1 0 27784 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_312
timestamp 1701704242
transform 1 0 29256 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_329
timestamp 1701704242
transform 1 0 30820 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1701704242
transform 1 0 828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_11
timestamp 1701704242
transform 1 0 1564 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_28
timestamp 1701704242
transform 1 0 3128 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_36
timestamp 1701704242
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp 1701704242
transform 1 0 5336 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_87
timestamp 1701704242
transform 1 0 8556 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_95
timestamp 1701704242
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_106
timestamp 1701704242
transform 1 0 10304 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1701704242
transform 1 0 10948 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_117
timestamp 1701704242
transform 1 0 11316 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_146
timestamp 1701704242
transform 1 0 13984 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_156
timestamp 1701704242
transform 1 0 14904 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_169
timestamp 1701704242
transform 1 0 16100 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_184
timestamp 1701704242
transform 1 0 17480 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_193
timestamp 1701704242
transform 1 0 18308 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_197
timestamp 1701704242
transform 1 0 18676 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_220
timestamp 1701704242
transform 1 0 20792 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_231
timestamp 1701704242
transform 1 0 21804 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_250
timestamp 1701704242
transform 1 0 23552 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_258
timestamp 1701704242
transform 1 0 24288 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_319
timestamp 1701704242
transform 1 0 29900 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_331
timestamp 1701704242
transform 1 0 31004 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_3
timestamp 1701704242
transform 1 0 828 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1701704242
transform 1 0 3220 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_49
timestamp 1701704242
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_54
timestamp 1701704242
transform 1 0 5520 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_61
timestamp 1701704242
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_72
timestamp 1701704242
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1701704242
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_117
timestamp 1701704242
transform 1 0 11316 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1701704242
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_152
timestamp 1701704242
transform 1 0 14536 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_168
timestamp 1701704242
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_175
timestamp 1701704242
transform 1 0 16652 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_179
timestamp 1701704242
transform 1 0 17020 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_185
timestamp 1701704242
transform 1 0 17572 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 1701704242
transform 1 0 18308 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_237
timestamp 1701704242
transform 1 0 22356 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_250
timestamp 1701704242
transform 1 0 23552 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_258
timestamp 1701704242
transform 1 0 24288 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_280
timestamp 1701704242
transform 1 0 26312 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_299
timestamp 1701704242
transform 1 0 28060 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1701704242
transform 1 0 28796 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_315
timestamp 1701704242
transform 1 0 29532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_327
timestamp 1701704242
transform 1 0 30636 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_331
timestamp 1701704242
transform 1 0 31004 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_3
timestamp 1701704242
transform 1 0 828 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_22
timestamp 1701704242
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_40
timestamp 1701704242
transform 1 0 4232 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_50
timestamp 1701704242
transform 1 0 5152 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_60
timestamp 1701704242
transform 1 0 6072 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_64
timestamp 1701704242
transform 1 0 6440 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1701704242
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_93
timestamp 1701704242
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1701704242
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_132
timestamp 1701704242
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_151
timestamp 1701704242
transform 1 0 14444 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_163
timestamp 1701704242
transform 1 0 15548 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1701704242
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1701704242
transform 1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_173
timestamp 1701704242
transform 1 0 16468 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_190
timestamp 1701704242
transform 1 0 18032 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_202
timestamp 1701704242
transform 1 0 19136 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_222
timestamp 1701704242
transform 1 0 20976 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_241
timestamp 1701704242
transform 1 0 22724 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_252
timestamp 1701704242
transform 1 0 23736 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_267
timestamp 1701704242
transform 1 0 25116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1701704242
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_287
timestamp 1701704242
transform 1 0 26956 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_331
timestamp 1701704242
transform 1 0 31004 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp 1701704242
transform 1 0 828 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_20
timestamp 1701704242
transform 1 0 2392 0 1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1701704242
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_41
timestamp 1701704242
transform 1 0 4324 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_60
timestamp 1701704242
transform 1 0 6072 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 1701704242
transform 1 0 8372 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_93
timestamp 1701704242
transform 1 0 9108 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_119
timestamp 1701704242
transform 1 0 11500 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_123
timestamp 1701704242
transform 1 0 11868 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_141
timestamp 1701704242
transform 1 0 13524 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_168
timestamp 1701704242
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1701704242
transform 1 0 18308 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_204
timestamp 1701704242
transform 1 0 19320 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_216
timestamp 1701704242
transform 1 0 20424 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_235
timestamp 1701704242
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_247
timestamp 1701704242
transform 1 0 23276 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1701704242
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_261
timestamp 1701704242
transform 1 0 24564 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_267
timestamp 1701704242
transform 1 0 25116 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_284
timestamp 1701704242
transform 1 0 26680 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_296
timestamp 1701704242
transform 1 0 27784 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1701704242
transform 1 0 30084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_329
timestamp 1701704242
transform 1 0 30820 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_3
timestamp 1701704242
transform 1 0 828 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_21
timestamp 1701704242
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1701704242
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_57
timestamp 1701704242
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_63
timestamp 1701704242
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_80
timestamp 1701704242
transform 1 0 7912 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_92
timestamp 1701704242
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1701704242
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 1701704242
transform 1 0 10948 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_135
timestamp 1701704242
transform 1 0 12972 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_141
timestamp 1701704242
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_164
timestamp 1701704242
transform 1 0 15640 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_169
timestamp 1701704242
transform 1 0 16100 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_187
timestamp 1701704242
transform 1 0 17756 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_203
timestamp 1701704242
transform 1 0 19228 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1701704242
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_225
timestamp 1701704242
transform 1 0 21252 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_231
timestamp 1701704242
transform 1 0 21804 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_248
timestamp 1701704242
transform 1 0 23368 0 -1 15776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_264
timestamp 1701704242
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_276
timestamp 1701704242
transform 1 0 25944 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_297
timestamp 1701704242
transform 1 0 27876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_314
timestamp 1701704242
transform 1 0 29440 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_331
timestamp 1701704242
transform 1 0 31004 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_3
timestamp 1701704242
transform 1 0 828 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_9
timestamp 1701704242
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 1701704242
transform 1 0 3220 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_36
timestamp 1701704242
transform 1 0 3864 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_64
timestamp 1701704242
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_76
timestamp 1701704242
transform 1 0 7544 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_116
timestamp 1701704242
transform 1 0 11224 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_120
timestamp 1701704242
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1701704242
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_185
timestamp 1701704242
transform 1 0 17572 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_193
timestamp 1701704242
transform 1 0 18308 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_209
timestamp 1701704242
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_229
timestamp 1701704242
transform 1 0 21620 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_233
timestamp 1701704242
transform 1 0 21988 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1701704242
transform 1 0 23552 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_288
timestamp 1701704242
transform 1 0 27048 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_292
timestamp 1701704242
transform 1 0 27416 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_315
timestamp 1701704242
transform 1 0 29532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_327
timestamp 1701704242
transform 1 0 30636 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_331
timestamp 1701704242
transform 1 0 31004 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1701704242
transform 1 0 828 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_11
timestamp 1701704242
transform 1 0 1564 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_17
timestamp 1701704242
transform 1 0 2116 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_44
timestamp 1701704242
transform 1 0 4600 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_48
timestamp 1701704242
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_79
timestamp 1701704242
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_97
timestamp 1701704242
transform 1 0 9476 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_103
timestamp 1701704242
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_107
timestamp 1701704242
transform 1 0 10396 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1701704242
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_113
timestamp 1701704242
transform 1 0 10948 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_120
timestamp 1701704242
transform 1 0 11592 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_124
timestamp 1701704242
transform 1 0 11960 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_131
timestamp 1701704242
transform 1 0 12604 0 -1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_153
timestamp 1701704242
transform 1 0 14628 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1701704242
transform 1 0 15732 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1701704242
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_181
timestamp 1701704242
transform 1 0 17204 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_203
timestamp 1701704242
transform 1 0 19228 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_207
timestamp 1701704242
transform 1 0 19596 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_217
timestamp 1701704242
transform 1 0 20516 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1701704242
transform 1 0 20976 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1701704242
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_249
timestamp 1701704242
transform 1 0 23460 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_266
timestamp 1701704242
transform 1 0 25024 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1701704242
transform 1 0 26128 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_281
timestamp 1701704242
transform 1 0 26404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_300
timestamp 1701704242
transform 1 0 28152 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_304
timestamp 1701704242
transform 1 0 28520 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_321
timestamp 1701704242
transform 1 0 30084 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_329
timestamp 1701704242
transform 1 0 30820 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_6
timestamp 1701704242
transform 1 0 1104 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_18
timestamp 1701704242
transform 1 0 2208 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1701704242
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3220 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_33
timestamp 1701704242
transform 1 0 3588 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_50
timestamp 1701704242
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_64
timestamp 1701704242
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_75
timestamp 1701704242
transform 1 0 7452 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1701704242
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1701704242
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_97
timestamp 1701704242
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_115
timestamp 1701704242
transform 1 0 11132 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 1701704242
transform 1 0 13064 0 1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1701704242
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_153
timestamp 1701704242
transform 1 0 14628 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_170
timestamp 1701704242
transform 1 0 16192 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1701704242
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1701704242
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_197
timestamp 1701704242
transform 1 0 18676 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_203
timestamp 1701704242
transform 1 0 19228 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_225
timestamp 1701704242
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_246
timestamp 1701704242
transform 1 0 23184 0 1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1701704242
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_296
timestamp 1701704242
transform 1 0 27784 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1701704242
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_321
timestamp 1701704242
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_329
timestamp 1701704242
transform 1 0 30820 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1701704242
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1701704242
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1701704242
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1701704242
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1701704242
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1701704242
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_57
timestamp 1701704242
transform 1 0 5796 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_72
timestamp 1701704242
transform 1 0 7176 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_82
timestamp 1701704242
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_100
timestamp 1701704242
transform 1 0 9752 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1701704242
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_125
timestamp 1701704242
transform 1 0 12052 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_141
timestamp 1701704242
transform 1 0 13524 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_158
timestamp 1701704242
transform 1 0 15088 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1701704242
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_191
timestamp 1701704242
transform 1 0 18124 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_195
timestamp 1701704242
transform 1 0 18492 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_211
timestamp 1701704242
transform 1 0 19964 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1701704242
transform 1 0 21068 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_263
timestamp 1701704242
transform 1 0 24748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1701704242
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1701704242
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1701704242
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1701704242
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1701704242
transform 1 0 29716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_329
timestamp 1701704242
transform 1 0 30820 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_6
timestamp 1701704242
transform 1 0 1104 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_18
timestamp 1701704242
transform 1 0 2208 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_26
timestamp 1701704242
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1701704242
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1701704242
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1701704242
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_65
timestamp 1701704242
transform 1 0 6532 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_72
timestamp 1701704242
transform 1 0 7176 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_88
timestamp 1701704242
transform 1 0 8648 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_92
timestamp 1701704242
transform 1 0 9016 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_118
timestamp 1701704242
transform 1 0 11408 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_131
timestamp 1701704242
transform 1 0 12604 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_136
timestamp 1701704242
transform 1 0 13064 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_150
timestamp 1701704242
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_168
timestamp 1701704242
transform 1 0 16008 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1701704242
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_201
timestamp 1701704242
transform 1 0 19044 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_214
timestamp 1701704242
transform 1 0 20240 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_220
timestamp 1701704242
transform 1 0 20792 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_224
timestamp 1701704242
transform 1 0 21160 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_232
timestamp 1701704242
transform 1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_238
timestamp 1701704242
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_256
timestamp 1701704242
transform 1 0 24104 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_260
timestamp 1701704242
transform 1 0 24472 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_266
timestamp 1701704242
transform 1 0 25024 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_278
timestamp 1701704242
transform 1 0 26128 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_290
timestamp 1701704242
transform 1 0 27232 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_302
timestamp 1701704242
transform 1 0 28336 0 1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1701704242
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1701704242
transform 1 0 30084 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_329
timestamp 1701704242
transform 1 0 30820 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_12
timestamp 1701704242
transform 1 0 1656 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_24
timestamp 1701704242
transform 1 0 2760 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1701704242
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1701704242
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1701704242
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 1701704242
transform 1 0 5796 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_68
timestamp 1701704242
transform 1 0 6808 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_75
timestamp 1701704242
transform 1 0 7452 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_82
timestamp 1701704242
transform 1 0 8096 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_88
timestamp 1701704242
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_96
timestamp 1701704242
transform 1 0 9384 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_113
timestamp 1701704242
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_131
timestamp 1701704242
transform 1 0 12604 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_139
timestamp 1701704242
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_141
timestamp 1701704242
transform 1 0 13524 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_158
timestamp 1701704242
transform 1 0 15088 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1701704242
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_185
timestamp 1701704242
transform 1 0 17572 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_193
timestamp 1701704242
transform 1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_197
timestamp 1701704242
transform 1 0 18676 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_216
timestamp 1701704242
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1701704242
transform 1 0 21068 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_228
timestamp 1701704242
transform 1 0 21528 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_237
timestamp 1701704242
transform 1 0 22356 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_243
timestamp 1701704242
transform 1 0 22908 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_251
timestamp 1701704242
transform 1 0 23644 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_269
timestamp 1701704242
transform 1 0 25300 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1701704242
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1701704242
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_293
timestamp 1701704242
transform 1 0 27508 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_299
timestamp 1701704242
transform 1 0 28060 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_306
timestamp 1701704242
transform 1 0 28704 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_309
timestamp 1701704242
transform 1 0 28980 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_321
timestamp 1701704242
transform 1 0 30084 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_325
timestamp 1701704242
transform 1 0 30452 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 31096 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1701704242
transform 1 0 15548 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1701704242
transform 1 0 16192 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 17572 0 1 544
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1701704242
transform 1 0 17480 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1701704242
transform 1 0 18124 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 31372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 31372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 31372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 31372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 31372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 31372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 31372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 31372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 31372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 31372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 31372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 31372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 31372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 31372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 31372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 31372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 31372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 31372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1701704242
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 31372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1701704242
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 31372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1701704242
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 31372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1701704242
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 31372 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1701704242
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 31372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1701704242
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 31372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1701704242
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 31372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1701704242
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 31372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1701704242
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 31372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1701704242
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 31372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1701704242
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 31372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1701704242
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 31372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1701704242
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 31372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1701704242
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 29256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer2
timestamp 1701704242
transform 1 0 30636 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer3
timestamp 1701704242
transform -1 0 29348 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer4
timestamp 1701704242
transform 1 0 30268 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer5
timestamp 1701704242
transform 1 0 28520 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer6
timestamp 1701704242
transform 1 0 29348 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1701704242
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1701704242
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1701704242
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1701704242
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1701704242
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1701704242
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1701704242
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1701704242
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_82
timestamp 1701704242
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp 1701704242
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 1701704242
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 1701704242
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 1701704242
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 1701704242
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 1701704242
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp 1701704242
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 1701704242
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_97
timestamp 1701704242
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 1701704242
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 1701704242
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 1701704242
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_101
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_103
timestamp 1701704242
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_104
timestamp 1701704242
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_105
timestamp 1701704242
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_108
timestamp 1701704242
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_109
timestamp 1701704242
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_110
timestamp 1701704242
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_111
timestamp 1701704242
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_112
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_113
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_114
timestamp 1701704242
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_115
timestamp 1701704242
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1701704242
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_117
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_118
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_119
timestamp 1701704242
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1701704242
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1701704242
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1701704242
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_123
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1701704242
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1701704242
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1701704242
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1701704242
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1701704242
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_132
timestamp 1701704242
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_133
timestamp 1701704242
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp 1701704242
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp 1701704242
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp 1701704242
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_140
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_141
timestamp 1701704242
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_142
timestamp 1701704242
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_143
timestamp 1701704242
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_144
timestamp 1701704242
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_145
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_146
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_147
timestamp 1701704242
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_148
timestamp 1701704242
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_149
timestamp 1701704242
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_150
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_152
timestamp 1701704242
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_153
timestamp 1701704242
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_154
timestamp 1701704242
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_155
timestamp 1701704242
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_156
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_157
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_158
timestamp 1701704242
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_159
timestamp 1701704242
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 1701704242
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_162
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_163
timestamp 1701704242
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 1701704242
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 1701704242
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 1701704242
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_167
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_168
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 1701704242
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_170
timestamp 1701704242
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 1701704242
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_172
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 1701704242
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 1701704242
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 1701704242
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 1701704242
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 1701704242
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 1701704242
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 1701704242
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_183
timestamp 1701704242
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_184
timestamp 1701704242
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_185
timestamp 1701704242
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 1701704242
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 1701704242
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 1701704242
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 1701704242
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_190
timestamp 1701704242
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_191
timestamp 1701704242
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_192
timestamp 1701704242
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 1701704242
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_194
timestamp 1701704242
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1701704242
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 1701704242
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 1701704242
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 1701704242
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 1701704242
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_200
timestamp 1701704242
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_201
timestamp 1701704242
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 1701704242
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 1701704242
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 1701704242
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_205
timestamp 1701704242
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 1701704242
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 1701704242
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 1701704242
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_209
timestamp 1701704242
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_210
timestamp 1701704242
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 1701704242
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 1701704242
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_213
timestamp 1701704242
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_214
timestamp 1701704242
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_215
timestamp 1701704242
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 1701704242
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 1701704242
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_218
timestamp 1701704242
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_219
timestamp 1701704242
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_220
timestamp 1701704242
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_221
timestamp 1701704242
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_222
timestamp 1701704242
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_223
timestamp 1701704242
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_224
timestamp 1701704242
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_225
timestamp 1701704242
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_226
timestamp 1701704242
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_227
timestamp 1701704242
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_228
timestamp 1701704242
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_229
timestamp 1701704242
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_230
timestamp 1701704242
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_231
timestamp 1701704242
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_232
timestamp 1701704242
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_233
timestamp 1701704242
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_234
timestamp 1701704242
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_235
timestamp 1701704242
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_236
timestamp 1701704242
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_237
timestamp 1701704242
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_238
timestamp 1701704242
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_239
timestamp 1701704242
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_240
timestamp 1701704242
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_241
timestamp 1701704242
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_242
timestamp 1701704242
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_243
timestamp 1701704242
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_244
timestamp 1701704242
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_245
timestamp 1701704242
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_246
timestamp 1701704242
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_247
timestamp 1701704242
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_248
timestamp 1701704242
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_249
timestamp 1701704242
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_250
timestamp 1701704242
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_251
timestamp 1701704242
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_252
timestamp 1701704242
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_253
timestamp 1701704242
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_254
timestamp 1701704242
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_255
timestamp 1701704242
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_256
timestamp 1701704242
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_257
timestamp 1701704242
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_258
timestamp 1701704242
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_259
timestamp 1701704242
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_260
timestamp 1701704242
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_261
timestamp 1701704242
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_262
timestamp 1701704242
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_263
timestamp 1701704242
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp 1701704242
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1701704242
transform 1 0 28888 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  tdc0.g_dly_chain_even\[0\].dly_stg1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 25116 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  tdc0.g_dly_chain_even\[0\].dly_stg2
timestamp 1701704242
transform 1 0 25852 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[1\].dly_stg1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 25852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[1\].dly_stg2
timestamp 1701704242
transform -1 0 25852 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[2\].dly_stg1
timestamp 1701704242
transform -1 0 27140 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[2\].dly_stg2
timestamp 1701704242
transform -1 0 27692 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[3\].dly_stg1
timestamp 1701704242
transform 1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[3\].dly_stg2
timestamp 1701704242
transform 1 0 27968 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[4\].dly_stg1
timestamp 1701704242
transform -1 0 27968 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[4\].dly_stg2
timestamp 1701704242
transform -1 0 28244 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[5\].dly_stg1
timestamp 1701704242
transform 1 0 28796 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[5\].dly_stg2
timestamp 1701704242
transform -1 0 28520 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[6\].dly_stg1
timestamp 1701704242
transform -1 0 28796 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[6\].dly_stg2
timestamp 1701704242
transform 1 0 28980 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[7\].dly_stg1
timestamp 1701704242
transform -1 0 29532 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[7\].dly_stg2
timestamp 1701704242
transform 1 0 30820 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[8\].dly_stg1
timestamp 1701704242
transform -1 0 29900 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[8\].dly_stg2
timestamp 1701704242
transform 1 0 29348 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[9\].dly_stg1
timestamp 1701704242
transform 1 0 28796 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[9\].dly_stg2
timestamp 1701704242
transform -1 0 28796 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[10\].dly_stg1
timestamp 1701704242
transform 1 0 30452 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[10\].dly_stg2
timestamp 1701704242
transform -1 0 29256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[11\].dly_stg1
timestamp 1701704242
transform -1 0 29164 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[11\].dly_stg2
timestamp 1701704242
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[12\].dly_stg1
timestamp 1701704242
transform -1 0 29532 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[12\].dly_stg2
timestamp 1701704242
transform -1 0 29808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[13\].dly_stg1
timestamp 1701704242
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[13\].dly_stg2
timestamp 1701704242
transform 1 0 28796 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[14\].dly_stg1
timestamp 1701704242
transform 1 0 30544 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[14\].dly_stg2
timestamp 1701704242
transform -1 0 30268 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[15\].dly_stg1
timestamp 1701704242
transform 1 0 30820 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[15\].dly_stg2
timestamp 1701704242
transform -1 0 28152 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[16\].dly_stg1
timestamp 1701704242
transform 1 0 30728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[16\].dly_stg2
timestamp 1701704242
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[17\].dly_stg1
timestamp 1701704242
transform -1 0 28612 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[17\].dly_stg2
timestamp 1701704242
transform 1 0 28704 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[18\].dly_stg1
timestamp 1701704242
transform 1 0 30820 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[18\].dly_stg2
timestamp 1701704242
transform -1 0 28336 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[19\].dly_stg1
timestamp 1701704242
transform -1 0 28796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[19\].dly_stg2
timestamp 1701704242
transform -1 0 27692 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[20\].dly_stg1
timestamp 1701704242
transform 1 0 27692 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[20\].dly_stg2
timestamp 1701704242
transform -1 0 26312 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[21\].dly_stg1
timestamp 1701704242
transform -1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[21\].dly_stg2
timestamp 1701704242
transform -1 0 27140 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[22\].dly_stg1
timestamp 1701704242
transform -1 0 25300 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[22\].dly_stg2
timestamp 1701704242
transform 1 0 26312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[23\].dly_stg1
timestamp 1701704242
transform -1 0 26036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[23\].dly_stg2
timestamp 1701704242
transform -1 0 24656 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[24\].dly_stg1
timestamp 1701704242
transform 1 0 23828 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[24\].dly_stg2
timestamp 1701704242
transform 1 0 24932 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[25\].dly_stg1
timestamp 1701704242
transform -1 0 24380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[25\].dly_stg2
timestamp 1701704242
transform 1 0 24380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[26\].dly_stg1
timestamp 1701704242
transform 1 0 22816 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[26\].dly_stg2
timestamp 1701704242
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[27\].dly_stg1
timestamp 1701704242
transform -1 0 22632 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[27\].dly_stg2
timestamp 1701704242
transform -1 0 22080 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[28\].dly_stg1
timestamp 1701704242
transform -1 0 21528 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[28\].dly_stg2
timestamp 1701704242
transform 1 0 21528 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[29\].dly_stg1
timestamp 1701704242
transform -1 0 22356 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[29\].dly_stg2
timestamp 1701704242
transform -1 0 22172 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[30\].dly_stg1
timestamp 1701704242
transform 1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[30\].dly_stg2
timestamp 1701704242
transform 1 0 22448 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[31\].dly_stg1
timestamp 1701704242
transform -1 0 22080 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[31\].dly_stg2
timestamp 1701704242
transform 1 0 22264 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[32\].dly_stg1
timestamp 1701704242
transform -1 0 22264 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[32\].dly_stg2
timestamp 1701704242
transform -1 0 21712 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[33\].dly_stg1
timestamp 1701704242
transform 1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[33\].dly_stg2
timestamp 1701704242
transform 1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[34\].dly_stg1
timestamp 1701704242
transform -1 0 22264 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[34\].dly_stg2
timestamp 1701704242
transform 1 0 22724 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[35\].dly_stg1
timestamp 1701704242
transform -1 0 22632 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[35\].dly_stg2
timestamp 1701704242
transform -1 0 22908 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[36\].dly_stg1
timestamp 1701704242
transform -1 0 23736 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[36\].dly_stg2
timestamp 1701704242
transform 1 0 23460 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[37\].dly_stg1
timestamp 1701704242
transform 1 0 24380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[37\].dly_stg2
timestamp 1701704242
transform -1 0 24932 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[38\].dly_stg1
timestamp 1701704242
transform -1 0 25024 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[38\].dly_stg2
timestamp 1701704242
transform -1 0 25300 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[39\].dly_stg1
timestamp 1701704242
transform 1 0 26680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[39\].dly_stg2
timestamp 1701704242
transform 1 0 26404 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[40\].dly_stg1
timestamp 1701704242
transform 1 0 26404 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[40\].dly_stg2
timestamp 1701704242
transform 1 0 27232 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[41\].dly_stg1
timestamp 1701704242
transform -1 0 28060 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[41\].dly_stg2
timestamp 1701704242
transform -1 0 27600 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[42\].dly_stg1
timestamp 1701704242
transform -1 0 28428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[42\].dly_stg2
timestamp 1701704242
transform -1 0 28704 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[43\].dly_stg1
timestamp 1701704242
transform -1 0 29532 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[43\].dly_stg2
timestamp 1701704242
transform 1 0 28980 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[44\].dly_stg1
timestamp 1701704242
transform -1 0 29532 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[44\].dly_stg2
timestamp 1701704242
transform 1 0 29532 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[45\].dly_stg1
timestamp 1701704242
transform -1 0 28612 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[45\].dly_stg2
timestamp 1701704242
transform -1 0 29532 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[46\].dly_stg1
timestamp 1701704242
transform -1 0 29164 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[46\].dly_stg2
timestamp 1701704242
transform 1 0 29164 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[47\].dly_stg1
timestamp 1701704242
transform -1 0 28612 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[47\].dly_stg2
timestamp 1701704242
transform -1 0 28336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[48\].dly_stg1
timestamp 1701704242
transform 1 0 27508 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[48\].dly_stg2
timestamp 1701704242
transform -1 0 28152 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[49\].dly_stg1
timestamp 1701704242
transform 1 0 26772 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[49\].dly_stg2
timestamp 1701704242
transform -1 0 27324 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[50\].dly_stg1
timestamp 1701704242
transform -1 0 26128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[50\].dly_stg2
timestamp 1701704242
transform 1 0 26036 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[51\].dly_stg1
timestamp 1701704242
transform -1 0 25208 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[51\].dly_stg2
timestamp 1701704242
transform 1 0 25760 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[52\].dly_stg1
timestamp 1701704242
transform -1 0 25668 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[52\].dly_stg2
timestamp 1701704242
transform -1 0 25944 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[53\].dly_stg1
timestamp 1701704242
transform -1 0 24748 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[53\].dly_stg2
timestamp 1701704242
transform -1 0 24472 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[54\].dly_stg1
timestamp 1701704242
transform -1 0 22908 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[54\].dly_stg2
timestamp 1701704242
transform 1 0 23460 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[55\].dly_stg1
timestamp 1701704242
transform -1 0 22448 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[55\].dly_stg2
timestamp 1701704242
transform -1 0 22356 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[56\].dly_stg1
timestamp 1701704242
transform 1 0 20792 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[56\].dly_stg2
timestamp 1701704242
transform 1 0 21252 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[57\].dly_stg1
timestamp 1701704242
transform -1 0 19964 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[57\].dly_stg2
timestamp 1701704242
transform -1 0 19688 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[58\].dly_stg1
timestamp 1701704242
transform -1 0 16836 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[58\].dly_stg2
timestamp 1701704242
transform -1 0 16376 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[59\].dly_stg1
timestamp 1701704242
transform -1 0 19136 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[59\].dly_stg2
timestamp 1701704242
transform 1 0 19688 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[60\].dly_stg1
timestamp 1701704242
transform 1 0 19320 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[60\].dly_stg2
timestamp 1701704242
transform -1 0 20148 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[61\].dly_stg1
timestamp 1701704242
transform 1 0 20148 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[61\].dly_stg2
timestamp 1701704242
transform 1 0 20700 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[62\].dly_stg1
timestamp 1701704242
transform -1 0 21252 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[62\].dly_stg2
timestamp 1701704242
transform -1 0 19964 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[63\].dly_stg1
timestamp 1701704242
transform -1 0 22356 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[63\].dly_stg2
timestamp 1701704242
transform -1 0 22080 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[64\].dly_stg1
timestamp 1701704242
transform -1 0 20516 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[64\].dly_stg2
timestamp 1701704242
transform 1 0 20700 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[65\].dly_stg1
timestamp 1701704242
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[65\].dly_stg2
timestamp 1701704242
transform -1 0 20792 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[66\].dly_stg1
timestamp 1701704242
transform -1 0 19780 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[66\].dly_stg2
timestamp 1701704242
transform -1 0 18400 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[67\].dly_stg1
timestamp 1701704242
transform -1 0 19228 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[67\].dly_stg2
timestamp 1701704242
transform -1 0 18676 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[68\].dly_stg1
timestamp 1701704242
transform -1 0 17480 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[68\].dly_stg2
timestamp 1701704242
transform -1 0 17204 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[69\].dly_stg1
timestamp 1701704242
transform -1 0 15180 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[69\].dly_stg2
timestamp 1701704242
transform 1 0 15732 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[70\].dly_stg1
timestamp 1701704242
transform -1 0 15364 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[70\].dly_stg2
timestamp 1701704242
transform -1 0 14904 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[71\].dly_stg1
timestamp 1701704242
transform -1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[71\].dly_stg2
timestamp 1701704242
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[72\].dly_stg1
timestamp 1701704242
transform 1 0 13156 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[72\].dly_stg2
timestamp 1701704242
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[73\].dly_stg1
timestamp 1701704242
transform -1 0 12696 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[73\].dly_stg2
timestamp 1701704242
transform -1 0 11684 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[74\].dly_stg1
timestamp 1701704242
transform 1 0 12144 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[74\].dly_stg2
timestamp 1701704242
transform 1 0 11868 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[75\].dly_stg1
timestamp 1701704242
transform 1 0 12512 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[75\].dly_stg2
timestamp 1701704242
transform -1 0 12236 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[76\].dly_stg1
timestamp 1701704242
transform -1 0 10856 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[76\].dly_stg2
timestamp 1701704242
transform -1 0 11316 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[77\].dly_stg1
timestamp 1701704242
transform -1 0 10304 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[77\].dly_stg2
timestamp 1701704242
transform -1 0 10396 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[78\].dly_stg1
timestamp 1701704242
transform -1 0 9752 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[78\].dly_stg2
timestamp 1701704242
transform -1 0 9476 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[79\].dly_stg1
timestamp 1701704242
transform 1 0 9292 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[79\].dly_stg2
timestamp 1701704242
transform -1 0 9292 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[80\].dly_stg1
timestamp 1701704242
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[80\].dly_stg2
timestamp 1701704242
transform 1 0 10120 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[81\].dly_stg1
timestamp 1701704242
transform -1 0 9752 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[81\].dly_stg2
timestamp 1701704242
transform -1 0 10028 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[82\].dly_stg1
timestamp 1701704242
transform -1 0 10120 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[82\].dly_stg2
timestamp 1701704242
transform -1 0 10396 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[83\].dly_stg1
timestamp 1701704242
transform -1 0 9752 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[83\].dly_stg2
timestamp 1701704242
transform 1 0 9752 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[84\].dly_stg1
timestamp 1701704242
transform -1 0 10488 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[84\].dly_stg2
timestamp 1701704242
transform -1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[85\].dly_stg1
timestamp 1701704242
transform -1 0 9384 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[85\].dly_stg2
timestamp 1701704242
transform 1 0 10120 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[86\].dly_stg1
timestamp 1701704242
transform -1 0 10948 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[86\].dly_stg2
timestamp 1701704242
transform -1 0 10396 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[87\].dly_stg1
timestamp 1701704242
transform -1 0 11592 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[87\].dly_stg2
timestamp 1701704242
transform -1 0 11316 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[88\].dly_stg1
timestamp 1701704242
transform 1 0 12328 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[88\].dly_stg2
timestamp 1701704242
transform 1 0 12512 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[89\].dly_stg1
timestamp 1701704242
transform -1 0 11960 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[89\].dly_stg2
timestamp 1701704242
transform 1 0 12788 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[90\].dly_stg1
timestamp 1701704242
transform -1 0 13248 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[90\].dly_stg2
timestamp 1701704242
transform -1 0 12696 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[91\].dly_stg1
timestamp 1701704242
transform -1 0 13800 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[91\].dly_stg2
timestamp 1701704242
transform 1 0 14076 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[92\].dly_stg1
timestamp 1701704242
transform -1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[92\].dly_stg2
timestamp 1701704242
transform 1 0 12328 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[93\].dly_stg1
timestamp 1701704242
transform -1 0 10304 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[93\].dly_stg2
timestamp 1701704242
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[94\].dly_stg1
timestamp 1701704242
transform -1 0 10028 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[94\].dly_stg2
timestamp 1701704242
transform -1 0 9752 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[95\].dly_stg1
timestamp 1701704242
transform -1 0 8648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[95\].dly_stg2
timestamp 1701704242
transform -1 0 8280 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[96\].dly_stg1
timestamp 1701704242
transform 1 0 7452 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[96\].dly_stg2
timestamp 1701704242
transform -1 0 7820 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[97\].dly_stg1
timestamp 1701704242
transform -1 0 6900 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[97\].dly_stg2
timestamp 1701704242
transform -1 0 7176 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[98\].dly_stg1
timestamp 1701704242
transform -1 0 7452 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[98\].dly_stg2
timestamp 1701704242
transform -1 0 6900 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[99\].dly_stg1
timestamp 1701704242
transform -1 0 6164 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[99\].dly_stg2
timestamp 1701704242
transform -1 0 5888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[100\].dly_stg1
timestamp 1701704242
transform -1 0 5704 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[100\].dly_stg2
timestamp 1701704242
transform -1 0 5428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[101\].dly_stg1
timestamp 1701704242
transform 1 0 3772 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[101\].dly_stg2
timestamp 1701704242
transform -1 0 4600 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[102\].dly_stg1
timestamp 1701704242
transform 1 0 3220 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[102\].dly_stg2
timestamp 1701704242
transform 1 0 3588 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[103\].dly_stg1
timestamp 1701704242
transform 1 0 2024 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[103\].dly_stg2
timestamp 1701704242
transform -1 0 2576 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[104\].dly_stg1
timestamp 1701704242
transform -1 0 2116 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[104\].dly_stg2
timestamp 1701704242
transform -1 0 1748 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[105\].dly_stg1
timestamp 1701704242
transform -1 0 1656 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[105\].dly_stg2
timestamp 1701704242
transform 1 0 2208 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[106\].dly_stg1
timestamp 1701704242
transform -1 0 2116 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[106\].dly_stg2
timestamp 1701704242
transform -1 0 1840 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[107\].dly_stg1
timestamp 1701704242
transform -1 0 2300 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[107\].dly_stg2
timestamp 1701704242
transform -1 0 2024 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[108\].dly_stg1
timestamp 1701704242
transform 1 0 1012 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[108\].dly_stg2
timestamp 1701704242
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[109\].dly_stg1
timestamp 1701704242
transform 1 0 1932 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[109\].dly_stg2
timestamp 1701704242
transform 1 0 1288 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[110\].dly_stg1
timestamp 1701704242
transform -1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[110\].dly_stg2
timestamp 1701704242
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[111\].dly_stg1
timestamp 1701704242
transform 1 0 1748 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[111\].dly_stg2
timestamp 1701704242
transform -1 0 1748 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[112\].dly_stg1
timestamp 1701704242
transform -1 0 1748 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[112\].dly_stg2
timestamp 1701704242
transform 1 0 1748 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[113\].dly_stg1
timestamp 1701704242
transform 1 0 2300 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[113\].dly_stg2
timestamp 1701704242
transform -1 0 1472 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[114\].dly_stg1
timestamp 1701704242
transform 1 0 1564 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[114\].dly_stg2
timestamp 1701704242
transform -1 0 1196 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[115\].dly_stg1
timestamp 1701704242
transform 1 0 2116 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[115\].dly_stg2
timestamp 1701704242
transform -1 0 2576 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[116\].dly_stg1
timestamp 1701704242
transform 1 0 2852 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[116\].dly_stg2
timestamp 1701704242
transform -1 0 3956 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[117\].dly_stg1
timestamp 1701704242
transform -1 0 3588 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[117\].dly_stg2
timestamp 1701704242
transform 1 0 4232 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[118\].dly_stg1
timestamp 1701704242
transform -1 0 3956 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[118\].dly_stg2
timestamp 1701704242
transform -1 0 3864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[119\].dly_stg1
timestamp 1701704242
transform 1 0 4416 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[119\].dly_stg2
timestamp 1701704242
transform -1 0 4324 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[120\].dly_stg1
timestamp 1701704242
transform -1 0 4324 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[120\].dly_stg2
timestamp 1701704242
transform 1 0 4600 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[121\].dly_stg1
timestamp 1701704242
transform -1 0 4508 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[121\].dly_stg2
timestamp 1701704242
transform -1 0 4232 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[122\].dly_stg1
timestamp 1701704242
transform -1 0 4232 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[122\].dly_stg2
timestamp 1701704242
transform 1 0 4508 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[123\].dly_stg1
timestamp 1701704242
transform 1 0 4784 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[123\].dly_stg2
timestamp 1701704242
transform -1 0 5152 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[124\].dly_stg1
timestamp 1701704242
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[124\].dly_stg2
timestamp 1701704242
transform 1 0 5612 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[125\].dly_stg1
timestamp 1701704242
transform -1 0 6900 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[125\].dly_stg2
timestamp 1701704242
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[126\].dly_stg1
timestamp 1701704242
transform -1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[126\].dly_stg2
timestamp 1701704242
transform -1 0 7544 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[127\].dly_stg1
timestamp 1701704242
transform -1 0 8188 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[127\].dly_stg2
timestamp 1701704242
transform 1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[128\].dly_stg1
timestamp 1701704242
transform 1 0 7176 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[128\].dly_stg2
timestamp 1701704242
transform -1 0 7728 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[129\].dly_stg1
timestamp 1701704242
transform 1 0 6900 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[129\].dly_stg2
timestamp 1701704242
transform 1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[130\].dly_stg1
timestamp 1701704242
transform -1 0 7452 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[130\].dly_stg2
timestamp 1701704242
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[131\].dly_stg1
timestamp 1701704242
transform 1 0 6992 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[131\].dly_stg2
timestamp 1701704242
transform 1 0 7544 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[132\].dly_stg1
timestamp 1701704242
transform -1 0 6348 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[132\].dly_stg2
timestamp 1701704242
transform -1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[133\].dly_stg1
timestamp 1701704242
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[133\].dly_stg2
timestamp 1701704242
transform -1 0 5704 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[134\].dly_stg1
timestamp 1701704242
transform -1 0 6348 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[134\].dly_stg2
timestamp 1701704242
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[135\].dly_stg1
timestamp 1701704242
transform -1 0 6348 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[135\].dly_stg2
timestamp 1701704242
transform -1 0 7636 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[136\].dly_stg1
timestamp 1701704242
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[136\].dly_stg2
timestamp 1701704242
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[137\].dly_stg1
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[137\].dly_stg2
timestamp 1701704242
transform 1 0 9200 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[138\].dly_stg1
timestamp 1701704242
transform -1 0 10028 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[138\].dly_stg2
timestamp 1701704242
transform -1 0 9752 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[139\].dly_stg1
timestamp 1701704242
transform 1 0 10672 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[139\].dly_stg2
timestamp 1701704242
transform 1 0 10396 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[140\].dly_stg1
timestamp 1701704242
transform -1 0 9844 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[140\].dly_stg2
timestamp 1701704242
transform 1 0 10120 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[141\].dly_stg1
timestamp 1701704242
transform -1 0 9016 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[141\].dly_stg2
timestamp 1701704242
transform -1 0 8740 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[142\].dly_stg1
timestamp 1701704242
transform -1 0 7728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[142\].dly_stg2
timestamp 1701704242
transform -1 0 8004 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[143\].dly_stg1
timestamp 1701704242
transform -1 0 7544 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[143\].dly_stg2
timestamp 1701704242
transform -1 0 6900 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[144\].dly_stg1
timestamp 1701704242
transform 1 0 5520 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[144\].dly_stg2
timestamp 1701704242
transform -1 0 6348 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[145\].dly_stg1
timestamp 1701704242
transform -1 0 4968 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[145\].dly_stg2
timestamp 1701704242
transform -1 0 5244 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[146\].dly_stg1
timestamp 1701704242
transform -1 0 4416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[146\].dly_stg2
timestamp 1701704242
transform -1 0 4416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[147\].dly_stg1
timestamp 1701704242
transform -1 0 3772 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[147\].dly_stg2
timestamp 1701704242
transform -1 0 3864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[148\].dly_stg1
timestamp 1701704242
transform 1 0 2392 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[148\].dly_stg2
timestamp 1701704242
transform -1 0 2668 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[149\].dly_stg1
timestamp 1701704242
transform -1 0 2944 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[149\].dly_stg2
timestamp 1701704242
transform -1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[150\].dly_stg1
timestamp 1701704242
transform -1 0 1932 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[150\].dly_stg2
timestamp 1701704242
transform -1 0 1564 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[151\].dly_stg1
timestamp 1701704242
transform -1 0 1932 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[151\].dly_stg2
timestamp 1701704242
transform 1 0 1932 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[152\].dly_stg1
timestamp 1701704242
transform -1 0 2760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[152\].dly_stg2
timestamp 1701704242
transform -1 0 1656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[153\].dly_stg1
timestamp 1701704242
transform 1 0 1288 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[153\].dly_stg2
timestamp 1701704242
transform 1 0 2392 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[154\].dly_stg1
timestamp 1701704242
transform -1 0 1932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[154\].dly_stg2
timestamp 1701704242
transform 1 0 2852 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[155\].dly_stg1
timestamp 1701704242
transform -1 0 2852 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[155\].dly_stg2
timestamp 1701704242
transform -1 0 2576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[156\].dly_stg1
timestamp 1701704242
transform -1 0 3128 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[156\].dly_stg2
timestamp 1701704242
transform 1 0 3128 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[157\].dly_stg1
timestamp 1701704242
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[157\].dly_stg2
timestamp 1701704242
transform -1 0 4508 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[158\].dly_stg1
timestamp 1701704242
transform 1 0 4600 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[158\].dly_stg2
timestamp 1701704242
transform -1 0 5152 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[159\].dly_stg1
timestamp 1701704242
transform -1 0 5980 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[159\].dly_stg2
timestamp 1701704242
transform -1 0 6256 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[160\].dly_stg1
timestamp 1701704242
transform 1 0 6532 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[160\].dly_stg2
timestamp 1701704242
transform -1 0 7360 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[161\].dly_stg1
timestamp 1701704242
transform -1 0 7544 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[161\].dly_stg2
timestamp 1701704242
transform 1 0 8004 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[162\].dly_stg1
timestamp 1701704242
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[162\].dly_stg2
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[163\].dly_stg1
timestamp 1701704242
transform -1 0 8648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[163\].dly_stg2
timestamp 1701704242
transform 1 0 8096 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[164\].dly_stg1
timestamp 1701704242
transform -1 0 9568 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[164\].dly_stg2
timestamp 1701704242
transform -1 0 9200 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[165\].dly_stg1
timestamp 1701704242
transform -1 0 10028 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[165\].dly_stg2
timestamp 1701704242
transform -1 0 9752 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[166\].dly_stg1
timestamp 1701704242
transform -1 0 10856 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[166\].dly_stg2
timestamp 1701704242
transform -1 0 10304 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[167\].dly_stg1
timestamp 1701704242
transform -1 0 12512 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[167\].dly_stg2
timestamp 1701704242
transform -1 0 12420 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[168\].dly_stg1
timestamp 1701704242
transform -1 0 13248 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[168\].dly_stg2
timestamp 1701704242
transform 1 0 12696 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[169\].dly_stg1
timestamp 1701704242
transform 1 0 13524 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[169\].dly_stg2
timestamp 1701704242
transform -1 0 14076 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[170\].dly_stg1
timestamp 1701704242
transform -1 0 14628 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[170\].dly_stg2
timestamp 1701704242
transform -1 0 14352 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[171\].dly_stg1
timestamp 1701704242
transform -1 0 15640 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[171\].dly_stg2
timestamp 1701704242
transform -1 0 15364 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[172\].dly_stg1
timestamp 1701704242
transform 1 0 15456 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[172\].dly_stg2
timestamp 1701704242
transform 1 0 15732 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[173\].dly_stg1
timestamp 1701704242
transform -1 0 17020 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[173\].dly_stg2
timestamp 1701704242
transform 1 0 17020 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[174\].dly_stg1
timestamp 1701704242
transform -1 0 18124 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[174\].dly_stg2
timestamp 1701704242
transform -1 0 17204 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[175\].dly_stg1
timestamp 1701704242
transform 1 0 18216 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[175\].dly_stg2
timestamp 1701704242
transform -1 0 19228 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[176\].dly_stg1
timestamp 1701704242
transform 1 0 19780 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[176\].dly_stg2
timestamp 1701704242
transform -1 0 20332 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[177\].dly_stg1
timestamp 1701704242
transform 1 0 19964 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[177\].dly_stg2
timestamp 1701704242
transform 1 0 20148 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[178\].dly_stg1
timestamp 1701704242
transform -1 0 21528 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[178\].dly_stg2
timestamp 1701704242
transform -1 0 20884 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[179\].dly_stg1
timestamp 1701704242
transform 1 0 21804 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[179\].dly_stg2
timestamp 1701704242
transform -1 0 21804 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[180\].dly_stg1
timestamp 1701704242
transform 1 0 21804 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[180\].dly_stg2
timestamp 1701704242
transform -1 0 22080 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[181\].dly_stg1
timestamp 1701704242
transform -1 0 24104 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[181\].dly_stg2
timestamp 1701704242
transform -1 0 23644 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[182\].dly_stg1
timestamp 1701704242
transform 1 0 23460 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[182\].dly_stg2
timestamp 1701704242
transform 1 0 24656 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[183\].dly_stg1
timestamp 1701704242
transform -1 0 24380 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[183\].dly_stg2
timestamp 1701704242
transform 1 0 24196 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[184\].dly_stg1
timestamp 1701704242
transform 1 0 25484 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[184\].dly_stg2
timestamp 1701704242
transform 1 0 26036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[185\].dly_stg1
timestamp 1701704242
transform -1 0 26128 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[185\].dly_stg2
timestamp 1701704242
transform -1 0 25484 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[186\].dly_stg1
timestamp 1701704242
transform 1 0 26772 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[186\].dly_stg2
timestamp 1701704242
transform -1 0 26772 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[187\].dly_stg1
timestamp 1701704242
transform 1 0 27048 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[187\].dly_stg2
timestamp 1701704242
transform 1 0 27416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[188\].dly_stg1
timestamp 1701704242
transform -1 0 27416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[188\].dly_stg2
timestamp 1701704242
transform 1 0 27692 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[189\].dly_stg1
timestamp 1701704242
transform 1 0 28336 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[189\].dly_stg2
timestamp 1701704242
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[190\].dly_stg1
timestamp 1701704242
transform -1 0 29256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[190\].dly_stg2
timestamp 1701704242
transform 1 0 29808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[191\].dly_stg1
timestamp 1701704242
transform 1 0 29256 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[191\].dly_stg2
timestamp 1701704242
transform 1 0 30084 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[192\].dly_stg1
timestamp 1701704242
transform 1 0 30636 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[192\].dly_stg2
timestamp 1701704242
transform 1 0 29808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[0\].dly_stg1
timestamp 1701704242
transform -1 0 25208 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[0\].dly_stg2
timestamp 1701704242
transform 1 0 25484 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[1\].dly_stg1
timestamp 1701704242
transform 1 0 26588 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[1\].dly_stg2
timestamp 1701704242
transform 1 0 26312 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[2\].dly_stg1
timestamp 1701704242
transform 1 0 27140 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[2\].dly_stg2
timestamp 1701704242
transform 1 0 27692 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[3\].dly_stg1
timestamp 1701704242
transform 1 0 27416 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[3\].dly_stg2
timestamp 1701704242
transform 1 0 27140 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[4\].dly_stg1
timestamp 1701704242
transform 1 0 28520 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[4\].dly_stg2
timestamp 1701704242
transform 1 0 28244 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[5\].dly_stg1
timestamp 1701704242
transform 1 0 28244 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[5\].dly_stg2
timestamp 1701704242
transform 1 0 29072 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[6\].dly_stg1
timestamp 1701704242
transform 1 0 28980 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[6\].dly_stg2
timestamp 1701704242
transform 1 0 29900 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[7\].dly_stg1
timestamp 1701704242
transform 1 0 29072 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[7\].dly_stg2
timestamp 1701704242
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[8\].dly_stg1
timestamp 1701704242
transform -1 0 30176 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[8\].dly_stg2
timestamp 1701704242
transform -1 0 29348 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[9\].dly_stg1
timestamp 1701704242
transform -1 0 29532 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[9\].dly_stg2
timestamp 1701704242
transform -1 0 29808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[10\].dly_stg1
timestamp 1701704242
transform -1 0 29440 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[10\].dly_stg2
timestamp 1701704242
transform -1 0 30452 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[11\].dly_stg1
timestamp 1701704242
transform 1 0 28336 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[11\].dly_stg2
timestamp 1701704242
transform -1 0 29256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[12\].dly_stg1
timestamp 1701704242
transform -1 0 30084 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[12\].dly_stg2
timestamp 1701704242
transform 1 0 30084 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[13\].dly_stg1
timestamp 1701704242
transform 1 0 29716 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[13\].dly_stg2
timestamp 1701704242
transform 1 0 29072 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[14\].dly_stg1
timestamp 1701704242
transform 1 0 30636 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[14\].dly_stg2
timestamp 1701704242
transform -1 0 29256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[15\].dly_stg1
timestamp 1701704242
transform -1 0 30636 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[15\].dly_stg2
timestamp 1701704242
transform -1 0 28796 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[16\].dly_stg1
timestamp 1701704242
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[16\].dly_stg2
timestamp 1701704242
transform -1 0 30728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[17\].dly_stg1
timestamp 1701704242
transform 1 0 28428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[17\].dly_stg2
timestamp 1701704242
transform 1 0 28980 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[18\].dly_stg1
timestamp 1701704242
transform -1 0 29256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[18\].dly_stg2
timestamp 1701704242
transform -1 0 27968 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[19\].dly_stg1
timestamp 1701704242
transform -1 0 28244 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[19\].dly_stg2
timestamp 1701704242
transform -1 0 28520 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[20\].dly_stg1
timestamp 1701704242
transform -1 0 27692 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[20\].dly_stg2
timestamp 1701704242
transform -1 0 26680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[21\].dly_stg1
timestamp 1701704242
transform -1 0 25576 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[21\].dly_stg2
timestamp 1701704242
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[22\].dly_stg1
timestamp 1701704242
transform -1 0 26312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[22\].dly_stg2
timestamp 1701704242
transform -1 0 24932 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[23\].dly_stg1
timestamp 1701704242
transform -1 0 25760 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[23\].dly_stg2
timestamp 1701704242
transform -1 0 25484 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[24\].dly_stg1
timestamp 1701704242
transform -1 0 23644 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[24\].dly_stg2
timestamp 1701704242
transform -1 0 24932 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[25\].dly_stg1
timestamp 1701704242
transform -1 0 23368 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[25\].dly_stg2
timestamp 1701704242
transform -1 0 24104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[26\].dly_stg1
timestamp 1701704242
transform 1 0 21988 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[26\].dly_stg2
timestamp 1701704242
transform -1 0 22356 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[27\].dly_stg1
timestamp 1701704242
transform -1 0 21252 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[27\].dly_stg2
timestamp 1701704242
transform -1 0 22540 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[28\].dly_stg1
timestamp 1701704242
transform 1 0 22356 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[28\].dly_stg2
timestamp 1701704242
transform 1 0 21528 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[29\].dly_stg1
timestamp 1701704242
transform -1 0 22080 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[29\].dly_stg2
timestamp 1701704242
transform -1 0 22448 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[30\].dly_stg1
timestamp 1701704242
transform 1 0 22080 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[30\].dly_stg2
timestamp 1701704242
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[31\].dly_stg1
timestamp 1701704242
transform 1 0 22540 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[31\].dly_stg2
timestamp 1701704242
transform -1 0 21988 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[32\].dly_stg1
timestamp 1701704242
transform 1 0 22264 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[32\].dly_stg2
timestamp 1701704242
transform 1 0 22540 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[33\].dly_stg1
timestamp 1701704242
transform 1 0 21344 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[33\].dly_stg2
timestamp 1701704242
transform 1 0 21712 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[34\].dly_stg1
timestamp 1701704242
transform 1 0 22080 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[34\].dly_stg2
timestamp 1701704242
transform 1 0 22816 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[35\].dly_stg1
timestamp 1701704242
transform 1 0 22908 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[35\].dly_stg2
timestamp 1701704242
transform 1 0 23184 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[36\].dly_stg1
timestamp 1701704242
transform 1 0 24012 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[36\].dly_stg2
timestamp 1701704242
transform -1 0 22724 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[37\].dly_stg1
timestamp 1701704242
transform 1 0 24472 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[37\].dly_stg2
timestamp 1701704242
transform 1 0 24932 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[38\].dly_stg1
timestamp 1701704242
transform 1 0 26036 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[38\].dly_stg2
timestamp 1701704242
transform 1 0 26404 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[39\].dly_stg1
timestamp 1701704242
transform 1 0 26680 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[39\].dly_stg2
timestamp 1701704242
transform 1 0 26956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[40\].dly_stg1
timestamp 1701704242
transform 1 0 27508 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[40\].dly_stg2
timestamp 1701704242
transform -1 0 26956 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[41\].dly_stg1
timestamp 1701704242
transform 1 0 27600 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[41\].dly_stg2
timestamp 1701704242
transform 1 0 27876 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[42\].dly_stg1
timestamp 1701704242
transform 1 0 28704 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[42\].dly_stg2
timestamp 1701704242
transform 1 0 28980 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[43\].dly_stg1
timestamp 1701704242
transform -1 0 29532 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[43\].dly_stg2
timestamp 1701704242
transform -1 0 29256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[44\].dly_stg1
timestamp 1701704242
transform 1 0 29808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[44\].dly_stg2
timestamp 1701704242
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[45\].dly_stg1
timestamp 1701704242
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[45\].dly_stg2
timestamp 1701704242
transform -1 0 29256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[46\].dly_stg1
timestamp 1701704242
transform -1 0 28612 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[46\].dly_stg2
timestamp 1701704242
transform -1 0 28336 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[47\].dly_stg1
timestamp 1701704242
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[47\].dly_stg2
timestamp 1701704242
transform -1 0 28060 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[48\].dly_stg1
timestamp 1701704242
transform -1 0 27048 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[48\].dly_stg2
timestamp 1701704242
transform -1 0 27876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[49\].dly_stg1
timestamp 1701704242
transform -1 0 25852 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[49\].dly_stg2
timestamp 1701704242
transform 1 0 27324 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[50\].dly_stg1
timestamp 1701704242
transform -1 0 25484 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[50\].dly_stg2
timestamp 1701704242
transform -1 0 25760 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[51\].dly_stg1
timestamp 1701704242
transform -1 0 26220 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[51\].dly_stg2
timestamp 1701704242
transform -1 0 25392 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[52\].dly_stg1
timestamp 1701704242
transform -1 0 24472 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[52\].dly_stg2
timestamp 1701704242
transform -1 0 25024 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[53\].dly_stg1
timestamp 1701704242
transform -1 0 22908 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[53\].dly_stg2
timestamp 1701704242
transform -1 0 24104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[54\].dly_stg1
timestamp 1701704242
transform -1 0 23460 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[54\].dly_stg2
timestamp 1701704242
transform -1 0 23184 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[55\].dly_stg1
timestamp 1701704242
transform -1 0 21160 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[55\].dly_stg2
timestamp 1701704242
transform -1 0 22080 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[56\].dly_stg1
timestamp 1701704242
transform -1 0 20240 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[56\].dly_stg2
timestamp 1701704242
transform -1 0 20792 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[57\].dly_stg1
timestamp 1701704242
transform -1 0 17112 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[57\].dly_stg2
timestamp 1701704242
transform -1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[58\].dly_stg1
timestamp 1701704242
transform 1 0 18584 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[58\].dly_stg2
timestamp 1701704242
transform 1 0 17848 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[59\].dly_stg1
timestamp 1701704242
transform 1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[59\].dly_stg2
timestamp 1701704242
transform -1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[60\].dly_stg1
timestamp 1701704242
transform 1 0 19596 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[60\].dly_stg2
timestamp 1701704242
transform 1 0 20424 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[61\].dly_stg1
timestamp 1701704242
transform -1 0 20240 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[61\].dly_stg2
timestamp 1701704242
transform -1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[62\].dly_stg1
timestamp 1701704242
transform 1 0 21436 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[62\].dly_stg2
timestamp 1701704242
transform 1 0 21252 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[63\].dly_stg1
timestamp 1701704242
transform 1 0 19964 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[63\].dly_stg2
timestamp 1701704242
transform -1 0 21804 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[64\].dly_stg1
timestamp 1701704242
transform -1 0 21344 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[64\].dly_stg2
timestamp 1701704242
transform 1 0 20792 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[65\].dly_stg1
timestamp 1701704242
transform -1 0 19504 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[65\].dly_stg2
timestamp 1701704242
transform -1 0 21068 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[66\].dly_stg1
timestamp 1701704242
transform -1 0 19228 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[66\].dly_stg2
timestamp 1701704242
transform -1 0 18952 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[67\].dly_stg1
timestamp 1701704242
transform -1 0 17756 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[67\].dly_stg2
timestamp 1701704242
transform -1 0 18952 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[68\].dly_stg1
timestamp 1701704242
transform -1 0 15640 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[68\].dly_stg2
timestamp 1701704242
transform -1 0 16928 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[69\].dly_stg1
timestamp 1701704242
transform -1 0 15732 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[69\].dly_stg2
timestamp 1701704242
transform -1 0 15456 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[70\].dly_stg1
timestamp 1701704242
transform -1 0 14628 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[70\].dly_stg2
timestamp 1701704242
transform -1 0 14352 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[71\].dly_stg1
timestamp 1701704242
transform -1 0 13156 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[71\].dly_stg2
timestamp 1701704242
transform 1 0 14720 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[72\].dly_stg1
timestamp 1701704242
transform -1 0 13708 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[72\].dly_stg2
timestamp 1701704242
transform -1 0 13432 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[73\].dly_stg1
timestamp 1701704242
transform -1 0 12512 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[73\].dly_stg2
timestamp 1701704242
transform -1 0 11684 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[74\].dly_stg1
timestamp 1701704242
transform -1 0 12512 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[74\].dly_stg2
timestamp 1701704242
transform -1 0 11960 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[75\].dly_stg1
timestamp 1701704242
transform -1 0 11592 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[75\].dly_stg2
timestamp 1701704242
transform -1 0 11960 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[76\].dly_stg1
timestamp 1701704242
transform -1 0 10856 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[76\].dly_stg2
timestamp 1701704242
transform -1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[77\].dly_stg1
timestamp 1701704242
transform -1 0 10028 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[77\].dly_stg2
timestamp 1701704242
transform -1 0 10028 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[78\].dly_stg1
timestamp 1701704242
transform -1 0 9844 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[78\].dly_stg2
timestamp 1701704242
transform -1 0 9660 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[79\].dly_stg1
timestamp 1701704242
transform 1 0 9844 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[79\].dly_stg2
timestamp 1701704242
transform 1 0 9568 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[80\].dly_stg1
timestamp 1701704242
transform 1 0 9200 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[80\].dly_stg2
timestamp 1701704242
transform -1 0 9752 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[81\].dly_stg1
timestamp 1701704242
transform 1 0 9568 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[81\].dly_stg2
timestamp 1701704242
transform 1 0 10028 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[82\].dly_stg1
timestamp 1701704242
transform -1 0 9568 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[82\].dly_stg2
timestamp 1701704242
transform 1 0 10396 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[83\].dly_stg1
timestamp 1701704242
transform -1 0 9476 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[83\].dly_stg2
timestamp 1701704242
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[84\].dly_stg1
timestamp 1701704242
transform -1 0 10212 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[84\].dly_stg2
timestamp 1701704242
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[85\].dly_stg1
timestamp 1701704242
transform -1 0 10672 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[85\].dly_stg2
timestamp 1701704242
transform 1 0 9844 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[86\].dly_stg1
timestamp 1701704242
transform -1 0 11592 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[86\].dly_stg2
timestamp 1701704242
transform 1 0 10948 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[87\].dly_stg1
timestamp 1701704242
transform 1 0 12052 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[87\].dly_stg2
timestamp 1701704242
transform 1 0 11684 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[88\].dly_stg1
timestamp 1701704242
transform -1 0 12236 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[88\].dly_stg2
timestamp 1701704242
transform 1 0 12236 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[89\].dly_stg1
timestamp 1701704242
transform -1 0 12972 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[89\].dly_stg2
timestamp 1701704242
transform -1 0 12420 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[90\].dly_stg1
timestamp 1701704242
transform 1 0 13248 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[90\].dly_stg2
timestamp 1701704242
transform -1 0 13064 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[91\].dly_stg1
timestamp 1701704242
transform -1 0 12328 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[91\].dly_stg2
timestamp 1701704242
transform 1 0 13800 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[92\].dly_stg1
timestamp 1701704242
transform -1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[92\].dly_stg2
timestamp 1701704242
transform -1 0 11776 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[93\].dly_stg1
timestamp 1701704242
transform -1 0 9660 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[93\].dly_stg2
timestamp 1701704242
transform -1 0 9936 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[94\].dly_stg1
timestamp 1701704242
transform -1 0 9016 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[94\].dly_stg2
timestamp 1701704242
transform -1 0 9384 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[95\].dly_stg1
timestamp 1701704242
transform -1 0 8004 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[95\].dly_stg2
timestamp 1701704242
transform -1 0 8648 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[96\].dly_stg1
timestamp 1701704242
transform -1 0 7544 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[96\].dly_stg2
timestamp 1701704242
transform 1 0 7820 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[97\].dly_stg1
timestamp 1701704242
transform -1 0 7176 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[97\].dly_stg2
timestamp 1701704242
transform -1 0 6624 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[98\].dly_stg1
timestamp 1701704242
transform -1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[98\].dly_stg2
timestamp 1701704242
transform -1 0 7176 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[99\].dly_stg1
timestamp 1701704242
transform -1 0 6348 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[99\].dly_stg2
timestamp 1701704242
transform -1 0 5612 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[100\].dly_stg1
timestamp 1701704242
transform -1 0 4968 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[100\].dly_stg2
timestamp 1701704242
transform -1 0 6072 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[101\].dly_stg1
timestamp 1701704242
transform -1 0 3772 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[101\].dly_stg2
timestamp 1701704242
transform -1 0 4324 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[102\].dly_stg1
timestamp 1701704242
transform -1 0 3128 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[102\].dly_stg2
timestamp 1701704242
transform -1 0 3588 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[103\].dly_stg1
timestamp 1701704242
transform -1 0 2024 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[103\].dly_stg2
timestamp 1701704242
transform -1 0 2852 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[104\].dly_stg1
timestamp 1701704242
transform -1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[104\].dly_stg2
timestamp 1701704242
transform 1 0 1932 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[105\].dly_stg1
timestamp 1701704242
transform -1 0 1932 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[105\].dly_stg2
timestamp 1701704242
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[106\].dly_stg1
timestamp 1701704242
transform -1 0 2576 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[106\].dly_stg2
timestamp 1701704242
transform -1 0 1472 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[107\].dly_stg1
timestamp 1701704242
transform -1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[107\].dly_stg2
timestamp 1701704242
transform -1 0 1748 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[108\].dly_stg1
timestamp 1701704242
transform 1 0 1012 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[108\].dly_stg2
timestamp 1701704242
transform 1 0 1288 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[109\].dly_stg1
timestamp 1701704242
transform -1 0 1656 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[109\].dly_stg2
timestamp 1701704242
transform -1 0 1932 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[110\].dly_stg1
timestamp 1701704242
transform 1 0 2024 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[110\].dly_stg2
timestamp 1701704242
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[111\].dly_stg1
timestamp 1701704242
transform 1 0 1196 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[111\].dly_stg2
timestamp 1701704242
transform 1 0 1472 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[112\].dly_stg1
timestamp 1701704242
transform 1 0 2024 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[112\].dly_stg2
timestamp 1701704242
transform -1 0 1472 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[113\].dly_stg1
timestamp 1701704242
transform -1 0 1748 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[113\].dly_stg2
timestamp 1701704242
transform -1 0 2024 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[114\].dly_stg1
timestamp 1701704242
transform 1 0 2576 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[114\].dly_stg2
timestamp 1701704242
transform 1 0 2024 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[115\].dly_stg1
timestamp 1701704242
transform -1 0 4232 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[115\].dly_stg2
timestamp 1701704242
transform 1 0 2576 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[116\].dly_stg1
timestamp 1701704242
transform 1 0 3128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[116\].dly_stg2
timestamp 1701704242
transform 1 0 3404 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[117\].dly_stg1
timestamp 1701704242
transform 1 0 3312 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[117\].dly_stg2
timestamp 1701704242
transform -1 0 4232 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[118\].dly_stg1
timestamp 1701704242
transform 1 0 4692 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[118\].dly_stg2
timestamp 1701704242
transform 1 0 3864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[119\].dly_stg1
timestamp 1701704242
transform 1 0 3864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[119\].dly_stg2
timestamp 1701704242
transform 1 0 4140 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[120\].dly_stg1
timestamp 1701704242
transform 1 0 4324 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[120\].dly_stg2
timestamp 1701704242
transform 1 0 4784 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[121\].dly_stg1
timestamp 1701704242
transform 1 0 5060 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[121\].dly_stg2
timestamp 1701704242
transform 1 0 4508 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[122\].dly_stg1
timestamp 1701704242
transform 1 0 4600 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[122\].dly_stg2
timestamp 1701704242
transform 1 0 4232 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[123\].dly_stg1
timestamp 1701704242
transform 1 0 5244 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[123\].dly_stg2
timestamp 1701704242
transform 1 0 5888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[124\].dly_stg1
timestamp 1701704242
transform 1 0 6348 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[124\].dly_stg2
timestamp 1701704242
transform 1 0 6164 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[125\].dly_stg1
timestamp 1701704242
transform -1 0 8556 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[125\].dly_stg2
timestamp 1701704242
transform 1 0 6900 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[126\].dly_stg1
timestamp 1701704242
transform -1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[126\].dly_stg2
timestamp 1701704242
transform -1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[127\].dly_stg1
timestamp 1701704242
transform -1 0 7728 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[127\].dly_stg2
timestamp 1701704242
transform -1 0 7268 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[128\].dly_stg1
timestamp 1701704242
transform -1 0 7452 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[128\].dly_stg2
timestamp 1701704242
transform 1 0 7728 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[129\].dly_stg1
timestamp 1701704242
transform -1 0 6900 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[129\].dly_stg2
timestamp 1701704242
transform -1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[130\].dly_stg1
timestamp 1701704242
transform -1 0 7176 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[130\].dly_stg2
timestamp 1701704242
transform -1 0 7544 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[131\].dly_stg1
timestamp 1701704242
transform -1 0 6716 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[131\].dly_stg2
timestamp 1701704242
transform -1 0 6992 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[132\].dly_stg1
timestamp 1701704242
transform -1 0 7636 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[132\].dly_stg2
timestamp 1701704242
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[133\].dly_stg1
timestamp 1701704242
transform -1 0 6164 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[133\].dly_stg2
timestamp 1701704242
transform -1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[134\].dly_stg1
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[134\].dly_stg2
timestamp 1701704242
transform -1 0 5888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[135\].dly_stg1
timestamp 1701704242
transform -1 0 8924 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[135\].dly_stg2
timestamp 1701704242
transform 1 0 7636 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[136\].dly_stg1
timestamp 1701704242
transform 1 0 8280 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[136\].dly_stg2
timestamp 1701704242
transform 1 0 9016 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[137\].dly_stg1
timestamp 1701704242
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[137\].dly_stg2
timestamp 1701704242
transform 1 0 8924 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[138\].dly_stg1
timestamp 1701704242
transform 1 0 10120 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[138\].dly_stg2
timestamp 1701704242
transform 1 0 9476 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[139\].dly_stg1
timestamp 1701704242
transform 1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[139\].dly_stg2
timestamp 1701704242
transform -1 0 10488 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[140\].dly_stg1
timestamp 1701704242
transform -1 0 10120 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[140\].dly_stg2
timestamp 1701704242
transform -1 0 10028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[141\].dly_stg1
timestamp 1701704242
transform -1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[141\].dly_stg2
timestamp 1701704242
transform -1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[142\].dly_stg1
timestamp 1701704242
transform -1 0 7912 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[142\].dly_stg2
timestamp 1701704242
transform -1 0 7452 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[143\].dly_stg1
timestamp 1701704242
transform -1 0 6624 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[143\].dly_stg2
timestamp 1701704242
transform -1 0 7176 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[144\].dly_stg1
timestamp 1701704242
transform -1 0 5520 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[144\].dly_stg2
timestamp 1701704242
transform -1 0 6072 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[145\].dly_stg1
timestamp 1701704242
transform -1 0 5336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[145\].dly_stg2
timestamp 1701704242
transform -1 0 5060 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[146\].dly_stg1
timestamp 1701704242
transform -1 0 4140 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[146\].dly_stg2
timestamp 1701704242
transform -1 0 4140 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[147\].dly_stg1
timestamp 1701704242
transform -1 0 2944 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[147\].dly_stg2
timestamp 1701704242
transform -1 0 3220 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[148\].dly_stg1
timestamp 1701704242
transform -1 0 2392 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[148\].dly_stg2
timestamp 1701704242
transform 1 0 2668 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[149\].dly_stg1
timestamp 1701704242
transform -1 0 1840 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[149\].dly_stg2
timestamp 1701704242
transform -1 0 2116 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[150\].dly_stg1
timestamp 1701704242
transform -1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[150\].dly_stg2
timestamp 1701704242
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[151\].dly_stg1
timestamp 1701704242
transform 1 0 2208 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[151\].dly_stg2
timestamp 1701704242
transform -1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[152\].dly_stg1
timestamp 1701704242
transform -1 0 2392 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[152\].dly_stg2
timestamp 1701704242
transform -1 0 2116 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[153\].dly_stg1
timestamp 1701704242
transform -1 0 2208 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[153\].dly_stg2
timestamp 1701704242
transform 1 0 1564 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[154\].dly_stg1
timestamp 1701704242
transform -1 0 2852 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[154\].dly_stg2
timestamp 1701704242
transform 1 0 2300 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[155\].dly_stg1
timestamp 1701704242
transform 1 0 2576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[155\].dly_stg2
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[156\].dly_stg1
timestamp 1701704242
transform 1 0 3956 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[156\].dly_stg2
timestamp 1701704242
transform 1 0 3404 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[157\].dly_stg1
timestamp 1701704242
transform -1 0 5336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[157\].dly_stg2
timestamp 1701704242
transform 1 0 4600 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[158\].dly_stg1
timestamp 1701704242
transform 1 0 5428 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[158\].dly_stg2
timestamp 1701704242
transform 1 0 5152 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[159\].dly_stg1
timestamp 1701704242
transform 1 0 6808 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[159\].dly_stg2
timestamp 1701704242
transform 1 0 6256 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[160\].dly_stg1
timestamp 1701704242
transform 1 0 7176 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[160\].dly_stg2
timestamp 1701704242
transform 1 0 7360 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[161\].dly_stg1
timestamp 1701704242
transform 1 0 7544 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[161\].dly_stg2
timestamp 1701704242
transform 1 0 7728 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[162\].dly_stg1
timestamp 1701704242
transform 1 0 7820 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[162\].dly_stg2
timestamp 1701704242
transform 1 0 8372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[163\].dly_stg1
timestamp 1701704242
transform -1 0 9568 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[163\].dly_stg2
timestamp 1701704242
transform 1 0 8648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[164\].dly_stg1
timestamp 1701704242
transform 1 0 9568 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[164\].dly_stg2
timestamp 1701704242
transform 1 0 9200 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[165\].dly_stg1
timestamp 1701704242
transform -1 0 10580 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[165\].dly_stg2
timestamp 1701704242
transform 1 0 9752 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[166\].dly_stg1
timestamp 1701704242
transform 1 0 11868 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[166\].dly_stg2
timestamp 1701704242
transform 1 0 10948 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[167\].dly_stg1
timestamp 1701704242
transform 1 0 12512 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[167\].dly_stg2
timestamp 1701704242
transform 1 0 12604 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[168\].dly_stg1
timestamp 1701704242
transform 1 0 13248 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[168\].dly_stg2
timestamp 1701704242
transform 1 0 12972 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[169\].dly_stg1
timestamp 1701704242
transform -1 0 14628 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[169\].dly_stg2
timestamp 1701704242
transform 1 0 14628 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[170\].dly_stg1
timestamp 1701704242
transform 1 0 14628 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[170\].dly_stg2
timestamp 1701704242
transform 1 0 14352 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[171\].dly_stg1
timestamp 1701704242
transform -1 0 16008 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[171\].dly_stg2
timestamp 1701704242
transform 1 0 15180 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[172\].dly_stg1
timestamp 1701704242
transform 1 0 16284 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[172\].dly_stg2
timestamp 1701704242
transform 1 0 16008 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[173\].dly_stg1
timestamp 1701704242
transform 1 0 17296 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[173\].dly_stg2
timestamp 1701704242
transform 1 0 17204 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[174\].dly_stg1
timestamp 1701704242
transform 1 0 18676 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[174\].dly_stg2
timestamp 1701704242
transform 1 0 17940 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[175\].dly_stg1
timestamp 1701704242
transform 1 0 19504 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[175\].dly_stg2
timestamp 1701704242
transform 1 0 19228 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[176\].dly_stg1
timestamp 1701704242
transform 1 0 19688 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[176\].dly_stg2
timestamp 1701704242
transform 1 0 20608 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[177\].dly_stg1
timestamp 1701704242
transform 1 0 20884 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[177\].dly_stg2
timestamp 1701704242
transform 1 0 20332 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[178\].dly_stg1
timestamp 1701704242
transform 1 0 21528 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[178\].dly_stg2
timestamp 1701704242
transform 1 0 21252 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[179\].dly_stg1
timestamp 1701704242
transform 1 0 22080 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[179\].dly_stg2
timestamp 1701704242
transform 1 0 22356 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[180\].dly_stg1
timestamp 1701704242
transform 1 0 22908 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[180\].dly_stg2
timestamp 1701704242
transform 1 0 22632 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[181\].dly_stg1
timestamp 1701704242
transform -1 0 24656 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[181\].dly_stg2
timestamp 1701704242
transform 1 0 24104 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[182\].dly_stg1
timestamp 1701704242
transform 1 0 23828 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[182\].dly_stg2
timestamp 1701704242
transform -1 0 24656 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[183\].dly_stg1
timestamp 1701704242
transform 1 0 25300 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[183\].dly_stg2
timestamp 1701704242
transform -1 0 24196 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[184\].dly_stg1
timestamp 1701704242
transform 1 0 25576 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[184\].dly_stg2
timestamp 1701704242
transform -1 0 26036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[185\].dly_stg1
timestamp 1701704242
transform 1 0 26128 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[185\].dly_stg2
timestamp 1701704242
transform 1 0 25300 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[186\].dly_stg1
timestamp 1701704242
transform 1 0 26496 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[186\].dly_stg2
timestamp 1701704242
transform 1 0 26772 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[187\].dly_stg1
timestamp 1701704242
transform 1 0 26772 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[187\].dly_stg2
timestamp 1701704242
transform 1 0 27416 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[188\].dly_stg1
timestamp 1701704242
transform 1 0 28980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[188\].dly_stg2
timestamp 1701704242
transform 1 0 27140 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[189\].dly_stg1
timestamp 1701704242
transform 1 0 28428 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[189\].dly_stg2
timestamp 1701704242
transform -1 0 29164 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[190\].dly_stg1
timestamp 1701704242
transform 1 0 29532 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[190\].dly_stg2
timestamp 1701704242
transform 1 0 29256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[191\].dly_stg1
timestamp 1701704242
transform -1 0 28980 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[191\].dly_stg2
timestamp 1701704242
transform 1 0 30360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 30820 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_8
timestamp 1701704242
transform -1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_9
timestamp 1701704242
transform -1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_10
timestamp 1701704242
transform -1 0 8096 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_11
timestamp 1701704242
transform 1 0 30820 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_12
timestamp 1701704242
transform 1 0 30820 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_13
timestamp 1701704242
transform -1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_14
timestamp 1701704242
transform 1 0 30544 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_15
timestamp 1701704242
transform 1 0 30820 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_16
timestamp 1701704242
transform -1 0 6808 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_17
timestamp 1701704242
transform -1 0 7452 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_18
timestamp 1701704242
transform -1 0 28704 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_19
timestamp 1701704242
transform -1 0 1656 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_20
timestamp 1701704242
transform -1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_21
timestamp 1701704242
transform -1 0 28060 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v1_22
timestamp 1701704242
transform 1 0 30820 0 -1 19040
box -38 -48 314 592
<< labels >>
flabel metal4 s 8096 496 8416 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15801 496 16121 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23506 496 23826 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 31211 496 31531 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4244 496 4564 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11949 496 12269 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19654 496 19974 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 27359 496 27679 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 1306 0 1362 400 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 18 0 74 400 0 FreeSans 224 90 0 0 ena
port 3 nsew signal input
flabel metal2 s 662 0 718 400 0 FreeSans 224 90 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 31600 10208 32000 10328 0 FreeSans 480 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal2 s 1950 0 2006 400 0 FreeSans 224 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal2 s 2594 0 2650 400 0 FreeSans 224 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal2 s 16118 0 16174 400 0 FreeSans 224 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal2 s 17406 0 17462 400 0 FreeSans 224 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal2 s 18050 0 18106 400 0 FreeSans 224 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal2 s 3238 0 3294 400 0 FreeSans 224 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal2 s 3882 0 3938 400 0 FreeSans 224 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal2 s 4526 0 4582 400 0 FreeSans 224 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal2 s 5170 0 5226 400 0 FreeSans 224 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal2 s 5814 0 5870 400 0 FreeSans 224 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal2 s 6458 0 6514 400 0 FreeSans 224 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal2 s 7102 0 7158 400 0 FreeSans 224 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal2 s 7746 0 7802 400 0 FreeSans 224 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 31600 2048 32000 2168 0 FreeSans 480 0 0 0 uio_oe[0]
port 21 nsew signal tristate
flabel metal3 s 0 17008 400 17128 0 FreeSans 480 0 0 0 uio_oe[1]
port 22 nsew signal tristate
flabel metal3 s 0 17688 400 17808 0 FreeSans 480 0 0 0 uio_oe[2]
port 23 nsew signal tristate
flabel metal2 s 7746 19600 7802 20000 0 FreeSans 224 90 0 0 uio_oe[3]
port 24 nsew signal tristate
flabel metal3 s 31600 1368 32000 1488 0 FreeSans 480 0 0 0 uio_oe[4]
port 25 nsew signal tristate
flabel metal3 s 31600 688 32000 808 0 FreeSans 480 0 0 0 uio_oe[5]
port 26 nsew signal tristate
flabel metal3 s 0 19728 400 19848 0 FreeSans 480 0 0 0 uio_oe[6]
port 27 nsew signal tristate
flabel metal3 s 31600 19048 32000 19168 0 FreeSans 480 0 0 0 uio_oe[7]
port 28 nsew signal tristate
flabel metal3 s 31600 2728 32000 2848 0 FreeSans 480 0 0 0 uio_out[0]
port 29 nsew signal tristate
flabel metal2 s 6458 19600 6514 20000 0 FreeSans 224 90 0 0 uio_out[1]
port 30 nsew signal tristate
flabel metal2 s 7102 19600 7158 20000 0 FreeSans 224 90 0 0 uio_out[2]
port 31 nsew signal tristate
flabel metal2 s 28354 19600 28410 20000 0 FreeSans 224 90 0 0 uio_out[3]
port 32 nsew signal tristate
flabel metal3 s 0 19048 400 19168 0 FreeSans 480 0 0 0 uio_out[4]
port 33 nsew signal tristate
flabel metal3 s 0 18368 400 18488 0 FreeSans 480 0 0 0 uio_out[5]
port 34 nsew signal tristate
flabel metal2 s 27710 19600 27766 20000 0 FreeSans 224 90 0 0 uio_out[6]
port 35 nsew signal tristate
flabel metal3 s 31600 18368 32000 18488 0 FreeSans 480 0 0 0 uio_out[7]
port 36 nsew signal tristate
flabel metal2 s 19982 19600 20038 20000 0 FreeSans 224 90 0 0 uo_out[0]
port 37 nsew signal tristate
flabel metal3 s 31600 9528 32000 9648 0 FreeSans 480 0 0 0 uo_out[1]
port 38 nsew signal tristate
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 224 90 0 0 uo_out[2]
port 39 nsew signal tristate
flabel metal2 s 18050 19600 18106 20000 0 FreeSans 224 90 0 0 uo_out[3]
port 40 nsew signal tristate
flabel metal2 s 18694 19600 18750 20000 0 FreeSans 224 90 0 0 uo_out[4]
port 41 nsew signal tristate
flabel metal3 s 31600 12248 32000 12368 0 FreeSans 480 0 0 0 uo_out[5]
port 42 nsew signal tristate
flabel metal2 s 19338 19600 19394 20000 0 FreeSans 224 90 0 0 uo_out[6]
port 43 nsew signal tristate
flabel metal2 s 20626 19600 20682 20000 0 FreeSans 224 90 0 0 uo_out[7]
port 44 nsew signal tristate
rlabel via1 16041 19040 16041 19040 0 VGND
rlabel metal1 15962 18496 15962 18496 0 VPWR
rlabel metal1 17802 6086 17802 6086 0 _000_
rlabel metal1 18676 7922 18676 7922 0 _001_
rlabel metal1 18814 8806 18814 8806 0 _002_
rlabel metal1 18998 12954 18998 12954 0 _003_
rlabel metal2 23046 12478 23046 12478 0 _004_
rlabel metal2 15502 4726 15502 4726 0 _005_
rlabel metal1 15594 7242 15594 7242 0 _006_
rlabel viali 13166 7276 13166 7276 0 _007_
rlabel metal1 5198 10472 5198 10472 0 _008_
rlabel metal1 17388 6902 17388 6902 0 _009_
rlabel metal1 24150 11594 24150 11594 0 _010_
rlabel metal1 19964 12750 19964 12750 0 _011_
rlabel metal1 16330 11220 16330 11220 0 _012_
rlabel metal1 15272 6902 15272 6902 0 _013_
rlabel metal2 20470 9537 20470 9537 0 _014_
rlabel metal2 19734 10489 19734 10489 0 _015_
rlabel metal2 20378 11220 20378 11220 0 _016_
rlabel metal1 20746 12954 20746 12954 0 _017_
rlabel metal1 17756 8058 17756 8058 0 _018_
rlabel metal2 17894 5865 17894 5865 0 _019_
rlabel metal1 17848 13430 17848 13430 0 _020_
rlabel metal2 16698 8228 16698 8228 0 _021_
rlabel metal1 15548 7922 15548 7922 0 _022_
rlabel metal1 12512 7922 12512 7922 0 _023_
rlabel metal1 13478 7752 13478 7752 0 _024_
rlabel metal1 12006 8874 12006 8874 0 _025_
rlabel metal1 15824 7446 15824 7446 0 _026_
rlabel metal1 9200 8806 9200 8806 0 _027_
rlabel metal1 8970 10472 8970 10472 0 _028_
rlabel metal1 18676 12342 18676 12342 0 _029_
rlabel metal1 17710 6256 17710 6256 0 _030_
rlabel metal1 23027 5814 23027 5814 0 _031_
rlabel metal2 17158 10200 17158 10200 0 _032_
rlabel metal1 18914 6086 18914 6086 0 _033_
rlabel metal1 17204 10778 17204 10778 0 _034_
rlabel metal1 14122 6834 14122 6834 0 _035_
rlabel metal1 17020 9690 17020 9690 0 _036_
rlabel metal1 16790 9690 16790 9690 0 _037_
rlabel metal1 19826 3366 19826 3366 0 _038_
rlabel metal2 19918 10285 19918 10285 0 _039_
rlabel metal1 14598 3978 14598 3978 0 _040_
rlabel metal1 13984 4794 13984 4794 0 _041_
rlabel metal1 16744 4726 16744 4726 0 _042_
rlabel metal1 14549 4998 14549 4998 0 _043_
rlabel metal1 13892 3706 13892 3706 0 _044_
rlabel via2 14030 6443 14030 6443 0 _045_
rlabel metal1 14352 6426 14352 6426 0 _046_
rlabel metal1 14490 7718 14490 7718 0 _047_
rlabel metal1 16928 13362 16928 13362 0 _048_
rlabel metal1 17112 13362 17112 13362 0 _049_
rlabel metal2 13478 4896 13478 4896 0 _050_
rlabel metal1 12160 3978 12160 3978 0 _051_
rlabel metal3 18055 12988 18055 12988 0 _052_
rlabel metal1 17342 13158 17342 13158 0 _053_
rlabel metal1 17204 8806 17204 8806 0 _054_
rlabel via1 23232 12274 23232 12274 0 _055_
rlabel metal1 14430 3604 14430 3604 0 _056_
rlabel metal1 16744 11798 16744 11798 0 _057_
rlabel metal1 14766 10744 14766 10744 0 _058_
rlabel viali 16974 12277 16974 12277 0 _059_
rlabel metal1 12834 6426 12834 6426 0 _060_
rlabel metal3 17411 11764 17411 11764 0 _061_
rlabel metal1 16606 11662 16606 11662 0 _062_
rlabel metal1 19918 11832 19918 11832 0 _063_
rlabel metal1 18722 10064 18722 10064 0 _064_
rlabel metal1 18262 9044 18262 9044 0 _065_
rlabel metal1 20148 15130 20148 15130 0 _066_
rlabel metal2 24150 12410 24150 12410 0 _067_
rlabel metal2 21482 14025 21482 14025 0 _068_
rlabel metal2 21068 9418 21068 9418 0 _069_
rlabel metal2 20562 9316 20562 9316 0 _070_
rlabel metal1 21206 9588 21206 9588 0 _071_
rlabel metal2 19136 8636 19136 8636 0 _072_
rlabel metal1 14674 3468 14674 3468 0 _073_
rlabel metal1 14260 9894 14260 9894 0 _074_
rlabel metal2 14812 9486 14812 9486 0 _075_
rlabel metal1 13164 12614 13164 12614 0 _076_
rlabel metal1 14996 6834 14996 6834 0 _077_
rlabel metal1 17112 5882 17112 5882 0 _078_
rlabel metal2 14582 5066 14582 5066 0 _079_
rlabel metal1 14720 6970 14720 6970 0 _080_
rlabel metal1 15364 9894 15364 9894 0 _081_
rlabel metal2 21344 6596 21344 6596 0 _082_
rlabel metal1 14628 6358 14628 6358 0 _083_
rlabel viali 14774 9554 14774 9554 0 _084_
rlabel metal1 12190 9486 12190 9486 0 _085_
rlabel metal1 12466 9554 12466 9554 0 _086_
rlabel metal2 12742 9316 12742 9316 0 _087_
rlabel metal2 11684 4522 11684 4522 0 _088_
rlabel metal1 13846 9418 13846 9418 0 _089_
rlabel metal2 19918 8925 19918 8925 0 _090_
rlabel metal1 9890 11730 9890 11730 0 _091_
rlabel metal3 16284 11288 16284 11288 0 _092_
rlabel metal2 16652 11186 16652 11186 0 _093_
rlabel metal1 17618 11220 17618 11220 0 _094_
rlabel metal1 18170 8806 18170 8806 0 _095_
rlabel metal1 18262 8058 18262 8058 0 _096_
rlabel metal1 17756 8398 17756 8398 0 _097_
rlabel metal1 14950 5338 14950 5338 0 _098_
rlabel metal1 15042 8534 15042 8534 0 _099_
rlabel metal1 15134 8602 15134 8602 0 _100_
rlabel metal1 16100 8466 16100 8466 0 _101_
rlabel metal1 16560 4182 16560 4182 0 _102_
rlabel metal1 21574 3706 21574 3706 0 _103_
rlabel metal1 17480 3706 17480 3706 0 _104_
rlabel metal1 17618 4250 17618 4250 0 _105_
rlabel metal2 25346 8704 25346 8704 0 _106_
rlabel metal1 24242 8500 24242 8500 0 _107_
rlabel metal1 24242 4250 24242 4250 0 _108_
rlabel metal1 20118 8364 20118 8364 0 _109_
rlabel metal1 17756 8602 17756 8602 0 _110_
rlabel metal1 18124 12410 18124 12410 0 _111_
rlabel metal2 17986 10846 17986 10846 0 _112_
rlabel metal1 16146 8908 16146 8908 0 _113_
rlabel metal2 16606 9792 16606 9792 0 _114_
rlabel metal1 18262 7888 18262 7888 0 _115_
rlabel metal1 13110 3434 13110 3434 0 _116_
rlabel metal1 14904 9078 14904 9078 0 _117_
rlabel metal2 19366 13532 19366 13532 0 _118_
rlabel metal1 14490 13260 14490 13260 0 _119_
rlabel metal1 14674 13362 14674 13362 0 _120_
rlabel metal2 14950 12716 14950 12716 0 _121_
rlabel metal1 12926 6732 12926 6732 0 _122_
rlabel metal2 15134 4607 15134 4607 0 _123_
rlabel metal2 12926 7616 12926 7616 0 _124_
rlabel metal1 13386 8058 13386 8058 0 _125_
rlabel metal1 23782 9894 23782 9894 0 _126_
rlabel metal2 24702 13333 24702 13333 0 _127_
rlabel metal1 23782 9962 23782 9962 0 _128_
rlabel via2 23230 9979 23230 9979 0 _129_
rlabel metal1 17526 9486 17526 9486 0 _130_
rlabel metal1 5842 11118 5842 11118 0 _131_
rlabel metal2 18446 11781 18446 11781 0 _132_
rlabel metal2 20562 5644 20562 5644 0 _133_
rlabel metal1 16652 10778 16652 10778 0 _134_
rlabel metal1 13386 5236 13386 5236 0 _135_
rlabel metal1 19918 5338 19918 5338 0 _136_
rlabel metal1 18446 11560 18446 11560 0 _137_
rlabel metal1 12788 13158 12788 13158 0 _138_
rlabel metal1 13340 13226 13340 13226 0 _139_
rlabel metal1 13938 13158 13938 13158 0 _140_
rlabel metal1 15272 13498 15272 13498 0 _141_
rlabel metal1 18446 4658 18446 4658 0 _142_
rlabel metal1 13846 4488 13846 4488 0 _143_
rlabel metal1 18308 4250 18308 4250 0 _144_
rlabel metal1 18400 11730 18400 11730 0 _145_
rlabel metal1 23276 14042 23276 14042 0 _146_
rlabel metal1 23000 14042 23000 14042 0 _147_
rlabel metal1 22862 13974 22862 13974 0 _148_
rlabel metal2 18262 11866 18262 11866 0 _149_
rlabel metal1 19090 11628 19090 11628 0 _150_
rlabel metal2 18262 14688 18262 14688 0 _151_
rlabel metal1 24334 14246 24334 14246 0 _152_
rlabel metal2 13662 4947 13662 4947 0 _153_
rlabel metal1 24150 12308 24150 12308 0 _154_
rlabel metal1 13754 8058 13754 8058 0 _155_
rlabel metal1 13662 8534 13662 8534 0 _156_
rlabel metal1 13800 8602 13800 8602 0 _157_
rlabel metal1 19320 8058 19320 8058 0 _158_
rlabel metal1 19596 8534 19596 8534 0 _159_
rlabel metal1 20056 8058 20056 8058 0 _160_
rlabel metal1 13800 8806 13800 8806 0 _161_
rlabel metal1 14536 4794 14536 4794 0 _162_
rlabel metal1 12926 2856 12926 2856 0 _163_
rlabel metal1 13248 6426 13248 6426 0 _164_
rlabel metal2 13110 7888 13110 7888 0 _165_
rlabel metal1 12742 8602 12742 8602 0 _166_
rlabel metal2 12098 5066 12098 5066 0 _167_
rlabel metal4 13708 6188 13708 6188 0 _168_
rlabel metal2 13018 8806 13018 8806 0 _169_
rlabel via2 13478 8891 13478 8891 0 _170_
rlabel metal1 5612 10778 5612 10778 0 _171_
rlabel metal2 19366 11951 19366 11951 0 _172_
rlabel metal2 15318 13022 15318 13022 0 _173_
rlabel metal1 19458 12240 19458 12240 0 _174_
rlabel metal1 19366 9554 19366 9554 0 _175_
rlabel metal1 20010 4182 20010 4182 0 _176_
rlabel metal1 19596 9486 19596 9486 0 _177_
rlabel metal1 13616 7514 13616 7514 0 _178_
rlabel metal2 13202 6358 13202 6358 0 _179_
rlabel metal1 13892 9622 13892 9622 0 _180_
rlabel metal2 14904 7820 14904 7820 0 _181_
rlabel metal1 14536 4182 14536 4182 0 _182_
rlabel metal1 21160 4250 21160 4250 0 _183_
rlabel metal1 20470 3706 20470 3706 0 _184_
rlabel metal1 19780 6222 19780 6222 0 _185_
rlabel metal1 24656 8806 24656 8806 0 _186_
rlabel metal1 24242 8806 24242 8806 0 _187_
rlabel metal2 23690 8738 23690 8738 0 _188_
rlabel metal1 21942 9384 21942 9384 0 _189_
rlabel metal1 19596 9622 19596 9622 0 _190_
rlabel metal1 8050 11322 8050 11322 0 _191_
rlabel metal3 14628 12920 14628 12920 0 _192_
rlabel metal2 24472 13668 24472 13668 0 _193_
rlabel metal1 20470 12716 20470 12716 0 _194_
rlabel metal2 15318 4743 15318 4743 0 _195_
rlabel metal1 20562 5338 20562 5338 0 _196_
rlabel metal1 19918 12682 19918 12682 0 _197_
rlabel metal1 13616 12886 13616 12886 0 _198_
rlabel metal3 14007 12580 14007 12580 0 _199_
rlabel metal2 14030 13328 14030 13328 0 _200_
rlabel metal1 15410 12954 15410 12954 0 _201_
rlabel metal3 19504 5644 19504 5644 0 _202_
rlabel metal2 13846 3672 13846 3672 0 _203_
rlabel metal2 19366 4080 19366 4080 0 _204_
rlabel metal1 19550 4794 19550 4794 0 _205_
rlabel metal1 15962 13940 15962 13940 0 _206_
rlabel metal1 20010 13974 20010 13974 0 _207_
rlabel metal1 19274 13974 19274 13974 0 _208_
rlabel metal2 19274 13226 19274 13226 0 _209_
rlabel metal1 20562 12784 20562 12784 0 _210_
rlabel metal2 1334 5260 1334 5260 0 clk
rlabel metal2 12466 7105 12466 7105 0 clknet_0_clk
rlabel metal1 1150 5780 1150 5780 0 clknet_4_0_0_clk
rlabel metal1 25208 2958 25208 2958 0 clknet_4_10_0_clk
rlabel metal1 28842 10030 28842 10030 0 clknet_4_11_0_clk
rlabel metal1 17848 16626 17848 16626 0 clknet_4_12_0_clk
rlabel metal1 16330 17646 16330 17646 0 clknet_4_13_0_clk
rlabel metal1 27278 12682 27278 12682 0 clknet_4_14_0_clk
rlabel metal1 29578 14450 29578 14450 0 clknet_4_15_0_clk
rlabel metal1 2070 6834 2070 6834 0 clknet_4_1_0_clk
rlabel metal1 14582 2516 14582 2516 0 clknet_4_2_0_clk
rlabel metal1 8878 7378 8878 7378 0 clknet_4_3_0_clk
rlabel metal2 1702 13022 1702 13022 0 clknet_4_4_0_clk
rlabel metal2 2714 14212 2714 14212 0 clknet_4_5_0_clk
rlabel metal1 14582 12750 14582 12750 0 clknet_4_6_0_clk
rlabel metal1 11546 15572 11546 15572 0 clknet_4_7_0_clk
rlabel metal2 20102 2448 20102 2448 0 clknet_4_8_0_clk
rlabel metal1 21344 5746 21344 5746 0 clknet_4_9_0_clk
rlabel metal1 25530 10642 25530 10642 0 net1
rlabel metal1 7820 18802 7820 18802 0 net10
rlabel metal3 31380 1428 31380 1428 0 net11
rlabel metal3 31380 748 31380 748 0 net12
rlabel metal2 1150 19261 1150 19261 0 net13
rlabel metal1 31234 18802 31234 18802 0 net14
rlabel via2 31702 2788 31702 2788 0 net15
rlabel metal1 6532 18802 6532 18802 0 net16
rlabel metal1 7176 18802 7176 18802 0 net17
rlabel metal1 28428 18802 28428 18802 0 net18
rlabel metal1 1104 18802 1104 18802 0 net19
rlabel metal1 18078 5576 18078 5576 0 net2
rlabel metal3 590 18428 590 18428 0 net20
rlabel metal1 27784 18802 27784 18802 0 net21
rlabel metal3 31380 18428 31380 18428 0 net22
rlabel via1 29297 5134 29297 5134 0 net23
rlabel metal1 30600 5746 30600 5746 0 net24
rlabel metal1 29844 6222 29844 6222 0 net25
rlabel metal2 30314 7786 30314 7786 0 net26
rlabel metal1 28198 7514 28198 7514 0 net27
rlabel metal1 28300 5746 28300 5746 0 net28
rlabel metal1 16882 5780 16882 5780 0 net3
rlabel metal1 17572 7310 17572 7310 0 net4
rlabel metal1 17894 6222 17894 6222 0 net5
rlabel metal1 18492 5610 18492 5610 0 net6
rlabel metal3 31380 2108 31380 2108 0 net7
rlabel metal3 590 17068 590 17068 0 net8
rlabel metal3 590 17748 590 17748 0 net9
rlabel metal1 21367 11730 21367 11730 0 tdc0.o_result\[0\]
rlabel metal2 6118 17238 6118 17238 0 tdc0.o_result\[100\]
rlabel metal2 19182 8449 19182 8449 0 tdc0.o_result\[101\]
rlabel metal1 5704 15334 5704 15334 0 tdc0.o_result\[102\]
rlabel metal2 6394 14149 6394 14149 0 tdc0.o_result\[103\]
rlabel metal2 16790 13447 16790 13447 0 tdc0.o_result\[104\]
rlabel metal1 4784 14586 4784 14586 0 tdc0.o_result\[105\]
rlabel metal2 13846 11713 13846 11713 0 tdc0.o_result\[106\]
rlabel metal2 3082 12461 3082 12461 0 tdc0.o_result\[107\]
rlabel metal1 4830 11254 4830 11254 0 tdc0.o_result\[108\]
rlabel metal1 2346 6120 2346 6120 0 tdc0.o_result\[109\]
rlabel metal1 26128 9078 26128 9078 0 tdc0.o_result\[10\]
rlabel metal1 5290 10608 5290 10608 0 tdc0.o_result\[110\]
rlabel metal2 15594 13515 15594 13515 0 tdc0.o_result\[111\]
rlabel metal1 4186 9894 4186 9894 0 tdc0.o_result\[112\]
rlabel metal1 11454 7480 11454 7480 0 tdc0.o_result\[113\]
rlabel metal1 5658 9112 5658 9112 0 tdc0.o_result\[114\]
rlabel metal1 12650 7956 12650 7956 0 tdc0.o_result\[115\]
rlabel viali 5934 11186 5934 11186 0 tdc0.o_result\[116\]
rlabel metal1 13340 8262 13340 8262 0 tdc0.o_result\[117\]
rlabel viali 5750 11662 5750 11662 0 tdc0.o_result\[118\]
rlabel viali 6302 12274 6302 12274 0 tdc0.o_result\[119\]
rlabel metal2 24426 10608 24426 10608 0 tdc0.o_result\[11\]
rlabel metal1 9338 9078 9338 9078 0 tdc0.o_result\[120\]
rlabel via2 18722 14909 18722 14909 0 tdc0.o_result\[121\]
rlabel metal1 7406 13158 7406 13158 0 tdc0.o_result\[122\]
rlabel metal1 7958 14552 7958 14552 0 tdc0.o_result\[123\]
rlabel metal1 12742 13736 12742 13736 0 tdc0.o_result\[124\]
rlabel metal2 17710 14977 17710 14977 0 tdc0.o_result\[125\]
rlabel metal1 13110 9350 13110 9350 0 tdc0.o_result\[126\]
rlabel metal1 13754 12784 13754 12784 0 tdc0.o_result\[127\]
rlabel metal1 8234 10574 8234 10574 0 tdc0.o_result\[128\]
rlabel metal1 11178 9112 11178 9112 0 tdc0.o_result\[129\]
rlabel metal1 23966 5304 23966 5304 0 tdc0.o_result\[12\]
rlabel metal1 11454 8466 11454 8466 0 tdc0.o_result\[130\]
rlabel metal1 11362 7242 11362 7242 0 tdc0.o_result\[131\]
rlabel metal1 5796 8602 5796 8602 0 tdc0.o_result\[132\]
rlabel metal1 8602 6936 8602 6936 0 tdc0.o_result\[133\]
rlabel metal1 11546 7208 11546 7208 0 tdc0.o_result\[134\]
rlabel metal1 8096 7446 8096 7446 0 tdc0.o_result\[135\]
rlabel metal1 8418 6392 8418 6392 0 tdc0.o_result\[136\]
rlabel metal1 12374 7820 12374 7820 0 tdc0.o_result\[137\]
rlabel metal1 10994 4148 10994 4148 0 tdc0.o_result\[138\]
rlabel metal3 14375 12852 14375 12852 0 tdc0.o_result\[139\]
rlabel via2 19734 7973 19734 7973 0 tdc0.o_result\[13\]
rlabel metal1 13570 13362 13570 13362 0 tdc0.o_result\[140\]
rlabel metal1 13018 4556 13018 4556 0 tdc0.o_result\[141\]
rlabel metal2 13110 5797 13110 5797 0 tdc0.o_result\[142\]
rlabel metal2 11362 4420 11362 4420 0 tdc0.o_result\[143\]
rlabel metal1 15272 5610 15272 5610 0 tdc0.o_result\[144\]
rlabel metal1 7222 5848 7222 5848 0 tdc0.o_result\[145\]
rlabel metal1 7406 6086 7406 6086 0 tdc0.o_result\[146\]
rlabel metal2 4646 6035 4646 6035 0 tdc0.o_result\[147\]
rlabel via2 4922 4539 4922 4539 0 tdc0.o_result\[148\]
rlabel metal1 12742 5848 12742 5848 0 tdc0.o_result\[149\]
rlabel metal2 26542 8806 26542 8806 0 tdc0.o_result\[14\]
rlabel metal2 3542 8568 3542 8568 0 tdc0.o_result\[150\]
rlabel metal2 7222 4743 7222 4743 0 tdc0.o_result\[151\]
rlabel metal2 3450 4352 3450 4352 0 tdc0.o_result\[152\]
rlabel metal1 5980 3910 5980 3910 0 tdc0.o_result\[153\]
rlabel metal1 8510 3638 8510 3638 0 tdc0.o_result\[154\]
rlabel metal2 5290 2873 5290 2873 0 tdc0.o_result\[155\]
rlabel metal1 8602 2822 8602 2822 0 tdc0.o_result\[156\]
rlabel metal1 8096 3910 8096 3910 0 tdc0.o_result\[157\]
rlabel metal2 12006 3553 12006 3553 0 tdc0.o_result\[158\]
rlabel metal1 9890 3162 9890 3162 0 tdc0.o_result\[159\]
rlabel via2 19918 5797 19918 5797 0 tdc0.o_result\[15\]
rlabel metal2 13478 3570 13478 3570 0 tdc0.o_result\[160\]
rlabel metal2 14214 2958 14214 2958 0 tdc0.o_result\[161\]
rlabel metal1 13110 5032 13110 5032 0 tdc0.o_result\[162\]
rlabel metal1 11224 2618 11224 2618 0 tdc0.o_result\[163\]
rlabel metal2 13018 3570 13018 3570 0 tdc0.o_result\[164\]
rlabel metal1 13064 2618 13064 2618 0 tdc0.o_result\[165\]
rlabel metal1 12742 1530 12742 1530 0 tdc0.o_result\[166\]
rlabel metal1 12696 3162 12696 3162 0 tdc0.o_result\[167\]
rlabel metal1 16146 2618 16146 2618 0 tdc0.o_result\[168\]
rlabel metal1 14858 3638 14858 3638 0 tdc0.o_result\[169\]
rlabel via2 19734 6885 19734 6885 0 tdc0.o_result\[16\]
rlabel metal1 17112 3638 17112 3638 0 tdc0.o_result\[170\]
rlabel metal2 14950 3366 14950 3366 0 tdc0.o_result\[171\]
rlabel metal1 17940 3978 17940 3978 0 tdc0.o_result\[172\]
rlabel metal1 17066 3162 17066 3162 0 tdc0.o_result\[173\]
rlabel metal1 19964 3638 19964 3638 0 tdc0.o_result\[174\]
rlabel metal1 19734 3604 19734 3604 0 tdc0.o_result\[175\]
rlabel metal1 19228 3638 19228 3638 0 tdc0.o_result\[176\]
rlabel metal1 21620 3638 21620 3638 0 tdc0.o_result\[177\]
rlabel metal1 22080 3638 22080 3638 0 tdc0.o_result\[178\]
rlabel metal1 24242 4012 24242 4012 0 tdc0.o_result\[179\]
rlabel metal1 19642 5814 19642 5814 0 tdc0.o_result\[17\]
rlabel metal1 23828 1530 23828 1530 0 tdc0.o_result\[180\]
rlabel metal1 15318 4726 15318 4726 0 tdc0.o_result\[181\]
rlabel metal1 22402 2040 22402 2040 0 tdc0.o_result\[182\]
rlabel metal2 23368 5746 23368 5746 0 tdc0.o_result\[183\]
rlabel metal1 23368 3978 23368 3978 0 tdc0.o_result\[184\]
rlabel metal1 20511 9418 20511 9418 0 tdc0.o_result\[185\]
rlabel metal1 24656 3978 24656 3978 0 tdc0.o_result\[186\]
rlabel metal1 23322 3604 23322 3604 0 tdc0.o_result\[187\]
rlabel metal2 20010 4828 20010 4828 0 tdc0.o_result\[188\]
rlabel via2 22954 3995 22954 3995 0 tdc0.o_result\[189\]
rlabel metal2 18998 7905 18998 7905 0 tdc0.o_result\[18\]
rlabel metal1 23966 3128 23966 3128 0 tdc0.o_result\[190\]
rlabel metal1 20930 5032 20930 5032 0 tdc0.o_result\[191\]
rlabel metal1 23204 7480 23204 7480 0 tdc0.o_result\[19\]
rlabel metal1 25472 9486 25472 9486 0 tdc0.o_result\[1\]
rlabel metal1 22754 5576 22754 5576 0 tdc0.o_result\[20\]
rlabel metal1 21942 7820 21942 7820 0 tdc0.o_result\[21\]
rlabel metal1 24886 8296 24886 8296 0 tdc0.o_result\[22\]
rlabel metal1 20838 5848 20838 5848 0 tdc0.o_result\[23\]
rlabel metal3 18883 6732 18883 6732 0 tdc0.o_result\[24\]
rlabel metal2 15318 6630 15318 6630 0 tdc0.o_result\[25\]
rlabel metal1 24472 8058 24472 8058 0 tdc0.o_result\[26\]
rlabel metal1 17710 7514 17710 7514 0 tdc0.o_result\[27\]
rlabel metal1 22954 5202 22954 5202 0 tdc0.o_result\[28\]
rlabel metal1 20608 8330 20608 8330 0 tdc0.o_result\[29\]
rlabel metal1 20378 11254 20378 11254 0 tdc0.o_result\[2\]
rlabel metal1 24242 9146 24242 9146 0 tdc0.o_result\[30\]
rlabel metal2 23046 5236 23046 5236 0 tdc0.o_result\[31\]
rlabel metal2 20102 10778 20102 10778 0 tdc0.o_result\[32\]
rlabel metal1 15410 10064 15410 10064 0 tdc0.o_result\[33\]
rlabel metal1 21068 10982 21068 10982 0 tdc0.o_result\[34\]
rlabel metal2 23874 10336 23874 10336 0 tdc0.o_result\[35\]
rlabel metal2 23414 13600 23414 13600 0 tdc0.o_result\[36\]
rlabel metal1 22356 12614 22356 12614 0 tdc0.o_result\[37\]
rlabel metal2 19918 12223 19918 12223 0 tdc0.o_result\[38\]
rlabel metal1 19734 13872 19734 13872 0 tdc0.o_result\[39\]
rlabel metal1 19147 10098 19147 10098 0 tdc0.o_result\[3\]
rlabel metal1 17986 13464 17986 13464 0 tdc0.o_result\[40\]
rlabel metal1 24840 15130 24840 15130 0 tdc0.o_result\[41\]
rlabel via2 17066 11203 17066 11203 0 tdc0.o_result\[42\]
rlabel metal2 20378 13583 20378 13583 0 tdc0.o_result\[43\]
rlabel metal1 29486 14552 29486 14552 0 tdc0.o_result\[44\]
rlabel metal1 24334 14416 24334 14416 0 tdc0.o_result\[45\]
rlabel metal1 22871 4760 22871 4760 0 tdc0.o_result\[46\]
rlabel metal1 25254 14858 25254 14858 0 tdc0.o_result\[47\]
rlabel metal1 24702 11730 24702 11730 0 tdc0.o_result\[48\]
rlabel metal1 24628 15538 24628 15538 0 tdc0.o_result\[49\]
rlabel via1 19722 11662 19722 11662 0 tdc0.o_result\[4\]
rlabel metal4 17204 8908 17204 8908 0 tdc0.o_result\[50\]
rlabel metal1 25024 14518 25024 14518 0 tdc0.o_result\[51\]
rlabel metal2 23230 16014 23230 16014 0 tdc0.o_result\[52\]
rlabel via1 24058 14450 24058 14450 0 tdc0.o_result\[53\]
rlabel metal2 21252 11356 21252 11356 0 tdc0.o_result\[54\]
rlabel metal2 20838 15266 20838 15266 0 tdc0.o_result\[55\]
rlabel metal1 17296 18598 17296 18598 0 tdc0.o_result\[56\]
rlabel metal1 18998 14994 18998 14994 0 tdc0.o_result\[57\]
rlabel metal3 18331 16660 18331 16660 0 tdc0.o_result\[58\]
rlabel metal1 18022 12784 18022 12784 0 tdc0.o_result\[59\]
rlabel metal1 25932 12274 25932 12274 0 tdc0.o_result\[5\]
rlabel metal2 19182 14926 19182 14926 0 tdc0.o_result\[60\]
rlabel metal2 23138 14654 23138 14654 0 tdc0.o_result\[61\]
rlabel metal2 23874 14603 23874 14603 0 tdc0.o_result\[62\]
rlabel via1 23966 14926 23966 14926 0 tdc0.o_result\[63\]
rlabel metal1 17112 13770 17112 13770 0 tdc0.o_result\[64\]
rlabel metal2 20838 9486 20838 9486 0 tdc0.o_result\[65\]
rlabel metal1 21988 13770 21988 13770 0 tdc0.o_result\[66\]
rlabel metal3 16353 15980 16353 15980 0 tdc0.o_result\[67\]
rlabel metal1 22374 14518 22374 14518 0 tdc0.o_result\[68\]
rlabel metal1 17986 14824 17986 14824 0 tdc0.o_result\[69\]
rlabel metal1 22494 12172 22494 12172 0 tdc0.o_result\[6\]
rlabel metal2 18032 12852 18032 12852 0 tdc0.o_result\[70\]
rlabel metal2 13662 14280 13662 14280 0 tdc0.o_result\[71\]
rlabel metal1 16514 12648 16514 12648 0 tdc0.o_result\[72\]
rlabel metal1 12374 9350 12374 9350 0 tdc0.o_result\[73\]
rlabel metal1 13478 11662 13478 11662 0 tdc0.o_result\[74\]
rlabel metal1 16236 9486 16236 9486 0 tdc0.o_result\[75\]
rlabel viali 16330 10575 16330 10575 0 tdc0.o_result\[76\]
rlabel metal1 12466 8432 12466 8432 0 tdc0.o_result\[77\]
rlabel metal1 10718 10064 10718 10064 0 tdc0.o_result\[78\]
rlabel metal1 8786 11152 8786 11152 0 tdc0.o_result\[79\]
rlabel metal1 22218 12852 22218 12852 0 tdc0.o_result\[7\]
rlabel metal2 16652 10506 16652 10506 0 tdc0.o_result\[80\]
rlabel metal1 11546 12682 11546 12682 0 tdc0.o_result\[81\]
rlabel metal2 13938 13260 13938 13260 0 tdc0.o_result\[82\]
rlabel metal2 13754 14450 13754 14450 0 tdc0.o_result\[83\]
rlabel metal1 11730 13464 11730 13464 0 tdc0.o_result\[84\]
rlabel metal2 12972 12308 12972 12308 0 tdc0.o_result\[85\]
rlabel via1 15121 13770 15121 13770 0 tdc0.o_result\[86\]
rlabel metal1 13156 12682 13156 12682 0 tdc0.o_result\[87\]
rlabel viali 17710 13362 17710 13362 0 tdc0.o_result\[88\]
rlabel metal1 14444 10506 14444 10506 0 tdc0.o_result\[89\]
rlabel metal1 29578 11288 29578 11288 0 tdc0.o_result\[8\]
rlabel metal2 14582 11832 14582 11832 0 tdc0.o_result\[90\]
rlabel via3 15019 18020 15019 18020 0 tdc0.o_result\[91\]
rlabel metal1 16055 10608 16055 10608 0 tdc0.o_result\[92\]
rlabel metal2 12558 14552 12558 14552 0 tdc0.o_result\[93\]
rlabel metal2 14858 15062 14858 15062 0 tdc0.o_result\[94\]
rlabel metal3 15548 13668 15548 13668 0 tdc0.o_result\[95\]
rlabel metal1 14582 17544 14582 17544 0 tdc0.o_result\[96\]
rlabel metal2 9430 13702 9430 13702 0 tdc0.o_result\[97\]
rlabel metal2 7774 14421 7774 14421 0 tdc0.o_result\[98\]
rlabel via2 17802 12733 17802 12733 0 tdc0.o_result\[99\]
rlabel metal2 24150 9129 24150 9129 0 tdc0.o_result\[9\]
rlabel metal1 7774 16966 7774 16966 0 tdc0.w_dly_sig\[100\]
rlabel metal1 5382 16762 5382 16762 0 tdc0.w_dly_sig\[101\]
rlabel metal1 6256 16422 6256 16422 0 tdc0.w_dly_sig\[102\]
rlabel metal1 2070 16048 2070 16048 0 tdc0.w_dly_sig\[103\]
rlabel metal1 2254 16626 2254 16626 0 tdc0.w_dly_sig\[104\]
rlabel metal1 2714 15640 2714 15640 0 tdc0.w_dly_sig\[105\]
rlabel metal1 2208 15334 2208 15334 0 tdc0.w_dly_sig\[106\]
rlabel metal1 1978 14790 1978 14790 0 tdc0.w_dly_sig\[107\]
rlabel metal1 1472 14314 1472 14314 0 tdc0.w_dly_sig\[108\]
rlabel metal1 1564 14042 1564 14042 0 tdc0.w_dly_sig\[109\]
rlabel metal1 28934 9894 28934 9894 0 tdc0.w_dly_sig\[10\]
rlabel metal1 1288 12614 1288 12614 0 tdc0.w_dly_sig\[110\]
rlabel metal1 1334 11866 1334 11866 0 tdc0.w_dly_sig\[111\]
rlabel metal1 1876 13362 1876 13362 0 tdc0.w_dly_sig\[112\]
rlabel metal1 1748 9690 1748 9690 0 tdc0.w_dly_sig\[113\]
rlabel metal1 1380 9146 1380 9146 0 tdc0.w_dly_sig\[114\]
rlabel metal1 1472 8874 1472 8874 0 tdc0.w_dly_sig\[115\]
rlabel metal2 2438 8772 2438 8772 0 tdc0.w_dly_sig\[116\]
rlabel metal1 3358 10132 3358 10132 0 tdc0.w_dly_sig\[117\]
rlabel metal1 4554 9690 4554 9690 0 tdc0.w_dly_sig\[118\]
rlabel via1 3721 11662 3721 11662 0 tdc0.w_dly_sig\[119\]
rlabel metal1 29394 9622 29394 9622 0 tdc0.w_dly_sig\[11\]
rlabel metal1 4232 12750 4232 12750 0 tdc0.w_dly_sig\[120\]
rlabel metal1 4876 12614 4876 12614 0 tdc0.w_dly_sig\[121\]
rlabel metal1 4646 14484 4646 14484 0 tdc0.w_dly_sig\[122\]
rlabel metal1 5382 13838 5382 13838 0 tdc0.w_dly_sig\[123\]
rlabel metal2 5014 14144 5014 14144 0 tdc0.w_dly_sig\[124\]
rlabel metal1 5888 13702 5888 13702 0 tdc0.w_dly_sig\[125\]
rlabel metal1 6210 14246 6210 14246 0 tdc0.w_dly_sig\[126\]
rlabel metal1 7222 13702 7222 13702 0 tdc0.w_dly_sig\[127\]
rlabel metal1 7038 12614 7038 12614 0 tdc0.w_dly_sig\[128\]
rlabel metal1 7033 10506 7033 10506 0 tdc0.w_dly_sig\[129\]
rlabel metal1 29987 10166 29987 10166 0 tdc0.w_dly_sig\[12\]
rlabel metal1 7406 9044 7406 9044 0 tdc0.w_dly_sig\[130\]
rlabel metal2 7866 8636 7866 8636 0 tdc0.w_dly_sig\[131\]
rlabel metal1 7590 7956 7590 7956 0 tdc0.w_dly_sig\[132\]
rlabel metal1 5842 7956 5842 7956 0 tdc0.w_dly_sig\[133\]
rlabel metal1 5612 7718 5612 7718 0 tdc0.w_dly_sig\[134\]
rlabel metal1 8924 7310 8924 7310 0 tdc0.w_dly_sig\[135\]
rlabel metal1 6378 7242 6378 7242 0 tdc0.w_dly_sig\[136\]
rlabel metal1 8786 6222 8786 6222 0 tdc0.w_dly_sig\[137\]
rlabel metal1 10258 6222 10258 6222 0 tdc0.w_dly_sig\[138\]
rlabel metal1 10166 5542 10166 5542 0 tdc0.w_dly_sig\[139\]
rlabel metal1 29624 7310 29624 7310 0 tdc0.w_dly_sig\[13\]
rlabel metal2 10534 6630 10534 6630 0 tdc0.w_dly_sig\[140\]
rlabel metal2 10350 5984 10350 5984 0 tdc0.w_dly_sig\[141\]
rlabel via1 9517 4726 9517 4726 0 tdc0.w_dly_sig\[142\]
rlabel metal1 9752 4998 9752 4998 0 tdc0.w_dly_sig\[143\]
rlabel metal1 7360 4998 7360 4998 0 tdc0.w_dly_sig\[144\]
rlabel metal1 8142 5338 8142 5338 0 tdc0.w_dly_sig\[145\]
rlabel metal1 4232 6222 4232 6222 0 tdc0.w_dly_sig\[146\]
rlabel metal1 3726 6256 3726 6256 0 tdc0.w_dly_sig\[147\]
rlabel metal1 2438 5100 2438 5100 0 tdc0.w_dly_sig\[148\]
rlabel metal2 1978 4964 1978 4964 0 tdc0.w_dly_sig\[149\]
rlabel metal1 29378 7990 29378 7990 0 tdc0.w_dly_sig\[14\]
rlabel metal1 1324 5746 1324 5746 0 tdc0.w_dly_sig\[150\]
rlabel metal1 2116 5338 2116 5338 0 tdc0.w_dly_sig\[151\]
rlabel metal1 1794 4250 1794 4250 0 tdc0.w_dly_sig\[152\]
rlabel metal1 1242 4046 1242 4046 0 tdc0.w_dly_sig\[153\]
rlabel metal2 2530 3842 2530 3842 0 tdc0.w_dly_sig\[154\]
rlabel metal2 2806 2176 2806 2176 0 tdc0.w_dly_sig\[155\]
rlabel metal2 2438 2720 2438 2720 0 tdc0.w_dly_sig\[156\]
rlabel metal1 5336 2482 5336 2482 0 tdc0.w_dly_sig\[157\]
rlabel metal1 4646 1836 4646 1836 0 tdc0.w_dly_sig\[158\]
rlabel metal1 5934 1938 5934 1938 0 tdc0.w_dly_sig\[159\]
rlabel metal1 29670 6970 29670 6970 0 tdc0.w_dly_sig\[15\]
rlabel metal1 7130 2482 7130 2482 0 tdc0.w_dly_sig\[160\]
rlabel metal1 6808 2074 6808 2074 0 tdc0.w_dly_sig\[161\]
rlabel metal1 8188 2074 8188 2074 0 tdc0.w_dly_sig\[162\]
rlabel metal1 9200 1802 9200 1802 0 tdc0.w_dly_sig\[163\]
rlabel metal1 9660 1870 9660 1870 0 tdc0.w_dly_sig\[164\]
rlabel metal1 10580 1394 10580 1394 0 tdc0.w_dly_sig\[165\]
rlabel metal1 11822 782 11822 782 0 tdc0.w_dly_sig\[166\]
rlabel metal1 12512 1870 12512 1870 0 tdc0.w_dly_sig\[167\]
rlabel metal1 13110 782 13110 782 0 tdc0.w_dly_sig\[168\]
rlabel metal1 14168 782 14168 782 0 tdc0.w_dly_sig\[169\]
rlabel metal1 28566 7378 28566 7378 0 tdc0.w_dly_sig\[16\]
rlabel metal1 13156 1530 13156 1530 0 tdc0.w_dly_sig\[170\]
rlabel metal1 14490 918 14490 918 0 tdc0.w_dly_sig\[171\]
rlabel metal1 14444 1258 14444 1258 0 tdc0.w_dly_sig\[172\]
rlabel metal1 15594 1938 15594 1938 0 tdc0.w_dly_sig\[173\]
rlabel metal1 16141 2890 16141 2890 0 tdc0.w_dly_sig\[174\]
rlabel metal2 19550 1088 19550 1088 0 tdc0.w_dly_sig\[175\]
rlabel metal1 19826 1428 19826 1428 0 tdc0.w_dly_sig\[176\]
rlabel metal1 20010 1836 20010 1836 0 tdc0.w_dly_sig\[177\]
rlabel metal2 20286 2754 20286 2754 0 tdc0.w_dly_sig\[178\]
rlabel metal2 20470 1598 20470 1598 0 tdc0.w_dly_sig\[179\]
rlabel metal1 28566 6834 28566 6834 0 tdc0.w_dly_sig\[17\]
rlabel metal1 22673 782 22673 782 0 tdc0.w_dly_sig\[180\]
rlabel metal1 22264 1530 22264 1530 0 tdc0.w_dly_sig\[181\]
rlabel metal1 22816 1530 22816 1530 0 tdc0.w_dly_sig\[182\]
rlabel metal1 24288 1870 24288 1870 0 tdc0.w_dly_sig\[183\]
rlabel metal2 24518 2176 24518 2176 0 tdc0.w_dly_sig\[184\]
rlabel metal2 24058 2754 24058 2754 0 tdc0.w_dly_sig\[185\]
rlabel metal1 25622 2346 25622 2346 0 tdc0.w_dly_sig\[186\]
rlabel metal1 25530 2822 25530 2822 0 tdc0.w_dly_sig\[187\]
rlabel metal1 28811 2890 28811 2890 0 tdc0.w_dly_sig\[188\]
rlabel metal1 27784 3706 27784 3706 0 tdc0.w_dly_sig\[189\]
rlabel metal1 29578 6256 29578 6256 0 tdc0.w_dly_sig\[18\]
rlabel metal1 27512 3978 27512 3978 0 tdc0.w_dly_sig\[190\]
rlabel metal1 28980 3706 28980 3706 0 tdc0.w_dly_sig\[191\]
rlabel metal1 30682 4080 30682 4080 0 tdc0.w_dly_sig\[192\]
rlabel metal1 30222 3162 30222 3162 0 tdc0.w_dly_sig\[193\]
rlabel metal1 28934 5746 28934 5746 0 tdc0.w_dly_sig\[19\]
rlabel metal1 25913 11594 25913 11594 0 tdc0.w_dly_sig\[1\]
rlabel metal2 27554 7106 27554 7106 0 tdc0.w_dly_sig\[20\]
rlabel metal1 27416 6222 27416 6222 0 tdc0.w_dly_sig\[21\]
rlabel metal1 26174 6222 26174 6222 0 tdc0.w_dly_sig\[22\]
rlabel metal1 25760 6222 25760 6222 0 tdc0.w_dly_sig\[23\]
rlabel metal1 23920 5746 23920 5746 0 tdc0.w_dly_sig\[24\]
rlabel metal1 24334 6256 24334 6256 0 tdc0.w_dly_sig\[25\]
rlabel metal1 22034 6256 22034 6256 0 tdc0.w_dly_sig\[26\]
rlabel metal1 22586 6732 22586 6732 0 tdc0.w_dly_sig\[27\]
rlabel metal2 21482 7412 21482 7412 0 tdc0.w_dly_sig\[28\]
rlabel metal2 21712 5814 21712 5814 0 tdc0.w_dly_sig\[29\]
rlabel metal1 25668 10030 25668 10030 0 tdc0.w_dly_sig\[2\]
rlabel via1 22130 8330 22130 8330 0 tdc0.w_dly_sig\[30\]
rlabel metal1 22034 8976 22034 8976 0 tdc0.w_dly_sig\[31\]
rlabel metal1 21850 7752 21850 7752 0 tdc0.w_dly_sig\[32\]
rlabel metal1 21390 10608 21390 10608 0 tdc0.w_dly_sig\[33\]
rlabel metal1 22172 9894 22172 9894 0 tdc0.w_dly_sig\[34\]
rlabel metal1 22222 11186 22222 11186 0 tdc0.w_dly_sig\[35\]
rlabel metal1 23690 11696 23690 11696 0 tdc0.w_dly_sig\[36\]
rlabel metal2 24426 13056 24426 13056 0 tdc0.w_dly_sig\[37\]
rlabel metal1 25024 13362 25024 13362 0 tdc0.w_dly_sig\[38\]
rlabel metal1 25116 13158 25116 13158 0 tdc0.w_dly_sig\[39\]
rlabel metal1 25392 11118 25392 11118 0 tdc0.w_dly_sig\[3\]
rlabel metal1 27048 13702 27048 13702 0 tdc0.w_dly_sig\[40\]
rlabel metal1 28014 13804 28014 13804 0 tdc0.w_dly_sig\[41\]
rlabel metal2 26818 14722 26818 14722 0 tdc0.w_dly_sig\[42\]
rlabel metal1 28290 14246 28290 14246 0 tdc0.w_dly_sig\[43\]
rlabel metal1 29302 13702 29302 13702 0 tdc0.w_dly_sig\[44\]
rlabel metal2 29670 14654 29670 14654 0 tdc0.w_dly_sig\[45\]
rlabel metal1 28612 15538 28612 15538 0 tdc0.w_dly_sig\[46\]
rlabel metal1 29164 16218 29164 16218 0 tdc0.w_dly_sig\[47\]
rlabel metal1 27278 16014 27278 16014 0 tdc0.w_dly_sig\[48\]
rlabel metal1 26818 16592 26818 16592 0 tdc0.w_dly_sig\[49\]
rlabel metal1 27922 11220 27922 11220 0 tdc0.w_dly_sig\[4\]
rlabel metal2 25438 16524 25438 16524 0 tdc0.w_dly_sig\[50\]
rlabel via1 27466 17034 27466 17034 0 tdc0.w_dly_sig\[51\]
rlabel metal1 24380 17714 24380 17714 0 tdc0.w_dly_sig\[52\]
rlabel metal1 23372 17782 23372 17782 0 tdc0.w_dly_sig\[53\]
rlabel metal1 23322 18190 23322 18190 0 tdc0.w_dly_sig\[54\]
rlabel metal1 23782 18054 23782 18054 0 tdc0.w_dly_sig\[55\]
rlabel metal1 20838 18836 20838 18836 0 tdc0.w_dly_sig\[56\]
rlabel metal1 17020 18190 17020 18190 0 tdc0.w_dly_sig\[57\]
rlabel metal1 20102 18054 20102 18054 0 tdc0.w_dly_sig\[58\]
rlabel metal1 16642 17714 16642 17714 0 tdc0.w_dly_sig\[59\]
rlabel metal2 27278 11458 27278 11458 0 tdc0.w_dly_sig\[5\]
rlabel metal1 19826 17102 19826 17102 0 tdc0.w_dly_sig\[60\]
rlabel metal2 19274 17102 19274 17102 0 tdc0.w_dly_sig\[61\]
rlabel metal1 20700 17034 20700 17034 0 tdc0.w_dly_sig\[62\]
rlabel metal1 22356 16626 22356 16626 0 tdc0.w_dly_sig\[63\]
rlabel metal1 21988 16422 21988 16422 0 tdc0.w_dly_sig\[64\]
rlabel metal1 20274 16422 20274 16422 0 tdc0.w_dly_sig\[65\]
rlabel metal1 20792 15878 20792 15878 0 tdc0.w_dly_sig\[66\]
rlabel metal2 20930 15181 20930 15181 0 tdc0.w_dly_sig\[67\]
rlabel metal1 15548 15538 15548 15538 0 tdc0.w_dly_sig\[68\]
rlabel metal2 19826 14756 19826 14756 0 tdc0.w_dly_sig\[69\]
rlabel metal1 28750 11696 28750 11696 0 tdc0.w_dly_sig\[6\]
rlabel metal1 16647 14926 16647 14926 0 tdc0.w_dly_sig\[70\]
rlabel metal1 14490 15130 14490 15130 0 tdc0.w_dly_sig\[71\]
rlabel metal2 14214 14688 14214 14688 0 tdc0.w_dly_sig\[72\]
rlabel metal1 12558 14450 12558 14450 0 tdc0.w_dly_sig\[73\]
rlabel metal1 11403 9486 11403 9486 0 tdc0.w_dly_sig\[74\]
rlabel metal1 11776 12342 11776 12342 0 tdc0.w_dly_sig\[75\]
rlabel metal1 12006 10982 12006 10982 0 tdc0.w_dly_sig\[76\]
rlabel metal1 12006 11118 12006 11118 0 tdc0.w_dly_sig\[77\]
rlabel metal2 10258 9384 10258 9384 0 tdc0.w_dly_sig\[78\]
rlabel metal1 9798 11798 9798 11798 0 tdc0.w_dly_sig\[79\]
rlabel metal1 29210 12614 29210 12614 0 tdc0.w_dly_sig\[7\]
rlabel metal2 9200 12750 9200 12750 0 tdc0.w_dly_sig\[80\]
rlabel metal1 9706 13328 9706 13328 0 tdc0.w_dly_sig\[81\]
rlabel metal1 9982 14450 9982 14450 0 tdc0.w_dly_sig\[82\]
rlabel via1 10161 13770 10161 13770 0 tdc0.w_dly_sig\[83\]
rlabel metal1 10437 14858 10437 14858 0 tdc0.w_dly_sig\[84\]
rlabel metal1 9338 15504 9338 15504 0 tdc0.w_dly_sig\[85\]
rlabel metal1 10902 16048 10902 16048 0 tdc0.w_dly_sig\[86\]
rlabel metal1 13202 15504 13202 15504 0 tdc0.w_dly_sig\[87\]
rlabel metal1 11132 16422 11132 16422 0 tdc0.w_dly_sig\[88\]
rlabel metal1 12934 17170 12934 17170 0 tdc0.w_dly_sig\[89\]
rlabel metal1 30548 11594 30548 11594 0 tdc0.w_dly_sig\[8\]
rlabel metal1 13186 16694 13186 16694 0 tdc0.w_dly_sig\[90\]
rlabel metal1 13830 17782 13830 17782 0 tdc0.w_dly_sig\[91\]
rlabel metal2 14214 18598 14214 18598 0 tdc0.w_dly_sig\[92\]
rlabel metal1 9614 18292 9614 18292 0 tdc0.w_dly_sig\[93\]
rlabel metal1 9982 18734 9982 18734 0 tdc0.w_dly_sig\[94\]
rlabel metal1 8280 18802 8280 18802 0 tdc0.w_dly_sig\[95\]
rlabel metal2 9246 17544 9246 17544 0 tdc0.w_dly_sig\[96\]
rlabel via1 8586 17782 8586 17782 0 tdc0.w_dly_sig\[97\]
rlabel metal2 7958 17068 7958 17068 0 tdc0.w_dly_sig\[98\]
rlabel metal1 6624 17306 6624 17306 0 tdc0.w_dly_sig\[99\]
rlabel via1 30686 11186 30686 11186 0 tdc0.w_dly_sig\[9\]
rlabel metal1 25898 10540 25898 10540 0 tdc0.w_dly_sig_n\[0\]
rlabel metal1 6118 16626 6118 16626 0 tdc0.w_dly_sig_n\[100\]
rlabel metal1 4094 16626 4094 16626 0 tdc0.w_dly_sig_n\[101\]
rlabel metal1 3496 16422 3496 16422 0 tdc0.w_dly_sig_n\[102\]
rlabel metal1 2346 16014 2346 16014 0 tdc0.w_dly_sig_n\[103\]
rlabel metal1 1932 16218 1932 16218 0 tdc0.w_dly_sig_n\[104\]
rlabel metal1 1380 15334 1380 15334 0 tdc0.w_dly_sig_n\[105\]
rlabel metal1 1886 15130 1886 15130 0 tdc0.w_dly_sig_n\[106\]
rlabel metal1 2300 14314 2300 14314 0 tdc0.w_dly_sig_n\[107\]
rlabel metal1 1426 13872 1426 13872 0 tdc0.w_dly_sig_n\[108\]
rlabel metal1 1242 12750 1242 12750 0 tdc0.w_dly_sig_n\[109\]
rlabel metal1 30406 9520 30406 9520 0 tdc0.w_dly_sig_n\[10\]
rlabel metal1 1472 11662 1472 11662 0 tdc0.w_dly_sig_n\[110\]
rlabel metal1 2024 10438 2024 10438 0 tdc0.w_dly_sig_n\[111\]
rlabel metal1 1334 9486 1334 9486 0 tdc0.w_dly_sig_n\[112\]
rlabel metal1 2300 9350 2300 9350 0 tdc0.w_dly_sig_n\[113\]
rlabel metal1 1380 8942 1380 8942 0 tdc0.w_dly_sig_n\[114\]
rlabel metal1 2438 9010 2438 9010 0 tdc0.w_dly_sig_n\[115\]
rlabel metal1 3450 8976 3450 8976 0 tdc0.w_dly_sig_n\[116\]
rlabel metal1 3358 9350 3358 9350 0 tdc0.w_dly_sig_n\[117\]
rlabel metal1 3634 10098 3634 10098 0 tdc0.w_dly_sig_n\[118\]
rlabel metal1 4232 10098 4232 10098 0 tdc0.w_dly_sig_n\[119\]
rlabel metal1 29164 8806 29164 8806 0 tdc0.w_dly_sig_n\[11\]
rlabel metal1 4646 12784 4646 12784 0 tdc0.w_dly_sig_n\[120\]
rlabel metal1 4278 13158 4278 13158 0 tdc0.w_dly_sig_n\[121\]
rlabel metal1 4554 13770 4554 13770 0 tdc0.w_dly_sig_n\[122\]
rlabel metal1 5060 13838 5060 13838 0 tdc0.w_dly_sig_n\[123\]
rlabel metal1 6072 14450 6072 14450 0 tdc0.w_dly_sig_n\[124\]
rlabel metal1 7314 14042 7314 14042 0 tdc0.w_dly_sig_n\[125\]
rlabel metal1 7590 13838 7590 13838 0 tdc0.w_dly_sig_n\[126\]
rlabel metal1 7172 12272 7172 12272 0 tdc0.w_dly_sig_n\[127\]
rlabel metal1 7452 9894 7452 9894 0 tdc0.w_dly_sig_n\[128\]
rlabel metal1 7176 9350 7176 9350 0 tdc0.w_dly_sig_n\[129\]
rlabel metal1 28934 8602 28934 8602 0 tdc0.w_dly_sig_n\[12\]
rlabel metal1 7038 9078 7038 9078 0 tdc0.w_dly_sig_n\[130\]
rlabel metal1 7084 8602 7084 8602 0 tdc0.w_dly_sig_n\[131\]
rlabel metal1 6486 8398 6486 8398 0 tdc0.w_dly_sig_n\[132\]
rlabel metal1 6716 7718 6716 7718 0 tdc0.w_dly_sig_n\[133\]
rlabel metal1 5934 7310 5934 7310 0 tdc0.w_dly_sig_n\[134\]
rlabel metal1 6072 6698 6072 6698 0 tdc0.w_dly_sig_n\[135\]
rlabel metal2 8694 7072 8694 7072 0 tdc0.w_dly_sig_n\[136\]
rlabel metal2 8510 6528 8510 6528 0 tdc0.w_dly_sig_n\[137\]
rlabel metal1 9522 6188 9522 6188 0 tdc0.w_dly_sig_n\[138\]
rlabel metal1 10488 6222 10488 6222 0 tdc0.w_dly_sig_n\[139\]
rlabel metal1 29348 8330 29348 8330 0 tdc0.w_dly_sig_n\[13\]
rlabel metal1 9844 5338 9844 5338 0 tdc0.w_dly_sig_n\[140\]
rlabel metal1 9246 5168 9246 5168 0 tdc0.w_dly_sig_n\[141\]
rlabel metal1 8050 5134 8050 5134 0 tdc0.w_dly_sig_n\[142\]
rlabel metal1 7590 5542 7590 5542 0 tdc0.w_dly_sig_n\[143\]
rlabel metal1 5842 5134 5842 5134 0 tdc0.w_dly_sig_n\[144\]
rlabel metal1 4922 5338 4922 5338 0 tdc0.w_dly_sig_n\[145\]
rlabel metal1 4278 5134 4278 5134 0 tdc0.w_dly_sig_n\[146\]
rlabel metal1 3818 6086 3818 6086 0 tdc0.w_dly_sig_n\[147\]
rlabel metal2 2622 6052 2622 6052 0 tdc0.w_dly_sig_n\[148\]
rlabel metal1 2346 5202 2346 5202 0 tdc0.w_dly_sig_n\[149\]
rlabel metal1 30452 6834 30452 6834 0 tdc0.w_dly_sig_n\[14\]
rlabel metal1 1610 5134 1610 5134 0 tdc0.w_dly_sig_n\[150\]
rlabel metal1 1150 4658 1150 4658 0 tdc0.w_dly_sig_n\[151\]
rlabel metal1 2484 3910 2484 3910 0 tdc0.w_dly_sig_n\[152\]
rlabel metal1 1518 3570 1518 3570 0 tdc0.w_dly_sig_n\[153\]
rlabel metal1 1932 2890 1932 2890 0 tdc0.w_dly_sig_n\[154\]
rlabel metal1 2530 2516 2530 2516 0 tdc0.w_dly_sig_n\[155\]
rlabel metal1 3174 2448 3174 2448 0 tdc0.w_dly_sig_n\[156\]
rlabel metal1 3956 2414 3956 2414 0 tdc0.w_dly_sig_n\[157\]
rlabel via1 5194 1870 5194 1870 0 tdc0.w_dly_sig_n\[158\]
rlabel metal1 5704 1802 5704 1802 0 tdc0.w_dly_sig_n\[159\]
rlabel metal1 30866 7514 30866 7514 0 tdc0.w_dly_sig_n\[15\]
rlabel metal1 6808 1802 6808 1802 0 tdc0.w_dly_sig_n\[160\]
rlabel metal1 7360 1530 7360 1530 0 tdc0.w_dly_sig_n\[161\]
rlabel metal1 8326 1394 8326 1394 0 tdc0.w_dly_sig_n\[162\]
rlabel metal1 8050 1394 8050 1394 0 tdc0.w_dly_sig_n\[163\]
rlabel metal1 9246 1428 9246 1428 0 tdc0.w_dly_sig_n\[164\]
rlabel metal2 9706 1564 9706 1564 0 tdc0.w_dly_sig_n\[165\]
rlabel metal1 10856 1462 10856 1462 0 tdc0.w_dly_sig_n\[166\]
rlabel metal2 12374 1258 12374 1258 0 tdc0.w_dly_sig_n\[167\]
rlabel metal1 12696 1394 12696 1394 0 tdc0.w_dly_sig_n\[168\]
rlabel metal1 14030 1360 14030 1360 0 tdc0.w_dly_sig_n\[169\]
rlabel metal1 30544 5134 30544 5134 0 tdc0.w_dly_sig_n\[16\]
rlabel metal1 14444 1394 14444 1394 0 tdc0.w_dly_sig_n\[170\]
rlabel metal1 15226 1428 15226 1428 0 tdc0.w_dly_sig_n\[171\]
rlabel via1 15686 1870 15686 1870 0 tdc0.w_dly_sig_n\[172\]
rlabel metal1 16652 1734 16652 1734 0 tdc0.w_dly_sig_n\[173\]
rlabel metal1 17710 1870 17710 1870 0 tdc0.w_dly_sig_n\[174\]
rlabel metal2 18814 1632 18814 1632 0 tdc0.w_dly_sig_n\[175\]
rlabel metal1 19780 1258 19780 1258 0 tdc0.w_dly_sig_n\[176\]
rlabel metal1 20148 2074 20148 2074 0 tdc0.w_dly_sig_n\[177\]
rlabel metal1 21206 1190 21206 1190 0 tdc0.w_dly_sig_n\[178\]
rlabel metal1 22172 1326 22172 1326 0 tdc0.w_dly_sig_n\[179\]
rlabel metal2 28750 6086 28750 6086 0 tdc0.w_dly_sig_n\[17\]
rlabel metal1 22172 1190 22172 1190 0 tdc0.w_dly_sig_n\[180\]
rlabel metal1 23322 1394 23322 1394 0 tdc0.w_dly_sig_n\[181\]
rlabel metal1 24610 1904 24610 1904 0 tdc0.w_dly_sig_n\[182\]
rlabel metal1 24104 2074 24104 2074 0 tdc0.w_dly_sig_n\[183\]
rlabel metal1 25530 2278 25530 2278 0 tdc0.w_dly_sig_n\[184\]
rlabel metal1 25852 2822 25852 2822 0 tdc0.w_dly_sig_n\[185\]
rlabel metal1 26588 2890 26588 2890 0 tdc0.w_dly_sig_n\[186\]
rlabel metal1 27232 3094 27232 3094 0 tdc0.w_dly_sig_n\[187\]
rlabel metal2 27186 3094 27186 3094 0 tdc0.w_dly_sig_n\[188\]
rlabel metal1 28658 3570 28658 3570 0 tdc0.w_dly_sig_n\[189\]
rlabel metal1 29762 6698 29762 6698 0 tdc0.w_dly_sig_n\[18\]
rlabel metal1 28842 3978 28842 3978 0 tdc0.w_dly_sig_n\[190\]
rlabel metal2 29670 3808 29670 3808 0 tdc0.w_dly_sig_n\[191\]
rlabel metal1 29348 4590 29348 4590 0 tdc0.w_dly_sig_n\[192\]
rlabel metal1 28244 5882 28244 5882 0 tdc0.w_dly_sig_n\[19\]
rlabel metal1 25392 10778 25392 10778 0 tdc0.w_dly_sig_n\[1\]
rlabel metal1 26634 5780 26634 5780 0 tdc0.w_dly_sig_n\[20\]
rlabel metal1 27416 6154 27416 6154 0 tdc0.w_dly_sig_n\[21\]
rlabel metal1 25898 5882 25898 5882 0 tdc0.w_dly_sig_n\[22\]
rlabel metal1 24610 5780 24610 5780 0 tdc0.w_dly_sig_n\[23\]
rlabel metal1 24518 6154 24518 6154 0 tdc0.w_dly_sig_n\[24\]
rlabel metal1 23874 6426 23874 6426 0 tdc0.w_dly_sig_n\[25\]
rlabel metal1 22632 6426 22632 6426 0 tdc0.w_dly_sig_n\[26\]
rlabel metal1 22034 6800 22034 6800 0 tdc0.w_dly_sig_n\[27\]
rlabel metal1 21252 7174 21252 7174 0 tdc0.w_dly_sig_n\[28\]
rlabel metal1 22264 7922 22264 7922 0 tdc0.w_dly_sig_n\[29\]
rlabel metal1 26864 10506 26864 10506 0 tdc0.w_dly_sig_n\[2\]
rlabel metal1 21896 7514 21896 7514 0 tdc0.w_dly_sig_n\[30\]
rlabel metal1 22011 9486 22011 9486 0 tdc0.w_dly_sig_n\[31\]
rlabel metal2 21666 9894 21666 9894 0 tdc0.w_dly_sig_n\[32\]
rlabel metal1 21896 10098 21896 10098 0 tdc0.w_dly_sig_n\[33\]
rlabel metal1 22816 10098 22816 10098 0 tdc0.w_dly_sig_n\[34\]
rlabel metal1 22356 11662 22356 11662 0 tdc0.w_dly_sig_n\[35\]
rlabel metal1 22954 11798 22954 11798 0 tdc0.w_dly_sig_n\[36\]
rlabel metal1 24334 12682 24334 12682 0 tdc0.w_dly_sig_n\[37\]
rlabel metal1 25668 13498 25668 13498 0 tdc0.w_dly_sig_n\[38\]
rlabel metal1 26312 13838 26312 13838 0 tdc0.w_dly_sig_n\[39\]
rlabel metal1 27186 11152 27186 11152 0 tdc0.w_dly_sig_n\[3\]
rlabel metal1 26726 14450 26726 14450 0 tdc0.w_dly_sig_n\[40\]
rlabel metal1 27922 14416 27922 14416 0 tdc0.w_dly_sig_n\[41\]
rlabel metal1 28014 14518 28014 14518 0 tdc0.w_dly_sig_n\[42\]
rlabel metal1 29302 14586 29302 14586 0 tdc0.w_dly_sig_n\[43\]
rlabel metal2 29394 14416 29394 14416 0 tdc0.w_dly_sig_n\[44\]
rlabel metal1 29486 15130 29486 15130 0 tdc0.w_dly_sig_n\[45\]
rlabel metal1 28520 15470 28520 15470 0 tdc0.w_dly_sig_n\[46\]
rlabel metal2 28474 15776 28474 15776 0 tdc0.w_dly_sig_n\[47\]
rlabel metal1 28428 16626 28428 16626 0 tdc0.w_dly_sig_n\[48\]
rlabel metal2 26910 16320 26910 16320 0 tdc0.w_dly_sig_n\[49\]
rlabel metal1 27692 11050 27692 11050 0 tdc0.w_dly_sig_n\[4\]
rlabel metal1 25714 17136 25714 17136 0 tdc0.w_dly_sig_n\[50\]
rlabel metal2 25346 17510 25346 17510 0 tdc0.w_dly_sig_n\[51\]
rlabel metal1 25254 17850 25254 17850 0 tdc0.w_dly_sig_n\[52\]
rlabel metal1 24242 18190 24242 18190 0 tdc0.w_dly_sig_n\[53\]
rlabel metal2 22770 18496 22770 18496 0 tdc0.w_dly_sig_n\[54\]
rlabel metal1 22816 18122 22816 18122 0 tdc0.w_dly_sig_n\[55\]
rlabel metal1 21114 18802 21114 18802 0 tdc0.w_dly_sig_n\[56\]
rlabel metal1 19964 18122 19964 18122 0 tdc0.w_dly_sig_n\[57\]
rlabel metal2 16974 17884 16974 17884 0 tdc0.w_dly_sig_n\[58\]
rlabel metal1 18860 17646 18860 17646 0 tdc0.w_dly_sig_n\[59\]
rlabel metal1 29026 11186 29026 11186 0 tdc0.w_dly_sig_n\[5\]
rlabel metal1 19504 17306 19504 17306 0 tdc0.w_dly_sig_n\[60\]
rlabel metal1 20010 17238 20010 17238 0 tdc0.w_dly_sig_n\[61\]
rlabel metal1 21206 16626 21206 16626 0 tdc0.w_dly_sig_n\[62\]
rlabel metal1 21666 16626 21666 16626 0 tdc0.w_dly_sig_n\[63\]
rlabel viali 20842 16014 20842 16014 0 tdc0.w_dly_sig_n\[64\]
rlabel metal1 21344 15878 21344 15878 0 tdc0.w_dly_sig_n\[65\]
rlabel metal1 18630 16014 18630 16014 0 tdc0.w_dly_sig_n\[66\]
rlabel metal2 19090 15776 19090 15776 0 tdc0.w_dly_sig_n\[67\]
rlabel metal1 17480 15470 17480 15470 0 tdc0.w_dly_sig_n\[68\]
rlabel metal1 15456 14926 15456 14926 0 tdc0.w_dly_sig_n\[69\]
rlabel metal1 29762 12614 29762 12614 0 tdc0.w_dly_sig_n\[6\]
rlabel metal1 15502 15130 15502 15130 0 tdc0.w_dly_sig_n\[70\]
rlabel metal1 14628 14450 14628 14450 0 tdc0.w_dly_sig_n\[71\]
rlabel metal1 13754 14382 13754 14382 0 tdc0.w_dly_sig_n\[72\]
rlabel metal1 13064 14314 13064 14314 0 tdc0.w_dly_sig_n\[73\]
rlabel metal2 12282 12512 12282 12512 0 tdc0.w_dly_sig_n\[74\]
rlabel metal1 12512 11118 12512 11118 0 tdc0.w_dly_sig_n\[75\]
rlabel metal1 11362 11186 11362 11186 0 tdc0.w_dly_sig_n\[76\]
rlabel metal1 10350 10608 10350 10608 0 tdc0.w_dly_sig_n\[77\]
rlabel metal1 9752 11050 9752 11050 0 tdc0.w_dly_sig_n\[78\]
rlabel metal1 9660 11866 9660 11866 0 tdc0.w_dly_sig_n\[79\]
rlabel metal1 29072 11526 29072 11526 0 tdc0.w_dly_sig_n\[7\]
rlabel metal2 9706 12580 9706 12580 0 tdc0.w_dly_sig_n\[80\]
rlabel metal1 9476 13158 9476 13158 0 tdc0.w_dly_sig_n\[81\]
rlabel metal1 9844 14314 9844 14314 0 tdc0.w_dly_sig_n\[82\]
rlabel metal1 9660 14790 9660 14790 0 tdc0.w_dly_sig_n\[83\]
rlabel metal1 9568 15538 9568 15538 0 tdc0.w_dly_sig_n\[84\]
rlabel metal1 9890 16048 9890 16048 0 tdc0.w_dly_sig_n\[85\]
rlabel metal1 10902 15946 10902 15946 0 tdc0.w_dly_sig_n\[86\]
rlabel metal2 11454 16320 11454 16320 0 tdc0.w_dly_sig_n\[87\]
rlabel metal2 12466 16932 12466 16932 0 tdc0.w_dly_sig_n\[88\]
rlabel metal1 12834 17068 12834 17068 0 tdc0.w_dly_sig_n\[89\]
rlabel metal1 29578 10574 29578 10574 0 tdc0.w_dly_sig_n\[8\]
rlabel metal1 13064 17850 13064 17850 0 tdc0.w_dly_sig_n\[90\]
rlabel metal1 13524 18054 13524 18054 0 tdc0.w_dly_sig_n\[91\]
rlabel metal1 11822 18190 11822 18190 0 tdc0.w_dly_sig_n\[92\]
rlabel metal1 10028 18598 10028 18598 0 tdc0.w_dly_sig_n\[93\]
rlabel metal1 9798 18802 9798 18802 0 tdc0.w_dly_sig_n\[94\]
rlabel metal1 8556 18190 8556 18190 0 tdc0.w_dly_sig_n\[95\]
rlabel metal1 7728 18258 7728 18258 0 tdc0.w_dly_sig_n\[96\]
rlabel metal1 7084 17850 7084 17850 0 tdc0.w_dly_sig_n\[97\]
rlabel metal1 7176 17306 7176 17306 0 tdc0.w_dly_sig_n\[98\]
rlabel metal1 6164 17034 6164 17034 0 tdc0.w_dly_sig_n\[99\]
rlabel metal1 28842 10166 28842 10166 0 tdc0.w_dly_sig_n\[9\]
rlabel metal1 31326 10574 31326 10574 0 ui_in[0]
rlabel metal2 15502 415 15502 415 0 ui_in[3]
rlabel via1 16146 364 16146 364 0 ui_in[4]
rlabel metal2 16790 534 16790 534 0 ui_in[5]
rlabel metal2 17434 874 17434 874 0 ui_in[6]
rlabel metal2 18078 874 18078 874 0 ui_in[7]
rlabel metal2 20332 13260 20332 13260 0 uo_out[0]
rlabel metal3 28712 9588 28712 9588 0 uo_out[1]
rlabel metal2 18768 12852 18768 12852 0 uo_out[2]
rlabel metal1 18814 13804 18814 13804 0 uo_out[3]
rlabel metal2 19090 12716 19090 12716 0 uo_out[4]
rlabel metal3 30184 12308 30184 12308 0 uo_out[5]
rlabel metal1 20332 12206 20332 12206 0 uo_out[6]
rlabel metal1 21068 12818 21068 12818 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 32000 20000
<< end >>
