magic
tech sky130A
magscale 1 2
timestamp 1710401781
<< viali >>
rect 13185 18921 13219 18955
rect 14197 18921 14231 18955
rect 12909 18853 12943 18887
rect 1409 18785 1443 18819
rect 11437 18785 11471 18819
rect 11529 18785 11563 18819
rect 12081 18785 12115 18819
rect 12541 18785 12575 18819
rect 13001 18785 13035 18819
rect 13093 18785 13127 18819
rect 13737 18785 13771 18819
rect 13829 18785 13863 18819
rect 14105 18785 14139 18819
rect 14381 18785 14415 18819
rect 18521 18785 18555 18819
rect 1133 18717 1167 18751
rect 857 18581 891 18615
rect 12173 18581 12207 18615
rect 12633 18581 12667 18615
rect 13645 18581 13679 18615
rect 13921 18581 13955 18615
rect 14473 18581 14507 18615
rect 19073 18581 19107 18615
rect 10425 18377 10459 18411
rect 11989 18377 12023 18411
rect 12541 18377 12575 18411
rect 11713 18309 11747 18343
rect 3249 18241 3283 18275
rect 11069 18241 11103 18275
rect 857 18173 891 18207
rect 2697 18173 2731 18207
rect 3065 18173 3099 18207
rect 4721 18173 4755 18207
rect 4988 18173 5022 18207
rect 7573 18173 7607 18207
rect 8861 18173 8895 18207
rect 9128 18173 9162 18207
rect 10333 18173 10367 18207
rect 10977 18173 11011 18207
rect 11345 18173 11379 18207
rect 11805 18173 11839 18207
rect 12081 18173 12115 18207
rect 12357 18173 12391 18207
rect 12449 18173 12483 18207
rect 12725 18173 12759 18207
rect 13001 18173 13035 18207
rect 15117 18173 15151 18207
rect 15209 18173 15243 18207
rect 15476 18173 15510 18207
rect 18061 18173 18095 18207
rect 19073 18173 19107 18207
rect 3516 18105 3550 18139
rect 7328 18105 7362 18139
rect 11437 18105 11471 18139
rect 12265 18105 12299 18139
rect 14861 18105 14895 18139
rect 17816 18105 17850 18139
rect 2605 18037 2639 18071
rect 2973 18037 3007 18071
rect 4629 18037 4663 18071
rect 6101 18037 6135 18071
rect 6193 18037 6227 18071
rect 10241 18037 10275 18071
rect 12817 18037 12851 18071
rect 13093 18037 13127 18071
rect 13737 18037 13771 18071
rect 16589 18037 16623 18071
rect 16681 18037 16715 18071
rect 14381 17833 14415 17867
rect 2666 17765 2700 17799
rect 6469 17765 6503 17799
rect 10057 17765 10091 17799
rect 16497 17765 16531 17799
rect 2053 17697 2087 17731
rect 2329 17697 2363 17731
rect 4077 17697 4111 17731
rect 4169 17697 4203 17731
rect 4436 17697 4470 17731
rect 6193 17697 6227 17731
rect 6377 17697 6411 17731
rect 6561 17697 6595 17731
rect 7961 17697 7995 17731
rect 8217 17697 8251 17731
rect 8309 17697 8343 17731
rect 8576 17697 8610 17731
rect 9965 17697 9999 17731
rect 10149 17697 10183 17731
rect 10333 17697 10367 17731
rect 10793 17697 10827 17731
rect 10977 17697 11011 17731
rect 11161 17697 11195 17731
rect 11253 17697 11287 17731
rect 11345 17697 11379 17731
rect 11621 17697 11655 17731
rect 13010 17697 13044 17731
rect 13369 17697 13403 17731
rect 13461 17697 13495 17731
rect 13737 17697 13771 17731
rect 14013 17697 14047 17731
rect 14289 17697 14323 17731
rect 14821 17697 14855 17731
rect 16313 17697 16347 17731
rect 16405 17697 16439 17731
rect 16681 17697 16715 17731
rect 17049 17697 17083 17731
rect 18265 17697 18299 17731
rect 18521 17697 18555 17731
rect 18613 17697 18647 17731
rect 2421 17629 2455 17663
rect 13277 17629 13311 17663
rect 14565 17629 14599 17663
rect 3801 17561 3835 17595
rect 5549 17561 5583 17595
rect 11713 17561 11747 17595
rect 14105 17561 14139 17595
rect 1961 17493 1995 17527
rect 2237 17493 2271 17527
rect 3985 17493 4019 17527
rect 6745 17493 6779 17527
rect 6837 17493 6871 17527
rect 9689 17493 9723 17527
rect 9781 17493 9815 17527
rect 10701 17493 10735 17527
rect 11529 17493 11563 17527
rect 11897 17493 11931 17527
rect 13829 17493 13863 17527
rect 15945 17493 15979 17527
rect 16129 17493 16163 17527
rect 16957 17493 16991 17527
rect 17141 17493 17175 17527
rect 18705 17493 18739 17527
rect 1409 17289 1443 17323
rect 2973 17289 3007 17323
rect 4629 17289 4663 17323
rect 4905 17289 4939 17323
rect 8493 17289 8527 17323
rect 9413 17289 9447 17323
rect 9597 17289 9631 17323
rect 11437 17289 11471 17323
rect 11713 17289 11747 17323
rect 11989 17289 12023 17323
rect 13645 17289 13679 17323
rect 15485 17289 15519 17323
rect 16589 17289 16623 17323
rect 16865 17289 16899 17323
rect 18797 17289 18831 17323
rect 13277 17221 13311 17255
rect 17417 17221 17451 17255
rect 1593 17153 1627 17187
rect 5549 17153 5583 17187
rect 15209 17153 15243 17187
rect 17693 17153 17727 17187
rect 857 17085 891 17119
rect 1501 17085 1535 17119
rect 1860 17085 1894 17119
rect 3525 17085 3559 17119
rect 3801 17085 3835 17119
rect 4077 17085 4111 17119
rect 4353 17085 4387 17119
rect 4721 17085 4755 17119
rect 4813 17085 4847 17119
rect 7573 17085 7607 17119
rect 7849 17085 7883 17119
rect 7941 17085 7975 17119
rect 8585 17085 8619 17119
rect 9229 17085 9263 17119
rect 9689 17085 9723 17119
rect 10701 17085 10735 17119
rect 10793 17085 10827 17119
rect 11161 17085 11195 17119
rect 11253 17085 11287 17119
rect 11529 17085 11563 17119
rect 11805 17085 11839 17119
rect 11897 17085 11931 17119
rect 13369 17085 13403 17119
rect 13737 17085 13771 17119
rect 14197 17085 14231 17119
rect 14289 17085 14323 17119
rect 14749 17085 14783 17119
rect 14841 17085 14875 17119
rect 15301 17085 15335 17119
rect 15393 17085 15427 17119
rect 16681 17085 16715 17119
rect 16773 17085 16807 17119
rect 17049 17085 17083 17119
rect 17509 17085 17543 17119
rect 17785 17085 17819 17119
rect 18061 17085 18095 17119
rect 18153 17085 18187 17119
rect 18705 17087 18739 17121
rect 3433 17017 3467 17051
rect 5794 17017 5828 17051
rect 7757 17017 7791 17051
rect 17141 17017 17175 17051
rect 3709 16949 3743 16983
rect 3985 16949 4019 16983
rect 4261 16949 4295 16983
rect 6929 16949 6963 16983
rect 8125 16949 8159 16983
rect 14105 16949 14139 16983
rect 14381 16949 14415 16983
rect 14657 16949 14691 16983
rect 14933 16949 14967 16983
rect 17969 16949 18003 16983
rect 18245 16949 18279 16983
rect 1317 16745 1351 16779
rect 2421 16745 2455 16779
rect 2973 16745 3007 16779
rect 3249 16745 3283 16779
rect 4077 16745 4111 16779
rect 4629 16745 4663 16779
rect 5549 16745 5583 16779
rect 9505 16745 9539 16779
rect 11069 16745 11103 16779
rect 11621 16745 11655 16779
rect 11897 16745 11931 16779
rect 15485 16745 15519 16779
rect 15761 16745 15795 16779
rect 16681 16745 16715 16779
rect 16957 16745 16991 16779
rect 4905 16677 4939 16711
rect 5273 16677 5307 16711
rect 6377 16677 6411 16711
rect 15209 16677 15243 16711
rect 1409 16609 1443 16643
rect 1593 16609 1627 16643
rect 1685 16609 1719 16643
rect 1961 16609 1995 16643
rect 2053 16609 2087 16643
rect 2513 16609 2547 16643
rect 2697 16609 2731 16643
rect 2789 16609 2823 16643
rect 3065 16609 3099 16643
rect 3157 16609 3191 16643
rect 3709 16609 3743 16643
rect 4169 16609 4203 16643
rect 4261 16609 4295 16643
rect 4721 16609 4755 16643
rect 4997 16609 5031 16643
rect 5365 16609 5399 16643
rect 5641 16609 5675 16643
rect 6017 16609 6051 16643
rect 6121 16609 6155 16643
rect 6285 16609 6319 16643
rect 6469 16609 6503 16643
rect 6929 16609 6963 16643
rect 8125 16609 8159 16643
rect 8381 16609 8415 16643
rect 11161 16609 11195 16643
rect 11437 16609 11471 16643
rect 11529 16609 11563 16643
rect 11989 16609 12023 16643
rect 14105 16609 14139 16643
rect 14473 16609 14507 16643
rect 14749 16609 14783 16643
rect 15025 16609 15059 16643
rect 15117 16609 15151 16643
rect 15393 16609 15427 16643
rect 15669 16609 15703 16643
rect 16773 16609 16807 16643
rect 17049 16609 17083 16643
rect 18254 16609 18288 16643
rect 18521 16609 18555 16643
rect 18613 16609 18647 16643
rect 19073 16609 19107 16643
rect 5917 16541 5951 16575
rect 4353 16473 4387 16507
rect 11345 16473 11379 16507
rect 1869 16405 1903 16439
rect 2145 16405 2179 16439
rect 3617 16405 3651 16439
rect 6653 16405 6687 16439
rect 6837 16405 6871 16439
rect 14013 16405 14047 16439
rect 14381 16405 14415 16439
rect 14657 16405 14691 16439
rect 14933 16405 14967 16439
rect 17141 16405 17175 16439
rect 18705 16405 18739 16439
rect 5365 16201 5399 16235
rect 5641 16201 5675 16235
rect 6193 16201 6227 16235
rect 8033 16201 8067 16235
rect 14105 16201 14139 16235
rect 17601 16201 17635 16235
rect 17877 16201 17911 16235
rect 2605 16133 2639 16167
rect 9781 16133 9815 16167
rect 10701 16133 10735 16167
rect 14289 16133 14323 16167
rect 18429 16133 18463 16167
rect 5917 16065 5951 16099
rect 15669 16065 15703 16099
rect 1409 15997 1443 16031
rect 1869 15997 1903 16031
rect 1961 15997 1995 16031
rect 2421 15997 2455 16031
rect 2697 15997 2731 16031
rect 3249 15997 3283 16031
rect 5457 15997 5491 16031
rect 5733 15997 5767 16031
rect 5825 15997 5859 16031
rect 6285 15997 6319 16031
rect 6469 15997 6503 16031
rect 8125 15997 8159 16031
rect 8401 15997 8435 16031
rect 10149 15997 10183 16031
rect 10541 15997 10575 16031
rect 10793 15997 10827 16031
rect 11161 15997 11195 16031
rect 11529 15997 11563 16031
rect 13369 15997 13403 16031
rect 13921 15997 13955 16031
rect 14013 15997 14047 16031
rect 17693 15997 17727 16031
rect 17969 15997 18003 16031
rect 18061 15997 18095 16031
rect 18337 15997 18371 16031
rect 1501 15929 1535 15963
rect 3341 15929 3375 15963
rect 6736 15929 6770 15963
rect 8646 15929 8680 15963
rect 10333 15929 10367 15963
rect 10425 15929 10459 15963
rect 10977 15929 11011 15963
rect 11069 15929 11103 15963
rect 13277 15929 13311 15963
rect 15402 15929 15436 15963
rect 1777 15861 1811 15895
rect 2053 15861 2087 15895
rect 2329 15861 2363 15895
rect 7849 15861 7883 15895
rect 11345 15861 11379 15895
rect 11621 15861 11655 15895
rect 13829 15861 13863 15895
rect 18153 15861 18187 15895
rect 2789 15657 2823 15691
rect 5549 15657 5583 15691
rect 7021 15657 7055 15691
rect 7573 15657 7607 15691
rect 11069 15657 11103 15691
rect 12081 15657 12115 15691
rect 12357 15657 12391 15691
rect 13461 15657 13495 15691
rect 17325 15657 17359 15691
rect 17601 15657 17635 15691
rect 18613 15657 18647 15691
rect 11437 15589 11471 15623
rect 11529 15589 11563 15623
rect 12633 15589 12667 15623
rect 12909 15589 12943 15623
rect 14832 15589 14866 15623
rect 18981 15589 19015 15623
rect 1501 15521 1535 15555
rect 1777 15521 1811 15555
rect 2053 15521 2087 15555
rect 2145 15521 2179 15555
rect 2421 15521 2455 15555
rect 2881 15521 2915 15555
rect 3525 15521 3559 15555
rect 3781 15521 3815 15555
rect 5365 15521 5399 15555
rect 5641 15521 5675 15555
rect 6193 15521 6227 15555
rect 6469 15521 6503 15555
rect 6653 15521 6687 15555
rect 6745 15521 6779 15555
rect 6929 15521 6963 15555
rect 7389 15521 7423 15555
rect 7665 15521 7699 15555
rect 11161 15521 11195 15555
rect 11253 15521 11287 15555
rect 11621 15521 11655 15555
rect 12173 15521 12207 15555
rect 12265 15521 12299 15555
rect 12725 15521 12759 15555
rect 13001 15521 13035 15555
rect 13093 15521 13127 15555
rect 13553 15521 13587 15555
rect 13829 15521 13863 15555
rect 14105 15521 14139 15555
rect 14197 15521 14231 15555
rect 14565 15521 14599 15555
rect 17417 15521 17451 15555
rect 17693 15521 17727 15555
rect 17969 15521 18003 15555
rect 18429 15521 18463 15555
rect 18705 15521 18739 15555
rect 18889 15521 18923 15555
rect 1409 15453 1443 15487
rect 6377 15453 6411 15487
rect 14013 15453 14047 15487
rect 1961 15385 1995 15419
rect 2513 15385 2547 15419
rect 6101 15385 6135 15419
rect 7297 15385 7331 15419
rect 1685 15317 1719 15351
rect 2237 15317 2271 15351
rect 4905 15317 4939 15351
rect 5273 15317 5307 15351
rect 11805 15317 11839 15351
rect 13185 15317 13219 15351
rect 13737 15317 13771 15351
rect 14289 15317 14323 15351
rect 15945 15317 15979 15351
rect 17877 15317 17911 15351
rect 18337 15317 18371 15351
rect 6653 15113 6687 15147
rect 6929 15113 6963 15147
rect 7757 15113 7791 15147
rect 12541 15113 12575 15147
rect 18429 15113 18463 15147
rect 18981 15113 19015 15147
rect 2605 15045 2639 15079
rect 9137 15045 9171 15079
rect 13093 15045 13127 15079
rect 1225 14909 1259 14943
rect 1492 14909 1526 14943
rect 2697 14909 2731 14943
rect 3249 14909 3283 14943
rect 5089 14909 5123 14943
rect 6745 14909 6779 14943
rect 7021 14909 7055 14943
rect 7113 14909 7147 14943
rect 7481 14909 7515 14943
rect 7573 14909 7607 14943
rect 7849 14909 7883 14943
rect 8125 14909 8159 14943
rect 8677 14909 8711 14943
rect 8953 14909 8987 14943
rect 9229 14909 9263 14943
rect 9505 14911 9539 14945
rect 9689 14909 9723 14943
rect 9781 14909 9815 14943
rect 11078 14909 11112 14943
rect 11345 14909 11379 14943
rect 11713 14909 11747 14943
rect 12173 14909 12207 14943
rect 12633 14909 12667 14943
rect 12909 14909 12943 14943
rect 13185 14909 13219 14943
rect 14933 14909 14967 14943
rect 15025 14909 15059 14943
rect 15281 14909 15315 14943
rect 17610 14909 17644 14943
rect 17877 14909 17911 14943
rect 18153 14909 18187 14943
rect 18521 14909 18555 14943
rect 18889 14909 18923 14943
rect 3516 14841 3550 14875
rect 5356 14841 5390 14875
rect 8033 14841 8067 14875
rect 8861 14841 8895 14875
rect 14666 14841 14700 14875
rect 2789 14773 2823 14807
rect 4629 14773 4663 14807
rect 6469 14773 6503 14807
rect 7205 14773 7239 14807
rect 8585 14773 8619 14807
rect 9413 14773 9447 14807
rect 9965 14773 9999 14807
rect 11621 14773 11655 14807
rect 12081 14773 12115 14807
rect 12817 14773 12851 14807
rect 13553 14773 13587 14807
rect 16405 14773 16439 14807
rect 16497 14773 16531 14807
rect 18061 14773 18095 14807
rect 1133 14569 1167 14603
rect 1685 14569 1719 14603
rect 5917 14569 5951 14603
rect 6193 14569 6227 14603
rect 10701 14569 10735 14603
rect 17417 14569 17451 14603
rect 8677 14501 8711 14535
rect 13369 14501 13403 14535
rect 16405 14501 16439 14535
rect 18981 14501 19015 14535
rect 1225 14433 1259 14467
rect 1501 14433 1535 14467
rect 1593 14433 1627 14467
rect 2053 14423 2087 14457
rect 2145 14433 2179 14467
rect 2401 14433 2435 14467
rect 6009 14433 6043 14467
rect 6285 14433 6319 14467
rect 6377 14433 6411 14467
rect 6837 14433 6871 14467
rect 7113 14433 7147 14467
rect 7389 14433 7423 14467
rect 7665 14433 7699 14467
rect 9036 14433 9070 14467
rect 10517 14433 10551 14467
rect 10793 14433 10827 14467
rect 12101 14433 12135 14467
rect 13645 14433 13679 14467
rect 13912 14433 13946 14467
rect 16313 14433 16347 14467
rect 16497 14433 16531 14467
rect 16681 14433 16715 14467
rect 18541 14433 18575 14467
rect 18889 14433 18923 14467
rect 7941 14365 7975 14399
rect 8769 14365 8803 14399
rect 10425 14365 10459 14399
rect 12357 14365 12391 14399
rect 12541 14365 12575 14399
rect 18797 14365 18831 14399
rect 6469 14297 6503 14331
rect 7021 14297 7055 14331
rect 1409 14229 1443 14263
rect 1961 14229 1995 14263
rect 3525 14229 3559 14263
rect 6745 14229 6779 14263
rect 7297 14229 7331 14263
rect 7573 14229 7607 14263
rect 10149 14229 10183 14263
rect 10977 14229 11011 14263
rect 15025 14229 15059 14263
rect 16129 14229 16163 14263
rect 1593 14025 1627 14059
rect 1869 14025 1903 14059
rect 5089 14025 5123 14059
rect 8033 14025 8067 14059
rect 12725 14025 12759 14059
rect 13093 14025 13127 14059
rect 13921 14025 13955 14059
rect 16957 14025 16991 14059
rect 18797 14025 18831 14059
rect 8769 13957 8803 13991
rect 9045 13957 9079 13991
rect 3709 13889 3743 13923
rect 13645 13889 13679 13923
rect 14473 13889 14507 13923
rect 1685 13821 1719 13855
rect 1777 13821 1811 13855
rect 2053 13821 2087 13855
rect 2513 13821 2547 13855
rect 2789 13821 2823 13855
rect 2881 13821 2915 13855
rect 3433 13821 3467 13855
rect 5641 13821 5675 13855
rect 5908 13821 5942 13855
rect 7757 13821 7791 13855
rect 7849 13821 7883 13855
rect 8125 13821 8159 13855
rect 8493 13821 8527 13855
rect 8585 13821 8619 13855
rect 8861 13821 8895 13855
rect 9137 13821 9171 13855
rect 12817 13821 12851 13855
rect 13185 13821 13219 13855
rect 13553 13821 13587 13855
rect 13829 13821 13863 13855
rect 15209 13821 15243 13855
rect 15485 13821 15519 13855
rect 15577 13821 15611 13855
rect 15669 13821 15703 13855
rect 15853 13821 15887 13855
rect 16589 13821 16623 13855
rect 17049 13821 17083 13855
rect 18521 13821 18555 13855
rect 18705 13821 18739 13855
rect 3954 13753 3988 13787
rect 18254 13753 18288 13787
rect 2145 13685 2179 13719
rect 2421 13685 2455 13719
rect 2697 13685 2731 13719
rect 2973 13685 3007 13719
rect 3525 13685 3559 13719
rect 7021 13685 7055 13719
rect 15301 13685 15335 13719
rect 16497 13685 16531 13719
rect 17141 13685 17175 13719
rect 5641 13481 5675 13515
rect 14289 13481 14323 13515
rect 1400 13413 1434 13447
rect 3341 13413 3375 13447
rect 4169 13413 4203 13447
rect 6469 13413 6503 13447
rect 8922 13413 8956 13447
rect 12112 13413 12146 13447
rect 16497 13413 16531 13447
rect 17509 13413 17543 13447
rect 1133 13345 1167 13379
rect 2881 13345 2915 13379
rect 3157 13345 3191 13379
rect 4528 13345 4562 13379
rect 6009 13345 6043 13379
rect 6101 13345 6135 13379
rect 6193 13345 6227 13379
rect 6377 13345 6411 13379
rect 7481 13345 7515 13379
rect 7665 13345 7699 13379
rect 7757 13345 7791 13379
rect 7849 13345 7883 13379
rect 8677 13345 8711 13379
rect 13001 13345 13035 13379
rect 13277 13345 13311 13379
rect 13553 13345 13587 13379
rect 13829 13345 13863 13379
rect 13921 13345 13955 13379
rect 14381 13345 14415 13379
rect 15689 13345 15723 13379
rect 16313 13345 16347 13379
rect 18153 13345 18187 13379
rect 18337 13345 18371 13379
rect 18613 13345 18647 13379
rect 3065 13277 3099 13311
rect 4261 13277 4295 13311
rect 7205 13277 7239 13311
rect 12357 13277 12391 13311
rect 12909 13277 12943 13311
rect 13461 13277 13495 13311
rect 15945 13277 15979 13311
rect 17233 13277 17267 13311
rect 2513 13209 2547 13243
rect 13185 13209 13219 13243
rect 2789 13141 2823 13175
rect 5825 13141 5859 13175
rect 8033 13141 8067 13175
rect 10057 13141 10091 13175
rect 10977 13141 11011 13175
rect 13737 13141 13771 13175
rect 14013 13141 14047 13175
rect 14565 13141 14599 13175
rect 16221 13141 16255 13175
rect 2973 12937 3007 12971
rect 4997 12937 5031 12971
rect 6929 12937 6963 12971
rect 7297 12937 7331 12971
rect 8033 12937 8067 12971
rect 10701 12937 10735 12971
rect 13277 12937 13311 12971
rect 13921 12937 13955 12971
rect 14197 12937 14231 12971
rect 15393 12937 15427 12971
rect 18337 12937 18371 12971
rect 18797 12937 18831 12971
rect 6745 12869 6779 12903
rect 8953 12869 8987 12903
rect 4353 12801 4387 12835
rect 4721 12801 4755 12835
rect 5365 12801 5399 12835
rect 7021 12801 7055 12835
rect 7941 12801 7975 12835
rect 10793 12801 10827 12835
rect 14749 12801 14783 12835
rect 14933 12801 14967 12835
rect 2513 12733 2547 12767
rect 2605 12733 2639 12767
rect 3065 12733 3099 12767
rect 3341 12733 3375 12767
rect 3617 12733 3651 12767
rect 4629 12733 4663 12767
rect 4905 12733 4939 12767
rect 5621 12733 5655 12767
rect 7113 12733 7147 12767
rect 8033 12733 8067 12767
rect 8401 12733 8435 12767
rect 8769 12733 8803 12767
rect 9413 12733 9447 12767
rect 9689 12733 9723 12767
rect 9781 12733 9815 12767
rect 10885 12733 10919 12767
rect 12909 12733 12943 12767
rect 13369 12733 13403 12767
rect 13737 12733 13771 12767
rect 13829 12733 13863 12767
rect 14289 12733 14323 12767
rect 14657 12733 14691 12767
rect 15025 12733 15059 12767
rect 17141 12733 17175 12767
rect 17233 12733 17267 12767
rect 18429 12733 18463 12767
rect 18889 12733 18923 12767
rect 2697 12665 2731 12699
rect 6837 12665 6871 12699
rect 7757 12665 7791 12699
rect 8585 12665 8619 12699
rect 8677 12665 8711 12699
rect 9597 12665 9631 12699
rect 10333 12665 10367 12699
rect 10609 12665 10643 12699
rect 16874 12665 16908 12699
rect 18061 12665 18095 12699
rect 2421 12597 2455 12631
rect 3433 12597 3467 12631
rect 8217 12597 8251 12631
rect 9965 12597 9999 12631
rect 11069 12597 11103 12631
rect 13001 12597 13035 12631
rect 13645 12597 13679 12631
rect 15761 12597 15795 12631
rect 2329 12393 2363 12427
rect 3801 12393 3835 12427
rect 7205 12393 7239 12427
rect 9229 12393 9263 12427
rect 10793 12393 10827 12427
rect 17601 12393 17635 12427
rect 1216 12325 1250 12359
rect 2881 12325 2915 12359
rect 3525 12325 3559 12359
rect 5273 12325 5307 12359
rect 9593 12325 9627 12359
rect 10517 12325 10551 12359
rect 14289 12325 14323 12359
rect 2605 12257 2639 12291
rect 2789 12257 2823 12291
rect 2973 12257 3007 12291
rect 3249 12257 3283 12291
rect 3433 12257 3467 12291
rect 3617 12257 3651 12291
rect 4077 12257 4111 12291
rect 4261 12257 4295 12291
rect 4629 12257 4663 12291
rect 5089 12257 5123 12291
rect 5181 12257 5215 12291
rect 5825 12257 5859 12291
rect 6081 12257 6115 12291
rect 7849 12257 7883 12291
rect 8105 12257 8139 12291
rect 9321 12257 9355 12291
rect 9459 12257 9493 12291
rect 9689 12257 9723 12291
rect 10241 12257 10275 12291
rect 10425 12257 10459 12291
rect 10609 12257 10643 12291
rect 12101 12257 12135 12291
rect 12357 12257 12391 12291
rect 13573 12257 13607 12291
rect 13829 12257 13863 12291
rect 14105 12257 14139 12291
rect 14197 12257 14231 12291
rect 14933 12257 14967 12291
rect 15117 12257 15151 12291
rect 15577 12257 15611 12291
rect 15669 12257 15703 12291
rect 16129 12257 16163 12291
rect 16313 12257 16347 12291
rect 16681 12257 16715 12291
rect 17325 12257 17359 12291
rect 18714 12257 18748 12291
rect 18981 12257 19015 12291
rect 949 12189 983 12223
rect 16589 12189 16623 12223
rect 3157 12121 3191 12155
rect 4353 12121 4387 12155
rect 4997 12121 5031 12155
rect 15209 12121 15243 12155
rect 3985 12053 4019 12087
rect 4721 12053 4755 12087
rect 9873 12053 9907 12087
rect 10977 12053 11011 12087
rect 12449 12053 12483 12087
rect 14013 12053 14047 12087
rect 14933 12053 14967 12087
rect 15485 12053 15519 12087
rect 15761 12053 15795 12087
rect 2421 11849 2455 11883
rect 3893 11849 3927 11883
rect 10977 11849 11011 11883
rect 11713 11849 11747 11883
rect 12817 11849 12851 11883
rect 13921 11849 13955 11883
rect 14565 11849 14599 11883
rect 16497 11849 16531 11883
rect 18429 11849 18463 11883
rect 18797 11849 18831 11883
rect 11345 11781 11379 11815
rect 14841 11781 14875 11815
rect 17141 11781 17175 11815
rect 2605 11713 2639 11747
rect 11897 11713 11931 11747
rect 12357 11713 12391 11747
rect 13645 11713 13679 11747
rect 15393 11713 15427 11747
rect 1041 11645 1075 11679
rect 2513 11645 2547 11679
rect 3341 11645 3375 11679
rect 3433 11645 3467 11679
rect 3985 11645 4019 11679
rect 4077 11645 4111 11679
rect 4537 11645 4571 11679
rect 4629 11645 4663 11679
rect 4905 11645 4939 11679
rect 5181 11645 5215 11679
rect 5273 11645 5307 11679
rect 5641 11645 5675 11679
rect 5917 11645 5951 11679
rect 6009 11645 6043 11679
rect 8401 11645 8435 11679
rect 8585 11645 8619 11679
rect 8677 11645 8711 11679
rect 8769 11645 8803 11679
rect 9617 11645 9651 11679
rect 9873 11645 9907 11679
rect 9965 11645 9999 11679
rect 11069 11645 11103 11679
rect 11161 11645 11195 11679
rect 12081 11645 12115 11679
rect 12449 11645 12483 11679
rect 12909 11645 12943 11679
rect 13553 11645 13587 11679
rect 14013 11645 14047 11679
rect 14197 11645 14231 11679
rect 14289 11645 14323 11679
rect 14657 11645 14691 11679
rect 14933 11645 14967 11679
rect 15209 11645 15243 11679
rect 15485 11645 15519 11679
rect 15577 11645 15611 11679
rect 16037 11645 16071 11679
rect 16313 11645 16347 11679
rect 16589 11645 16623 11679
rect 16957 11645 16991 11679
rect 17233 11645 17267 11679
rect 17417 11645 17451 11679
rect 17509 11645 17543 11679
rect 17785 11645 17819 11679
rect 18245 11645 18279 11679
rect 18521 11645 18555 11679
rect 18889 11645 18923 11679
rect 1308 11577 1342 11611
rect 4169 11577 4203 11611
rect 4445 11577 4479 11611
rect 4721 11577 4755 11611
rect 4997 11577 5031 11611
rect 5549 11577 5583 11611
rect 9781 11577 9815 11611
rect 10885 11577 10919 11611
rect 15669 11577 15703 11611
rect 15945 11577 15979 11611
rect 5825 11509 5859 11543
rect 6101 11509 6135 11543
rect 8953 11509 8987 11543
rect 10149 11509 10183 11543
rect 15117 11509 15151 11543
rect 16221 11509 16255 11543
rect 17693 11509 17727 11543
rect 18153 11509 18187 11543
rect 1317 11305 1351 11339
rect 4813 11305 4847 11339
rect 7573 11305 7607 11339
rect 9045 11305 9079 11339
rect 9965 11305 9999 11339
rect 10517 11305 10551 11339
rect 14289 11305 14323 11339
rect 16497 11305 16531 11339
rect 7932 11237 7966 11271
rect 1409 11159 1443 11193
rect 1768 11169 1802 11203
rect 3433 11169 3467 11203
rect 3700 11169 3734 11203
rect 4905 11169 4939 11203
rect 5181 11169 5215 11203
rect 5273 11169 5307 11203
rect 5641 11169 5675 11203
rect 5917 11169 5951 11203
rect 6193 11169 6227 11203
rect 6449 11169 6483 11203
rect 7665 11169 7699 11203
rect 9505 11169 9539 11203
rect 9781 11169 9815 11203
rect 10057 11169 10091 11203
rect 10149 11169 10183 11203
rect 10333 11169 10367 11203
rect 11437 11169 11471 11203
rect 11805 11169 11839 11203
rect 13838 11169 13872 11203
rect 14381 11169 14415 11203
rect 14565 11169 14599 11203
rect 14657 11169 14691 11203
rect 15117 11169 15151 11203
rect 15393 11169 15427 11203
rect 15669 11169 15703 11203
rect 16221 11169 16255 11203
rect 16313 11169 16347 11203
rect 16589 11169 16623 11203
rect 16681 11169 16715 11203
rect 16773 11169 16807 11203
rect 17969 11169 18003 11203
rect 19073 11169 19107 11203
rect 1501 11101 1535 11135
rect 9689 11101 9723 11135
rect 11529 11101 11563 11135
rect 11713 11101 11747 11135
rect 12449 11101 12483 11135
rect 14105 11101 14139 11135
rect 15577 11101 15611 11135
rect 18613 11101 18647 11135
rect 12725 11033 12759 11067
rect 15025 11033 15059 11067
rect 2881 10965 2915 10999
rect 4997 10965 5031 10999
rect 5549 10965 5583 10999
rect 6009 10965 6043 10999
rect 9505 10965 9539 10999
rect 15301 10965 15335 10999
rect 17877 10965 17911 10999
rect 6469 10761 6503 10795
rect 7389 10761 7423 10795
rect 9689 10761 9723 10795
rect 11437 10761 11471 10795
rect 11897 10761 11931 10795
rect 11989 10761 12023 10795
rect 13921 10761 13955 10795
rect 14565 10761 14599 10795
rect 18337 10761 18371 10795
rect 4629 10693 4663 10727
rect 10793 10693 10827 10727
rect 3249 10625 3283 10659
rect 6653 10625 6687 10659
rect 18153 10625 18187 10659
rect 2513 10557 2547 10591
rect 2881 10557 2915 10591
rect 3505 10557 3539 10591
rect 5457 10557 5491 10591
rect 5825 10557 5859 10591
rect 6745 10557 6779 10591
rect 7297 10557 7331 10591
rect 9873 10557 9907 10591
rect 10057 10557 10091 10591
rect 10149 10557 10183 10591
rect 10241 10557 10275 10591
rect 10425 10557 10459 10591
rect 10517 10557 10551 10591
rect 10609 10557 10643 10591
rect 11437 10557 11471 10591
rect 11621 10557 11655 10591
rect 11713 10557 11747 10591
rect 12173 10557 12207 10591
rect 12265 10557 12299 10591
rect 13829 10557 13863 10591
rect 14657 10557 14691 10591
rect 15301 10557 15335 10591
rect 18245 10557 18279 10591
rect 18705 10557 18739 10591
rect 2697 10489 2731 10523
rect 2789 10489 2823 10523
rect 6469 10489 6503 10523
rect 11989 10489 12023 10523
rect 15568 10489 15602 10523
rect 17886 10489 17920 10523
rect 18797 10489 18831 10523
rect 3065 10421 3099 10455
rect 5549 10421 5583 10455
rect 5917 10421 5951 10455
rect 6929 10421 6963 10455
rect 11161 10421 11195 10455
rect 12449 10421 12483 10455
rect 16681 10421 16715 10455
rect 16773 10421 16807 10455
rect 6469 10217 6503 10251
rect 9321 10217 9355 10251
rect 12265 10217 12299 10251
rect 1492 10149 1526 10183
rect 10965 10149 10999 10183
rect 18622 10149 18656 10183
rect 1225 10081 1259 10115
rect 5457 10081 5491 10115
rect 6009 10081 6043 10115
rect 6101 10081 6135 10115
rect 6561 10081 6595 10115
rect 6745 10081 6779 10115
rect 7001 10081 7035 10115
rect 9505 10081 9539 10115
rect 9781 10081 9815 10115
rect 14482 10081 14516 10115
rect 14749 10081 14783 10115
rect 16313 10081 16347 10115
rect 16681 10081 16715 10115
rect 18889 10081 18923 10115
rect 9597 10013 9631 10047
rect 16405 10013 16439 10047
rect 16589 10013 16623 10047
rect 17233 10013 17267 10047
rect 2605 9945 2639 9979
rect 8125 9945 8159 9979
rect 5549 9877 5583 9911
rect 5917 9877 5951 9911
rect 6193 9877 6227 9911
rect 9781 9877 9815 9911
rect 13369 9877 13403 9911
rect 17509 9877 17543 9911
rect 2421 9673 2455 9707
rect 11621 9673 11655 9707
rect 18797 9673 18831 9707
rect 6285 9605 6319 9639
rect 12357 9537 12391 9571
rect 12541 9537 12575 9571
rect 15853 9537 15887 9571
rect 17141 9537 17175 9571
rect 1041 9469 1075 9503
rect 4721 9469 4755 9503
rect 4905 9469 4939 9503
rect 4997 9469 5031 9503
rect 5089 9469 5123 9503
rect 5457 9469 5491 9503
rect 5825 9469 5859 9503
rect 5917 9469 5951 9503
rect 6193 9469 6227 9503
rect 6653 9469 6687 9503
rect 9045 9469 9079 9503
rect 9301 9469 9335 9503
rect 11069 9469 11103 9503
rect 11253 9469 11287 9503
rect 11345 9469 11379 9503
rect 11437 9469 11471 9503
rect 12265 9469 12299 9503
rect 12633 9469 12667 9503
rect 13737 9469 13771 9503
rect 14013 9469 14047 9503
rect 14105 9469 14139 9503
rect 17049 9469 17083 9503
rect 17408 9469 17442 9503
rect 18705 9469 18739 9503
rect 1286 9401 1320 9435
rect 5273 9401 5307 9435
rect 5365 9401 5399 9435
rect 6898 9401 6932 9435
rect 13921 9401 13955 9435
rect 15586 9401 15620 9435
rect 16957 9401 16991 9435
rect 4629 9333 4663 9367
rect 5641 9333 5675 9367
rect 8033 9333 8067 9367
rect 10425 9333 10459 9367
rect 13185 9333 13219 9367
rect 14289 9333 14323 9367
rect 14473 9333 14507 9367
rect 18521 9333 18555 9367
rect 1409 9129 1443 9163
rect 5089 9129 5123 9163
rect 9597 9129 9631 9163
rect 12081 9129 12115 9163
rect 13277 9129 13311 9163
rect 14657 9129 14691 9163
rect 18153 9129 18187 9163
rect 18889 9129 18923 9163
rect 4721 9061 4755 9095
rect 7840 9061 7874 9095
rect 9321 9061 9355 9095
rect 11253 9061 11287 9095
rect 13737 9061 13771 9095
rect 16948 9061 16982 9095
rect 1317 8993 1351 9027
rect 1849 8993 1883 9027
rect 3065 8993 3099 9027
rect 3321 8993 3355 9027
rect 4537 8993 4571 9027
rect 4813 8993 4847 9027
rect 4905 8993 4939 9027
rect 5365 8993 5399 9027
rect 5549 8993 5583 9027
rect 5641 8993 5675 9027
rect 6009 8993 6043 9027
rect 6101 8993 6135 9027
rect 6561 8993 6595 9027
rect 7573 8993 7607 9027
rect 9045 8993 9079 9027
rect 9229 8993 9263 9027
rect 9413 8993 9447 9027
rect 10241 8993 10275 9027
rect 10425 8993 10459 9027
rect 10517 8993 10551 9027
rect 10609 8993 10643 9027
rect 10977 8993 11011 9027
rect 11161 8993 11195 9027
rect 11345 8993 11379 9027
rect 11621 8993 11655 9027
rect 11897 8993 11931 9027
rect 12265 8993 12299 9027
rect 12357 8993 12391 9027
rect 12725 8993 12759 9027
rect 12909 8993 12943 9027
rect 13461 8993 13495 9027
rect 13645 8993 13679 9027
rect 13829 8993 13863 9027
rect 14197 8993 14231 9027
rect 14381 8993 14415 9027
rect 14473 8993 14507 9027
rect 14749 8993 14783 9027
rect 14933 8993 14967 9027
rect 15301 8993 15335 9027
rect 15485 8993 15519 9027
rect 16681 8993 16715 9027
rect 18337 8993 18371 9027
rect 18429 8993 18463 9027
rect 18521 8993 18555 9027
rect 18705 8993 18739 9027
rect 18797 8993 18831 9027
rect 1593 8925 1627 8959
rect 11805 8925 11839 8959
rect 15945 8925 15979 8959
rect 5273 8857 5307 8891
rect 6193 8857 6227 8891
rect 8953 8857 8987 8891
rect 10793 8857 10827 8891
rect 18061 8857 18095 8891
rect 2973 8789 3007 8823
rect 4445 8789 4479 8823
rect 5917 8789 5951 8823
rect 6469 8789 6503 8823
rect 11529 8789 11563 8823
rect 11621 8789 11655 8823
rect 14013 8789 14047 8823
rect 14197 8789 14231 8823
rect 2329 8585 2363 8619
rect 9045 8585 9079 8619
rect 9505 8585 9539 8619
rect 10977 8585 11011 8619
rect 11805 8585 11839 8619
rect 12771 8585 12805 8619
rect 17693 8585 17727 8619
rect 7389 8517 7423 8551
rect 9781 8517 9815 8551
rect 18429 8517 18463 8551
rect 12081 8449 12115 8483
rect 12173 8449 12207 8483
rect 17417 8449 17451 8483
rect 1409 8381 1443 8415
rect 1685 8381 1719 8415
rect 1961 8381 1995 8415
rect 2421 8381 2455 8415
rect 4629 8381 4663 8415
rect 4905 8381 4939 8415
rect 5181 8381 5215 8415
rect 5457 8381 5491 8415
rect 5733 8381 5767 8415
rect 6009 8381 6043 8415
rect 6276 8381 6310 8415
rect 8401 8381 8435 8415
rect 8769 8381 8803 8415
rect 9045 8381 9079 8415
rect 9229 8381 9263 8415
rect 9321 8381 9355 8415
rect 9965 8381 9999 8415
rect 11253 8381 11287 8415
rect 11437 8381 11471 8415
rect 11529 8381 11563 8415
rect 11645 8381 11679 8415
rect 11989 8381 12023 8415
rect 12265 8381 12299 8415
rect 12541 8381 12575 8415
rect 13553 8381 13587 8415
rect 13820 8381 13854 8415
rect 16037 8381 16071 8415
rect 16313 8381 16347 8415
rect 16405 8381 16439 8415
rect 17877 8381 17911 8415
rect 18245 8381 18279 8415
rect 18337 8381 18371 8415
rect 18705 8381 18739 8415
rect 1317 8313 1351 8347
rect 1593 8313 1627 8347
rect 8585 8313 8619 8347
rect 8677 8313 8711 8347
rect 10057 8313 10091 8347
rect 10333 8313 10367 8347
rect 11069 8313 11103 8347
rect 12449 8313 12483 8347
rect 16221 8313 16255 8347
rect 16681 8313 16715 8347
rect 17969 8313 18003 8347
rect 18061 8313 18095 8347
rect 1869 8245 1903 8279
rect 4537 8245 4571 8279
rect 4813 8245 4847 8279
rect 5089 8245 5123 8279
rect 5365 8245 5399 8279
rect 5641 8245 5675 8279
rect 8953 8245 8987 8279
rect 10149 8245 10183 8279
rect 14933 8245 14967 8279
rect 16589 8245 16623 8279
rect 18797 8245 18831 8279
rect 1225 8041 1259 8075
rect 1777 8041 1811 8075
rect 2329 8041 2363 8075
rect 8861 8041 8895 8075
rect 10701 8041 10735 8075
rect 12357 8041 12391 8075
rect 13645 8041 13679 8075
rect 15393 8041 15427 8075
rect 16589 8041 16623 8075
rect 17693 8041 17727 8075
rect 7288 7973 7322 8007
rect 11161 7973 11195 8007
rect 12909 7973 12943 8007
rect 15025 7973 15059 8007
rect 17141 7973 17175 8007
rect 1041 7905 1075 7939
rect 1317 7905 1351 7939
rect 1409 7905 1443 7939
rect 1501 7905 1535 7939
rect 1685 7905 1719 7939
rect 2145 7905 2179 7939
rect 2421 7905 2455 7939
rect 2789 7905 2823 7939
rect 3157 7905 3191 7939
rect 3985 7905 4019 7939
rect 4353 7905 4387 7939
rect 4629 7905 4663 7939
rect 4905 7905 4939 7939
rect 5181 7905 5215 7939
rect 5457 7905 5491 7939
rect 7021 7905 7055 7939
rect 8953 7905 8987 7939
rect 9597 7905 9631 7939
rect 10057 7905 10091 7939
rect 10149 7905 10183 7939
rect 10241 7905 10275 7939
rect 10517 7905 10551 7939
rect 11529 7905 11563 7939
rect 11621 7905 11655 7939
rect 12081 7905 12115 7939
rect 12725 7905 12759 7939
rect 12817 7905 12851 7939
rect 13093 7905 13127 7939
rect 13277 7905 13311 7939
rect 13369 7905 13403 7939
rect 13829 7905 13863 7939
rect 14105 7905 14139 7939
rect 14289 7905 14323 7939
rect 14749 7905 14783 7939
rect 14933 7905 14967 7939
rect 15117 7905 15151 7939
rect 15577 7905 15611 7939
rect 15669 7905 15703 7939
rect 15761 7905 15795 7939
rect 15945 7905 15979 7939
rect 16129 7905 16163 7939
rect 16405 7905 16439 7939
rect 16865 7905 16899 7939
rect 17233 7905 17267 7939
rect 18806 7905 18840 7939
rect 19073 7905 19107 7939
rect 2697 7837 2731 7871
rect 9689 7837 9723 7871
rect 11069 7837 11103 7871
rect 12173 7837 12207 7871
rect 13921 7837 13955 7871
rect 14473 7837 14507 7871
rect 16313 7837 16347 7871
rect 949 7769 983 7803
rect 3065 7769 3099 7803
rect 5365 7769 5399 7803
rect 15301 7769 15335 7803
rect 2053 7701 2087 7735
rect 3893 7701 3927 7735
rect 4261 7701 4295 7735
rect 4537 7701 4571 7735
rect 4813 7701 4847 7735
rect 5089 7701 5123 7735
rect 8401 7701 8435 7735
rect 13093 7701 13127 7735
rect 13553 7701 13587 7735
rect 14013 7701 14047 7735
rect 16405 7701 16439 7735
rect 1041 7497 1075 7531
rect 1317 7497 1351 7531
rect 2145 7497 2179 7531
rect 2421 7497 2455 7531
rect 2697 7497 2731 7531
rect 7021 7497 7055 7531
rect 9965 7497 9999 7531
rect 14105 7497 14139 7531
rect 14473 7497 14507 7531
rect 14749 7497 14783 7531
rect 16313 7497 16347 7531
rect 18245 7497 18279 7531
rect 18889 7497 18923 7531
rect 4813 7429 4847 7463
rect 13553 7429 13587 7463
rect 4445 7361 4479 7395
rect 4997 7361 5031 7395
rect 7941 7361 7975 7395
rect 8861 7361 8895 7395
rect 11161 7361 11195 7395
rect 12173 7361 12207 7395
rect 13185 7361 13219 7395
rect 17969 7361 18003 7395
rect 1133 7293 1167 7327
rect 1409 7293 1443 7327
rect 1685 7293 1719 7327
rect 1961 7293 1995 7327
rect 2237 7293 2271 7327
rect 2513 7293 2547 7327
rect 2789 7293 2823 7327
rect 3065 7293 3099 7327
rect 3617 7293 3651 7327
rect 4905 7293 4939 7327
rect 6469 7293 6503 7327
rect 6653 7293 6687 7327
rect 6837 7293 6871 7327
rect 7205 7293 7239 7327
rect 9321 7293 9355 7327
rect 9781 7293 9815 7327
rect 10149 7293 10183 7327
rect 10425 7293 10459 7327
rect 10701 7293 10735 7327
rect 10885 7293 10919 7327
rect 11253 7293 11287 7327
rect 11621 7293 11655 7327
rect 11713 7293 11747 7327
rect 12265 7293 12299 7327
rect 12817 7293 12851 7327
rect 13921 7293 13955 7327
rect 14289 7293 14323 7327
rect 14841 7293 14875 7327
rect 15853 7271 15887 7305
rect 16129 7293 16163 7327
rect 17518 7293 17552 7327
rect 17785 7293 17819 7327
rect 17877 7293 17911 7327
rect 18337 7293 18371 7327
rect 18789 7293 18823 7327
rect 1869 7225 1903 7259
rect 3709 7225 3743 7259
rect 5264 7225 5298 7259
rect 6745 7225 6779 7259
rect 8769 7225 8803 7259
rect 8953 7225 8987 7259
rect 9229 7225 9263 7259
rect 12725 7225 12759 7259
rect 13277 7225 13311 7259
rect 13737 7225 13771 7259
rect 1593 7157 1627 7191
rect 2973 7157 3007 7191
rect 3525 7157 3559 7191
rect 6377 7157 6411 7191
rect 8585 7157 8619 7191
rect 9597 7157 9631 7191
rect 9689 7157 9723 7191
rect 10241 7157 10275 7191
rect 15945 7157 15979 7191
rect 16405 7157 16439 7191
rect 3341 6953 3375 6987
rect 9873 6953 9907 6987
rect 13369 6953 13403 6987
rect 17509 6953 17543 6987
rect 8677 6885 8711 6919
rect 11897 6885 11931 6919
rect 16497 6885 16531 6919
rect 1133 6817 1167 6851
rect 1409 6817 1443 6851
rect 1665 6817 1699 6851
rect 2965 6817 2999 6851
rect 3433 6817 3467 6851
rect 3709 6817 3743 6851
rect 4077 6817 4111 6851
rect 4169 6817 4203 6851
rect 4436 6817 4470 6851
rect 6184 6817 6218 6851
rect 7665 6817 7699 6851
rect 8401 6817 8435 6851
rect 8585 6817 8619 6851
rect 8769 6817 8803 6851
rect 9045 6817 9079 6851
rect 9229 6817 9263 6851
rect 9321 6817 9355 6851
rect 9413 6817 9447 6851
rect 9965 6817 9999 6851
rect 10241 6817 10275 6851
rect 10425 6817 10459 6851
rect 11437 6817 11471 6851
rect 11621 6817 11655 6851
rect 12541 6817 12575 6851
rect 12633 6817 12667 6851
rect 13185 6817 13219 6851
rect 13912 6817 13946 6851
rect 17233 6817 17267 6851
rect 18622 6817 18656 6851
rect 18889 6817 18923 6851
rect 5917 6749 5951 6783
rect 10793 6749 10827 6783
rect 11529 6749 11563 6783
rect 11713 6749 11747 6783
rect 12081 6749 12115 6783
rect 12173 6749 12207 6783
rect 13093 6749 13127 6783
rect 13645 6749 13679 6783
rect 2789 6681 2823 6715
rect 7573 6681 7607 6715
rect 1041 6613 1075 6647
rect 3065 6613 3099 6647
rect 3617 6613 3651 6647
rect 3985 6613 4019 6647
rect 5549 6613 5583 6647
rect 7297 6613 7331 6647
rect 8953 6613 8987 6647
rect 9597 6613 9631 6647
rect 15025 6613 15059 6647
rect 1225 6409 1259 6443
rect 2973 6409 3007 6443
rect 15853 6409 15887 6443
rect 16129 6409 16163 6443
rect 18153 6409 18187 6443
rect 18429 6409 18463 6443
rect 949 6341 983 6375
rect 9413 6341 9447 6375
rect 10977 6341 11011 6375
rect 16037 6341 16071 6375
rect 3525 6273 3559 6307
rect 6837 6273 6871 6307
rect 11437 6273 11471 6307
rect 12449 6273 12483 6307
rect 14657 6273 14691 6307
rect 18797 6273 18831 6307
rect 1041 6205 1075 6239
rect 1317 6205 1351 6239
rect 1593 6205 1627 6239
rect 1869 6205 1903 6239
rect 2145 6205 2179 6239
rect 3065 6205 3099 6239
rect 3433 6205 3467 6239
rect 3977 6205 4011 6239
rect 4997 6205 5031 6239
rect 5273 6205 5307 6239
rect 5641 6205 5675 6239
rect 5825 6205 5859 6239
rect 6009 6205 6043 6239
rect 7104 6205 7138 6239
rect 8861 6205 8895 6239
rect 9137 6205 9171 6239
rect 9229 6205 9263 6239
rect 11161 6205 11195 6239
rect 11897 6205 11931 6239
rect 14105 6205 14139 6239
rect 14197 6205 14231 6239
rect 14289 6205 14323 6239
rect 14473 6205 14507 6239
rect 15761 6205 15795 6239
rect 15853 6205 15887 6239
rect 16313 6205 16347 6239
rect 16405 6205 16439 6239
rect 16681 6205 16715 6239
rect 17233 6205 17267 6239
rect 17325 6205 17359 6239
rect 17785 6205 17819 6239
rect 17877 6205 17911 6239
rect 18245 6205 18279 6239
rect 18337 6205 18371 6239
rect 18705 6205 18739 6239
rect 1961 6137 1995 6171
rect 2237 6137 2271 6171
rect 4261 6137 4295 6171
rect 5917 6137 5951 6171
rect 9045 6137 9079 6171
rect 11529 6137 11563 6171
rect 11989 6137 12023 6171
rect 15485 6137 15519 6171
rect 15577 6137 15611 6171
rect 16497 6137 16531 6171
rect 1685 6069 1719 6103
rect 3893 6069 3927 6103
rect 5181 6069 5215 6103
rect 6193 6069 6227 6103
rect 8217 6069 8251 6103
rect 13921 6069 13955 6103
rect 1409 5865 1443 5899
rect 2973 5865 3007 5899
rect 6377 5865 6411 5899
rect 8401 5865 8435 5899
rect 15117 5865 15151 5899
rect 16681 5865 16715 5899
rect 17049 5865 17083 5899
rect 17877 5865 17911 5899
rect 18153 5865 18187 5899
rect 18429 5865 18463 5899
rect 6101 5797 6135 5831
rect 7266 5797 7300 5831
rect 8769 5797 8803 5831
rect 12265 5797 12299 5831
rect 13268 5797 13302 5831
rect 14749 5797 14783 5831
rect 17325 5797 17359 5831
rect 17601 5797 17635 5831
rect 1317 5729 1351 5763
rect 1777 5729 1811 5763
rect 1869 5729 1903 5763
rect 3065 5719 3099 5753
rect 3157 5729 3191 5763
rect 3424 5729 3458 5763
rect 4629 5729 4663 5763
rect 5825 5729 5859 5763
rect 6009 5729 6043 5763
rect 6193 5729 6227 5763
rect 7021 5729 7055 5763
rect 8493 5729 8527 5763
rect 8677 5729 8711 5763
rect 8861 5729 8895 5763
rect 9137 5729 9171 5763
rect 9321 5729 9355 5763
rect 9413 5729 9447 5763
rect 9505 5729 9539 5763
rect 11161 5729 11195 5763
rect 11345 5729 11379 5763
rect 11529 5729 11563 5763
rect 11713 5729 11747 5763
rect 12449 5729 12483 5763
rect 14565 5729 14599 5763
rect 14841 5729 14875 5763
rect 14933 5729 14967 5763
rect 15393 5729 15427 5763
rect 15485 5729 15519 5763
rect 15577 5729 15611 5763
rect 15761 5729 15795 5763
rect 16313 5729 16347 5763
rect 16497 5729 16531 5763
rect 16589 5729 16623 5763
rect 16865 5729 16899 5763
rect 17141 5729 17175 5763
rect 17417 5729 17451 5763
rect 17693 5729 17727 5763
rect 17969 5729 18003 5763
rect 18245 5729 18279 5763
rect 18521 5729 18555 5763
rect 13001 5661 13035 5695
rect 4721 5593 4755 5627
rect 9689 5593 9723 5627
rect 11989 5593 12023 5627
rect 14381 5593 14415 5627
rect 1685 5525 1719 5559
rect 1961 5525 1995 5559
rect 4537 5525 4571 5559
rect 9045 5525 9079 5559
rect 15209 5525 15243 5559
rect 16129 5525 16163 5559
rect 1409 5321 1443 5355
rect 3065 5321 3099 5355
rect 6561 5321 6595 5355
rect 9505 5321 9539 5355
rect 10977 5321 11011 5355
rect 13553 5321 13587 5355
rect 14105 5321 14139 5355
rect 15301 5321 15335 5355
rect 15117 5253 15151 5287
rect 1133 5185 1167 5219
rect 15485 5185 15519 5219
rect 1225 5117 1259 5151
rect 1317 5117 1351 5151
rect 1685 5117 1719 5151
rect 3709 5117 3743 5151
rect 5181 5117 5215 5151
rect 5448 5117 5482 5151
rect 9321 5117 9355 5151
rect 9689 5117 9723 5151
rect 10057 5117 10091 5151
rect 10425 5117 10459 5151
rect 10701 5117 10735 5151
rect 10793 5117 10827 5151
rect 11437 5117 11471 5151
rect 11529 5117 11563 5151
rect 11989 5117 12023 5151
rect 13369 5117 13403 5151
rect 13737 5117 13771 5151
rect 14013 5117 14047 5151
rect 14289 5117 14323 5151
rect 14565 5117 14599 5151
rect 15301 5117 15335 5151
rect 15577 5117 15611 5151
rect 18153 5117 18187 5151
rect 18245 5117 18279 5151
rect 18705 5117 18739 5151
rect 1952 5049 1986 5083
rect 3976 5049 4010 5083
rect 8585 5049 8619 5083
rect 9781 5049 9815 5083
rect 9873 5049 9907 5083
rect 10609 5049 10643 5083
rect 11345 5049 11379 5083
rect 11897 5049 11931 5083
rect 12541 5049 12575 5083
rect 17886 5049 17920 5083
rect 5089 4981 5123 5015
rect 13921 4981 13955 5015
rect 14473 4981 14507 5015
rect 16773 4981 16807 5015
rect 18337 4981 18371 5015
rect 18797 4981 18831 5015
rect 1409 4777 1443 4811
rect 2973 4777 3007 4811
rect 5273 4777 5307 4811
rect 7481 4777 7515 4811
rect 9413 4777 9447 4811
rect 12173 4777 12207 4811
rect 15945 4777 15979 4811
rect 17693 4777 17727 4811
rect 1838 4709 1872 4743
rect 9076 4709 9110 4743
rect 11805 4709 11839 4743
rect 12449 4709 12483 4743
rect 12541 4709 12575 4743
rect 17049 4709 17083 4743
rect 17417 4709 17451 4743
rect 1225 4641 1259 4675
rect 1501 4641 1535 4675
rect 4160 4641 4194 4675
rect 6368 4641 6402 4675
rect 10526 4641 10560 4675
rect 10977 4641 11011 4675
rect 11069 4641 11103 4675
rect 11253 4641 11287 4675
rect 11437 4641 11471 4675
rect 11529 4641 11563 4675
rect 11713 4641 11747 4675
rect 11897 4641 11931 4675
rect 12357 4641 12391 4675
rect 12725 4641 12759 4675
rect 14832 4641 14866 4675
rect 16957 4641 16991 4675
rect 17509 4641 17543 4675
rect 18806 4641 18840 4675
rect 19073 4641 19107 4675
rect 1593 4573 1627 4607
rect 3893 4573 3927 4607
rect 6101 4573 6135 4607
rect 9321 4573 9355 4607
rect 10793 4573 10827 4607
rect 14565 4573 14599 4607
rect 12081 4505 12115 4539
rect 1133 4437 1167 4471
rect 7941 4437 7975 4471
rect 1501 4233 1535 4267
rect 10149 4233 10183 4267
rect 10609 4233 10643 4267
rect 13553 4233 13587 4267
rect 18337 4233 18371 4267
rect 18797 4233 18831 4267
rect 17785 4165 17819 4199
rect 5089 4097 5123 4131
rect 6837 4097 6871 4131
rect 16313 4097 16347 4131
rect 18061 4097 18095 4131
rect 1409 4029 1443 4063
rect 1685 4029 1719 4063
rect 1961 4029 1995 4063
rect 8769 4029 8803 4063
rect 9036 4029 9070 4063
rect 10517 4029 10551 4063
rect 11621 4029 11655 4063
rect 14933 4029 14967 4063
rect 15485 4029 15519 4063
rect 15669 4029 15703 4063
rect 15761 4029 15795 4063
rect 16129 4029 16163 4063
rect 16221 4029 16255 4063
rect 16681 4029 16715 4063
rect 16957 4029 16991 4063
rect 17233 4029 17267 4063
rect 17417 4029 17451 4063
rect 17877 4029 17911 4063
rect 17969 4029 18003 4063
rect 18429 4029 18463 4063
rect 18705 4029 18739 4063
rect 1777 3961 1811 3995
rect 5356 3961 5390 3995
rect 7104 3961 7138 3995
rect 11888 3961 11922 3995
rect 14666 3961 14700 3995
rect 15393 3961 15427 3995
rect 16037 3961 16071 3995
rect 16865 3961 16899 3995
rect 17141 3961 17175 3995
rect 17509 3961 17543 3995
rect 2053 3893 2087 3927
rect 6469 3893 6503 3927
rect 8217 3893 8251 3927
rect 13001 3893 13035 3927
rect 16589 3893 16623 3927
rect 1133 3689 1167 3723
rect 4997 3689 5031 3723
rect 5457 3689 5491 3723
rect 8125 3689 8159 3723
rect 10609 3689 10643 3723
rect 14381 3689 14415 3723
rect 14841 3689 14875 3723
rect 15485 3689 15519 3723
rect 16221 3689 16255 3723
rect 16773 3689 16807 3723
rect 17049 3689 17083 3723
rect 17601 3689 17635 3723
rect 18714 3621 18748 3655
rect 1225 3553 1259 3587
rect 1317 3553 1351 3587
rect 1777 3553 1811 3587
rect 2228 3553 2262 3587
rect 3617 3553 3651 3587
rect 3873 3553 3907 3587
rect 5365 3553 5399 3587
rect 6285 3553 6319 3587
rect 7001 3553 7035 3587
rect 9485 3553 9519 3587
rect 13001 3553 13035 3587
rect 13257 3553 13291 3587
rect 14749 3553 14783 3587
rect 15577 3553 15611 3587
rect 15669 3553 15703 3587
rect 16129 3553 16163 3587
rect 16405 3553 16439 3587
rect 16865 3553 16899 3587
rect 16957 3553 16991 3587
rect 17233 3553 17267 3587
rect 18981 3553 19015 3587
rect 1961 3485 1995 3519
rect 6745 3485 6779 3519
rect 9229 3485 9263 3519
rect 1409 3417 1443 3451
rect 16497 3417 16531 3451
rect 1685 3349 1719 3383
rect 3341 3349 3375 3383
rect 6377 3349 6411 3383
rect 15761 3349 15795 3383
rect 17325 3349 17359 3383
rect 3065 3145 3099 3179
rect 7297 3145 7331 3179
rect 7757 3145 7791 3179
rect 8769 3145 8803 3179
rect 10885 3145 10919 3179
rect 12909 3145 12943 3179
rect 15117 3145 15151 3179
rect 15393 3145 15427 3179
rect 15761 3145 15795 3179
rect 16129 3145 16163 3179
rect 17141 3145 17175 3179
rect 12265 3009 12299 3043
rect 14841 3009 14875 3043
rect 18521 3009 18555 3043
rect 1317 2941 1351 2975
rect 1593 2941 1627 2975
rect 1685 2941 1719 2975
rect 3249 2941 3283 2975
rect 5733 2941 5767 2975
rect 7021 2941 7055 2975
rect 7205 2941 7239 2975
rect 7665 2941 7699 2975
rect 8677 2941 8711 2975
rect 12817 2941 12851 2975
rect 14749 2941 14783 2975
rect 15209 2941 15243 2975
rect 15301 2941 15335 2975
rect 15669 2941 15703 2975
rect 16221 2941 16255 2975
rect 16497 2941 16531 2975
rect 16589 2941 16623 2975
rect 17049 2941 17083 2975
rect 1952 2873 1986 2907
rect 3341 2873 3375 2907
rect 12020 2873 12054 2907
rect 18254 2873 18288 2907
rect 1225 2805 1259 2839
rect 1501 2805 1535 2839
rect 5825 2805 5859 2839
rect 6929 2805 6963 2839
rect 16405 2805 16439 2839
rect 16681 2805 16715 2839
rect 16957 2805 16991 2839
rect 1961 2601 1995 2635
rect 3801 2601 3835 2635
rect 5273 2601 5307 2635
rect 6377 2601 6411 2635
rect 10609 2601 10643 2635
rect 13829 2601 13863 2635
rect 15485 2601 15519 2635
rect 16773 2601 16807 2635
rect 17141 2601 17175 2635
rect 17601 2601 17635 2635
rect 1685 2533 1719 2567
rect 3157 2533 3191 2567
rect 4353 2533 4387 2567
rect 4905 2533 4939 2567
rect 6806 2533 6840 2567
rect 9597 2533 9631 2567
rect 10241 2533 10275 2567
rect 16497 2533 16531 2567
rect 1225 2465 1259 2499
rect 1501 2465 1535 2499
rect 1593 2465 1627 2499
rect 2053 2465 2087 2499
rect 2329 2465 2363 2499
rect 2421 2465 2455 2499
rect 2789 2465 2823 2499
rect 3065 2465 3099 2499
rect 3617 2465 3651 2499
rect 3709 2465 3743 2499
rect 4169 2465 4203 2499
rect 4261 2465 4295 2499
rect 4537 2465 4571 2499
rect 4997 2465 5031 2499
rect 5181 2465 5215 2499
rect 5641 2465 5675 2499
rect 6009 2465 6043 2499
rect 6285 2465 6319 2499
rect 6561 2465 6595 2499
rect 8309 2465 8343 2499
rect 8585 2465 8619 2499
rect 8769 2465 8803 2499
rect 9045 2465 9079 2499
rect 9413 2465 9447 2499
rect 9689 2465 9723 2499
rect 9781 2465 9815 2499
rect 10057 2465 10091 2499
rect 10333 2465 10367 2499
rect 10425 2465 10459 2499
rect 10977 2465 11011 2499
rect 11069 2465 11103 2499
rect 11437 2465 11471 2499
rect 12449 2465 12483 2499
rect 12716 2465 12750 2499
rect 13921 2465 13955 2499
rect 14177 2465 14211 2499
rect 15577 2465 15611 2499
rect 15669 2465 15703 2499
rect 16313 2465 16347 2499
rect 16405 2465 16439 2499
rect 16681 2465 16715 2499
rect 17049 2465 17083 2499
rect 17693 2465 17727 2499
rect 1133 2397 1167 2431
rect 4629 2397 4663 2431
rect 4077 2329 4111 2363
rect 7941 2329 7975 2363
rect 1409 2261 1443 2295
rect 2881 2261 2915 2295
rect 3525 2261 3559 2295
rect 5549 2261 5583 2295
rect 6101 2261 6135 2295
rect 8217 2261 8251 2295
rect 8493 2261 8527 2295
rect 8861 2261 8895 2295
rect 9137 2261 9171 2295
rect 9965 2261 9999 2295
rect 11345 2261 11379 2295
rect 15301 2261 15335 2295
rect 15761 2261 15795 2295
rect 16221 2261 16255 2295
rect 19073 2261 19107 2295
rect 1317 2057 1351 2091
rect 1869 2057 1903 2091
rect 2973 2057 3007 2091
rect 7021 2057 7055 2091
rect 7573 2057 7607 2091
rect 8585 2057 8619 2091
rect 10425 2057 10459 2091
rect 10701 2057 10735 2091
rect 12357 2057 12391 2091
rect 12541 2057 12575 2091
rect 12817 2057 12851 2091
rect 13277 2057 13311 2091
rect 14565 2057 14599 2091
rect 16681 2057 16715 2091
rect 18153 2057 18187 2091
rect 3433 1989 3467 2023
rect 7297 1989 7331 2023
rect 9045 1921 9079 1955
rect 10977 1921 11011 1955
rect 1133 1853 1167 1887
rect 1225 1853 1259 1887
rect 1501 1853 1535 1887
rect 1961 1853 1995 1887
rect 2053 1853 2087 1887
rect 2513 1853 2547 1887
rect 2605 1853 2639 1887
rect 2697 1853 2731 1887
rect 2881 1853 2915 1887
rect 3341 1853 3375 1887
rect 3617 1853 3651 1887
rect 3893 1853 3927 1887
rect 5365 1853 5399 1887
rect 5632 1853 5666 1887
rect 7113 1853 7147 1887
rect 7205 1853 7239 1887
rect 7481 1853 7515 1887
rect 7757 1853 7791 1887
rect 8217 1853 8251 1887
rect 8493 1853 8527 1887
rect 8769 1853 8803 1887
rect 10609 1853 10643 1887
rect 12449 1853 12483 1887
rect 12909 1853 12943 1887
rect 13369 1853 13403 1887
rect 13645 1853 13679 1887
rect 13737 1853 13771 1887
rect 13829 1853 13863 1887
rect 14105 1853 14139 1887
rect 14473 1853 14507 1887
rect 14749 1853 14783 1887
rect 15025 1863 15059 1897
rect 15301 1853 15335 1887
rect 16773 1853 16807 1887
rect 19073 1853 19107 1887
rect 1593 1785 1627 1819
rect 4138 1785 4172 1819
rect 7849 1785 7883 1819
rect 8125 1785 8159 1819
rect 9290 1785 9324 1819
rect 11244 1785 11278 1819
rect 15568 1785 15602 1819
rect 17018 1785 17052 1819
rect 1041 1717 1075 1751
rect 2145 1717 2179 1751
rect 2421 1717 2455 1751
rect 3709 1717 3743 1751
rect 5273 1717 5307 1751
rect 6745 1717 6779 1751
rect 8861 1717 8895 1751
rect 13921 1717 13955 1751
rect 14197 1717 14231 1751
rect 14841 1717 14875 1751
rect 15117 1717 15151 1751
rect 1501 1513 1535 1547
rect 3065 1513 3099 1547
rect 4813 1513 4847 1547
rect 4997 1513 5031 1547
rect 5273 1513 5307 1547
rect 5917 1513 5951 1547
rect 6469 1513 6503 1547
rect 8309 1513 8343 1547
rect 9781 1513 9815 1547
rect 10425 1513 10459 1547
rect 11069 1513 11103 1547
rect 11897 1513 11931 1547
rect 13277 1513 13311 1547
rect 14841 1513 14875 1547
rect 15301 1513 15335 1547
rect 15577 1513 15611 1547
rect 16221 1513 16255 1547
rect 17877 1513 17911 1547
rect 1930 1445 1964 1479
rect 3678 1445 3712 1479
rect 6193 1445 6227 1479
rect 8646 1445 8680 1479
rect 9965 1445 9999 1479
rect 1409 1377 1443 1411
rect 3157 1377 3191 1411
rect 5089 1377 5123 1411
rect 5181 1377 5215 1411
rect 5457 1377 5491 1411
rect 6009 1377 6043 1411
rect 6101 1377 6135 1411
rect 6377 1377 6411 1411
rect 6653 1377 6687 1411
rect 6745 1377 6779 1411
rect 7196 1377 7230 1411
rect 10057 1377 10091 1411
rect 10517 1377 10551 1411
rect 10609 1377 10643 1411
rect 10977 1377 11011 1411
rect 11253 1377 11287 1411
rect 11345 1377 11379 1411
rect 11529 1377 11563 1411
rect 11621 1377 11655 1411
rect 11989 1377 12023 1411
rect 12173 1377 12207 1411
rect 12265 1377 12299 1411
rect 12357 1377 12391 1411
rect 12633 1377 12667 1411
rect 12909 1377 12943 1411
rect 13185 1377 13219 1411
rect 13461 1377 13495 1411
rect 13717 1377 13751 1411
rect 14933 1377 14967 1411
rect 15393 1377 15427 1411
rect 15669 1377 15703 1411
rect 15761 1377 15795 1411
rect 15853 1377 15887 1411
rect 16313 1377 16347 1411
rect 16497 1377 16531 1411
rect 16753 1377 16787 1411
rect 1685 1309 1719 1343
rect 3249 1309 3283 1343
rect 3433 1309 3467 1343
rect 5549 1309 5583 1343
rect 6929 1309 6963 1343
rect 8401 1309 8435 1343
rect 10701 1309 10735 1343
rect 12725 1309 12759 1343
rect 12449 1241 12483 1275
rect 13001 1241 13035 1275
rect 15025 1173 15059 1207
rect 2237 969 2271 1003
rect 4169 969 4203 1003
rect 7205 969 7239 1003
rect 10609 969 10643 1003
rect 13185 969 13219 1003
rect 13645 969 13679 1003
rect 13921 969 13955 1003
rect 14197 969 14231 1003
rect 14473 969 14507 1003
rect 15669 969 15703 1003
rect 16221 969 16255 1003
rect 16497 969 16531 1003
rect 2421 901 2455 935
rect 11989 901 12023 935
rect 12909 901 12943 935
rect 857 765 891 799
rect 1409 765 1443 799
rect 2329 765 2363 799
rect 4077 765 4111 799
rect 7297 765 7331 799
rect 10425 765 10459 799
rect 13737 765 13771 799
rect 13829 765 13863 799
rect 14289 765 14323 799
rect 14381 765 14415 799
rect 15761 765 15795 799
rect 16129 765 16163 799
rect 16589 765 16623 799
rect 18521 765 18555 799
rect 19073 765 19107 799
rect 11805 697 11839 731
rect 12725 697 12759 731
rect 13093 697 13127 731
<< metal1 >>
rect 552 19066 19571 19088
rect 552 19014 5112 19066
rect 5164 19014 5176 19066
rect 5228 19014 5240 19066
rect 5292 19014 5304 19066
rect 5356 19014 5368 19066
rect 5420 19014 9827 19066
rect 9879 19014 9891 19066
rect 9943 19014 9955 19066
rect 10007 19014 10019 19066
rect 10071 19014 10083 19066
rect 10135 19014 14542 19066
rect 14594 19014 14606 19066
rect 14658 19014 14670 19066
rect 14722 19014 14734 19066
rect 14786 19014 14798 19066
rect 14850 19014 19257 19066
rect 19309 19014 19321 19066
rect 19373 19014 19385 19066
rect 19437 19014 19449 19066
rect 19501 19014 19513 19066
rect 19565 19014 19571 19066
rect 552 18992 19571 19014
rect 13173 18955 13231 18961
rect 13173 18921 13185 18955
rect 13219 18952 13231 18955
rect 13538 18952 13544 18964
rect 13219 18924 13544 18952
rect 13219 18921 13231 18924
rect 13173 18915 13231 18921
rect 13538 18912 13544 18924
rect 13596 18952 13602 18964
rect 14185 18955 14243 18961
rect 14185 18952 14197 18955
rect 13596 18924 14197 18952
rect 13596 18912 13602 18924
rect 14185 18921 14197 18924
rect 14231 18952 14243 18955
rect 15378 18952 15384 18964
rect 14231 18924 15384 18952
rect 14231 18921 14243 18924
rect 14185 18915 14243 18921
rect 15378 18912 15384 18924
rect 15436 18912 15442 18964
rect 10410 18844 10416 18896
rect 10468 18884 10474 18896
rect 12897 18887 12955 18893
rect 12897 18884 12909 18887
rect 10468 18856 12909 18884
rect 10468 18844 10474 18856
rect 12897 18853 12909 18856
rect 12943 18884 12955 18887
rect 12943 18856 13768 18884
rect 12943 18853 12955 18856
rect 12897 18847 12955 18853
rect 750 18776 756 18828
rect 808 18816 814 18828
rect 1397 18819 1455 18825
rect 1397 18816 1409 18819
rect 808 18788 1409 18816
rect 808 18776 814 18788
rect 1397 18785 1409 18788
rect 1443 18785 1455 18819
rect 1397 18779 1455 18785
rect 11425 18819 11483 18825
rect 11425 18785 11437 18819
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 11517 18819 11575 18825
rect 11517 18785 11529 18819
rect 11563 18816 11575 18819
rect 11974 18816 11980 18828
rect 11563 18788 11980 18816
rect 11563 18785 11575 18788
rect 11517 18779 11575 18785
rect 1118 18708 1124 18760
rect 1176 18708 1182 18760
rect 11440 18624 11468 18779
rect 11974 18776 11980 18788
rect 12032 18816 12038 18828
rect 12069 18819 12127 18825
rect 12069 18816 12081 18819
rect 12032 18788 12081 18816
rect 12032 18776 12038 18788
rect 12069 18785 12081 18788
rect 12115 18816 12127 18819
rect 12529 18819 12587 18825
rect 12529 18816 12541 18819
rect 12115 18788 12541 18816
rect 12115 18785 12127 18788
rect 12069 18779 12127 18785
rect 12529 18785 12541 18788
rect 12575 18785 12587 18819
rect 12529 18779 12587 18785
rect 12986 18776 12992 18828
rect 13044 18776 13050 18828
rect 13740 18825 13768 18856
rect 13081 18819 13139 18825
rect 13081 18785 13093 18819
rect 13127 18785 13139 18819
rect 13081 18779 13139 18785
rect 13725 18819 13783 18825
rect 13725 18785 13737 18819
rect 13771 18816 13783 18819
rect 13817 18819 13875 18825
rect 13817 18816 13829 18819
rect 13771 18788 13829 18816
rect 13771 18785 13783 18788
rect 13725 18779 13783 18785
rect 13817 18785 13829 18788
rect 13863 18785 13875 18819
rect 13817 18779 13875 18785
rect 14093 18819 14151 18825
rect 14093 18785 14105 18819
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 13096 18748 13124 18779
rect 13998 18748 14004 18760
rect 12544 18720 13124 18748
rect 13648 18720 14004 18748
rect 12544 18624 12572 18720
rect 842 18572 848 18624
rect 900 18572 906 18624
rect 11422 18572 11428 18624
rect 11480 18572 11486 18624
rect 12161 18615 12219 18621
rect 12161 18581 12173 18615
rect 12207 18612 12219 18615
rect 12526 18612 12532 18624
rect 12207 18584 12532 18612
rect 12207 18581 12219 18584
rect 12161 18575 12219 18581
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 13648 18621 13676 18720
rect 13998 18708 14004 18720
rect 14056 18748 14062 18760
rect 14108 18748 14136 18779
rect 14182 18776 14188 18828
rect 14240 18816 14246 18828
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 14240 18788 14381 18816
rect 14240 18776 14246 18788
rect 14369 18785 14381 18788
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 18506 18776 18512 18828
rect 18564 18776 18570 18828
rect 14056 18720 14136 18748
rect 14056 18708 14062 18720
rect 12621 18615 12679 18621
rect 12621 18581 12633 18615
rect 12667 18612 12679 18615
rect 13633 18615 13691 18621
rect 13633 18612 13645 18615
rect 12667 18584 13645 18612
rect 12667 18581 12679 18584
rect 12621 18575 12679 18581
rect 13633 18581 13645 18584
rect 13679 18581 13691 18615
rect 13633 18575 13691 18581
rect 13906 18572 13912 18624
rect 13964 18572 13970 18624
rect 14366 18572 14372 18624
rect 14424 18612 14430 18624
rect 14461 18615 14519 18621
rect 14461 18612 14473 18615
rect 14424 18584 14473 18612
rect 14424 18572 14430 18584
rect 14461 18581 14473 18584
rect 14507 18581 14519 18615
rect 14461 18575 14519 18581
rect 19058 18572 19064 18624
rect 19116 18572 19122 18624
rect 552 18522 19412 18544
rect 552 18470 2755 18522
rect 2807 18470 2819 18522
rect 2871 18470 2883 18522
rect 2935 18470 2947 18522
rect 2999 18470 3011 18522
rect 3063 18470 7470 18522
rect 7522 18470 7534 18522
rect 7586 18470 7598 18522
rect 7650 18470 7662 18522
rect 7714 18470 7726 18522
rect 7778 18470 12185 18522
rect 12237 18470 12249 18522
rect 12301 18470 12313 18522
rect 12365 18470 12377 18522
rect 12429 18470 12441 18522
rect 12493 18470 16900 18522
rect 16952 18470 16964 18522
rect 17016 18470 17028 18522
rect 17080 18470 17092 18522
rect 17144 18470 17156 18522
rect 17208 18470 19412 18522
rect 552 18448 19412 18470
rect 10410 18368 10416 18420
rect 10468 18368 10474 18420
rect 10502 18368 10508 18420
rect 10560 18408 10566 18420
rect 11422 18408 11428 18420
rect 10560 18380 11428 18408
rect 10560 18368 10566 18380
rect 11422 18368 11428 18380
rect 11480 18408 11486 18420
rect 11977 18411 12035 18417
rect 11977 18408 11989 18411
rect 11480 18380 11989 18408
rect 11480 18368 11486 18380
rect 11977 18377 11989 18380
rect 12023 18377 12035 18411
rect 11977 18371 12035 18377
rect 12526 18368 12532 18420
rect 12584 18368 12590 18420
rect 10428 18340 10456 18368
rect 11701 18343 11759 18349
rect 11701 18340 11713 18343
rect 10244 18312 10456 18340
rect 10520 18312 11713 18340
rect 2406 18232 2412 18284
rect 2464 18272 2470 18284
rect 3237 18275 3295 18281
rect 3237 18272 3249 18275
rect 2464 18244 3249 18272
rect 2464 18232 2470 18244
rect 3237 18241 3249 18244
rect 3283 18241 3295 18275
rect 3237 18235 3295 18241
rect 842 18164 848 18216
rect 900 18164 906 18216
rect 2682 18164 2688 18216
rect 2740 18164 2746 18216
rect 3053 18207 3111 18213
rect 3053 18173 3065 18207
rect 3099 18173 3111 18207
rect 3252 18204 3280 18235
rect 4709 18207 4767 18213
rect 4709 18204 4721 18207
rect 3252 18176 4721 18204
rect 3053 18167 3111 18173
rect 3068 18136 3096 18167
rect 4172 18148 4200 18176
rect 4709 18173 4721 18176
rect 4755 18173 4767 18207
rect 4709 18167 4767 18173
rect 4976 18207 5034 18213
rect 4976 18173 4988 18207
rect 5022 18204 5034 18207
rect 7561 18207 7619 18213
rect 5022 18176 7236 18204
rect 5022 18173 5034 18176
rect 4976 18167 5034 18173
rect 3504 18139 3562 18145
rect 3504 18136 3516 18139
rect 3068 18108 3516 18136
rect 3504 18105 3516 18108
rect 3550 18136 3562 18139
rect 3786 18136 3792 18148
rect 3550 18108 3792 18136
rect 3550 18105 3562 18108
rect 3504 18099 3562 18105
rect 3786 18096 3792 18108
rect 3844 18096 3850 18148
rect 4154 18096 4160 18148
rect 4212 18096 4218 18148
rect 2590 18028 2596 18080
rect 2648 18068 2654 18080
rect 2961 18071 3019 18077
rect 2961 18068 2973 18071
rect 2648 18040 2973 18068
rect 2648 18028 2654 18040
rect 2961 18037 2973 18040
rect 3007 18037 3019 18071
rect 2961 18031 3019 18037
rect 4617 18071 4675 18077
rect 4617 18037 4629 18071
rect 4663 18068 4675 18071
rect 5718 18068 5724 18080
rect 4663 18040 5724 18068
rect 4663 18037 4675 18040
rect 4617 18031 4675 18037
rect 5718 18028 5724 18040
rect 5776 18028 5782 18080
rect 6086 18028 6092 18080
rect 6144 18028 6150 18080
rect 6181 18071 6239 18077
rect 6181 18037 6193 18071
rect 6227 18068 6239 18071
rect 6270 18068 6276 18080
rect 6227 18040 6276 18068
rect 6227 18037 6239 18040
rect 6181 18031 6239 18037
rect 6270 18028 6276 18040
rect 6328 18028 6334 18080
rect 7208 18068 7236 18176
rect 7561 18173 7573 18207
rect 7607 18204 7619 18207
rect 8386 18204 8392 18216
rect 7607 18176 8392 18204
rect 7607 18173 7619 18176
rect 7561 18167 7619 18173
rect 8386 18164 8392 18176
rect 8444 18204 8450 18216
rect 8849 18207 8907 18213
rect 8849 18204 8861 18207
rect 8444 18176 8861 18204
rect 8444 18164 8450 18176
rect 8849 18173 8861 18176
rect 8895 18173 8907 18207
rect 8849 18167 8907 18173
rect 9116 18207 9174 18213
rect 9116 18173 9128 18207
rect 9162 18204 9174 18207
rect 10244 18204 10272 18312
rect 9162 18176 10272 18204
rect 9162 18173 9174 18176
rect 9116 18167 9174 18173
rect 10318 18164 10324 18216
rect 10376 18164 10382 18216
rect 10520 18204 10548 18312
rect 11701 18309 11713 18312
rect 11747 18340 11759 18343
rect 11747 18312 12388 18340
rect 11747 18309 11759 18312
rect 11701 18303 11759 18309
rect 11057 18275 11115 18281
rect 11057 18241 11069 18275
rect 11103 18272 11115 18275
rect 11103 18244 11836 18272
rect 11103 18241 11115 18244
rect 11057 18235 11115 18241
rect 11808 18216 11836 18244
rect 10965 18207 11023 18213
rect 10965 18204 10977 18207
rect 10428 18176 10548 18204
rect 10704 18176 10977 18204
rect 7316 18139 7374 18145
rect 7316 18105 7328 18139
rect 7362 18136 7374 18139
rect 8478 18136 8484 18148
rect 7362 18108 8484 18136
rect 7362 18105 7374 18108
rect 7316 18099 7374 18105
rect 8478 18096 8484 18108
rect 8536 18136 8542 18148
rect 10428 18136 10456 18176
rect 8536 18108 10456 18136
rect 8536 18096 8542 18108
rect 10704 18080 10732 18176
rect 10965 18173 10977 18176
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 11333 18207 11391 18213
rect 11333 18173 11345 18207
rect 11379 18173 11391 18207
rect 11333 18167 11391 18173
rect 11348 18080 11376 18167
rect 11790 18164 11796 18216
rect 11848 18164 11854 18216
rect 12360 18213 12388 18312
rect 12544 18272 12572 18368
rect 12544 18244 13032 18272
rect 13004 18213 13032 18244
rect 12069 18207 12127 18213
rect 12069 18173 12081 18207
rect 12115 18173 12127 18207
rect 12345 18207 12403 18213
rect 12345 18204 12357 18207
rect 12303 18176 12357 18204
rect 12069 18167 12127 18173
rect 12345 18173 12357 18176
rect 12391 18204 12403 18207
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12391 18176 12449 18204
rect 12391 18173 12403 18176
rect 12345 18167 12403 18173
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12713 18207 12771 18213
rect 12713 18173 12725 18207
rect 12759 18173 12771 18207
rect 12713 18167 12771 18173
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18173 13047 18207
rect 12989 18167 13047 18173
rect 11425 18139 11483 18145
rect 11425 18105 11437 18139
rect 11471 18136 11483 18139
rect 12084 18136 12112 18167
rect 12253 18139 12311 18145
rect 12253 18136 12265 18139
rect 11471 18108 12265 18136
rect 11471 18105 11483 18108
rect 11425 18099 11483 18105
rect 12253 18105 12265 18108
rect 12299 18136 12311 18139
rect 12728 18136 12756 18167
rect 14458 18164 14464 18216
rect 14516 18204 14522 18216
rect 15105 18207 15163 18213
rect 15105 18204 15117 18207
rect 14516 18176 15117 18204
rect 14516 18164 14522 18176
rect 15105 18173 15117 18176
rect 15151 18173 15163 18207
rect 15105 18167 15163 18173
rect 15197 18207 15255 18213
rect 15197 18173 15209 18207
rect 15243 18204 15255 18207
rect 15286 18204 15292 18216
rect 15243 18176 15292 18204
rect 15243 18173 15255 18176
rect 15197 18167 15255 18173
rect 15286 18164 15292 18176
rect 15344 18164 15350 18216
rect 15464 18207 15522 18213
rect 15464 18173 15476 18207
rect 15510 18173 15522 18207
rect 18046 18204 18052 18216
rect 15464 18167 15522 18173
rect 16500 18176 18052 18204
rect 12299 18108 12756 18136
rect 12299 18105 12311 18108
rect 12253 18099 12311 18105
rect 13906 18096 13912 18148
rect 13964 18136 13970 18148
rect 14826 18136 14832 18148
rect 14884 18145 14890 18148
rect 14884 18139 14907 18145
rect 13964 18108 14832 18136
rect 13964 18096 13970 18108
rect 14826 18096 14832 18108
rect 14895 18105 14907 18139
rect 14884 18099 14907 18105
rect 14884 18096 14890 18099
rect 9582 18068 9588 18080
rect 7208 18040 9588 18068
rect 9582 18028 9588 18040
rect 9640 18068 9646 18080
rect 10134 18068 10140 18080
rect 9640 18040 10140 18068
rect 9640 18028 9646 18040
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10226 18028 10232 18080
rect 10284 18028 10290 18080
rect 10686 18028 10692 18080
rect 10744 18028 10750 18080
rect 11330 18028 11336 18080
rect 11388 18028 11394 18080
rect 12805 18071 12863 18077
rect 12805 18037 12817 18071
rect 12851 18068 12863 18071
rect 12986 18068 12992 18080
rect 12851 18040 12992 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 12986 18028 12992 18040
rect 13044 18068 13050 18080
rect 13081 18071 13139 18077
rect 13081 18068 13093 18071
rect 13044 18040 13093 18068
rect 13044 18028 13050 18040
rect 13081 18037 13093 18040
rect 13127 18068 13139 18071
rect 13354 18068 13360 18080
rect 13127 18040 13360 18068
rect 13127 18037 13139 18040
rect 13081 18031 13139 18037
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 13722 18028 13728 18080
rect 13780 18028 13786 18080
rect 15304 18068 15332 18164
rect 15378 18096 15384 18148
rect 15436 18136 15442 18148
rect 15488 18136 15516 18167
rect 15436 18108 15516 18136
rect 15436 18096 15442 18108
rect 16500 18068 16528 18176
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 19058 18164 19064 18216
rect 19116 18164 19122 18216
rect 17804 18139 17862 18145
rect 17804 18105 17816 18139
rect 17850 18136 17862 18139
rect 18230 18136 18236 18148
rect 17850 18108 18236 18136
rect 17850 18105 17862 18108
rect 17804 18099 17862 18105
rect 18230 18096 18236 18108
rect 18288 18096 18294 18148
rect 15304 18040 16528 18068
rect 16574 18028 16580 18080
rect 16632 18028 16638 18080
rect 16666 18028 16672 18080
rect 16724 18028 16730 18080
rect 552 17978 19571 18000
rect 552 17926 5112 17978
rect 5164 17926 5176 17978
rect 5228 17926 5240 17978
rect 5292 17926 5304 17978
rect 5356 17926 5368 17978
rect 5420 17926 9827 17978
rect 9879 17926 9891 17978
rect 9943 17926 9955 17978
rect 10007 17926 10019 17978
rect 10071 17926 10083 17978
rect 10135 17926 14542 17978
rect 14594 17926 14606 17978
rect 14658 17926 14670 17978
rect 14722 17926 14734 17978
rect 14786 17926 14798 17978
rect 14850 17926 19257 17978
rect 19309 17926 19321 17978
rect 19373 17926 19385 17978
rect 19437 17926 19449 17978
rect 19501 17926 19513 17978
rect 19565 17926 19571 17978
rect 552 17904 19571 17926
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 9858 17864 9864 17876
rect 4396 17836 9864 17864
rect 4396 17824 4402 17836
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 9968 17836 11100 17864
rect 2590 17796 2596 17808
rect 2056 17768 2596 17796
rect 2056 17737 2084 17768
rect 2590 17756 2596 17768
rect 2648 17805 2654 17808
rect 2648 17799 2712 17805
rect 2648 17765 2666 17799
rect 2700 17765 2712 17799
rect 2648 17759 2712 17765
rect 4080 17768 4292 17796
rect 2648 17756 2654 17759
rect 2041 17731 2099 17737
rect 2041 17728 2053 17731
rect 1504 17700 2053 17728
rect 1504 17672 1532 17700
rect 2041 17697 2053 17700
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 2314 17688 2320 17740
rect 2372 17688 2378 17740
rect 4080 17737 4108 17768
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17697 4123 17731
rect 4065 17691 4123 17697
rect 4154 17688 4160 17740
rect 4212 17688 4218 17740
rect 4264 17728 4292 17768
rect 6270 17756 6276 17808
rect 6328 17796 6334 17808
rect 6457 17799 6515 17805
rect 6457 17796 6469 17799
rect 6328 17768 6469 17796
rect 6328 17756 6334 17768
rect 6457 17765 6469 17768
rect 6503 17765 6515 17799
rect 6457 17759 6515 17765
rect 9398 17756 9404 17808
rect 9456 17796 9462 17808
rect 9968 17796 9996 17836
rect 9456 17768 9996 17796
rect 9456 17756 9462 17768
rect 4430 17737 4436 17740
rect 4424 17728 4436 17737
rect 4264 17700 4436 17728
rect 4424 17691 4436 17700
rect 4430 17688 4436 17691
rect 4488 17688 4494 17740
rect 6181 17731 6239 17737
rect 6181 17728 6193 17731
rect 5552 17700 6193 17728
rect 1486 17620 1492 17672
rect 1544 17620 1550 17672
rect 1578 17620 1584 17672
rect 1636 17660 1642 17672
rect 2406 17660 2412 17672
rect 1636 17632 2412 17660
rect 1636 17620 1642 17632
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 5552 17601 5580 17700
rect 6181 17697 6193 17700
rect 6227 17697 6239 17731
rect 6365 17731 6423 17737
rect 6365 17728 6377 17731
rect 6181 17691 6239 17697
rect 6288 17700 6377 17728
rect 6288 17604 6316 17700
rect 6365 17697 6377 17700
rect 6411 17697 6423 17731
rect 6365 17691 6423 17697
rect 6546 17688 6552 17740
rect 6604 17688 6610 17740
rect 7949 17731 8007 17737
rect 7949 17697 7961 17731
rect 7995 17728 8007 17731
rect 8110 17728 8116 17740
rect 7995 17700 8116 17728
rect 7995 17697 8007 17700
rect 7949 17691 8007 17697
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 8205 17731 8263 17737
rect 8205 17697 8217 17731
rect 8251 17728 8263 17731
rect 8297 17731 8355 17737
rect 8297 17728 8309 17731
rect 8251 17700 8309 17728
rect 8251 17697 8263 17700
rect 8205 17691 8263 17697
rect 8297 17697 8309 17700
rect 8343 17728 8355 17731
rect 8386 17728 8392 17740
rect 8343 17700 8392 17728
rect 8343 17697 8355 17700
rect 8297 17691 8355 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 8564 17731 8622 17737
rect 8564 17697 8576 17731
rect 8610 17728 8622 17731
rect 9674 17728 9680 17740
rect 8610 17700 9680 17728
rect 8610 17697 8622 17700
rect 8564 17691 8622 17697
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 9968 17737 9996 17768
rect 10045 17799 10103 17805
rect 10045 17765 10057 17799
rect 10091 17796 10103 17799
rect 10226 17796 10232 17808
rect 10091 17768 10232 17796
rect 10091 17765 10103 17768
rect 10045 17759 10103 17765
rect 10226 17756 10232 17768
rect 10284 17756 10290 17808
rect 11072 17796 11100 17836
rect 11238 17824 11244 17876
rect 11296 17864 11302 17876
rect 13722 17864 13728 17876
rect 11296 17836 13728 17864
rect 11296 17824 11302 17836
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 13906 17824 13912 17876
rect 13964 17864 13970 17876
rect 14369 17867 14427 17873
rect 14369 17864 14381 17867
rect 13964 17836 14381 17864
rect 13964 17824 13970 17836
rect 14369 17833 14381 17836
rect 14415 17833 14427 17867
rect 14369 17827 14427 17833
rect 18230 17824 18236 17876
rect 18288 17864 18294 17876
rect 18288 17836 18644 17864
rect 18288 17824 18294 17836
rect 16485 17799 16543 17805
rect 16485 17796 16497 17799
rect 10612 17768 11008 17796
rect 11072 17768 16497 17796
rect 9953 17731 10011 17737
rect 9953 17697 9965 17731
rect 9999 17697 10011 17731
rect 9953 17691 10011 17697
rect 10134 17688 10140 17740
rect 10192 17688 10198 17740
rect 10321 17731 10379 17737
rect 10321 17697 10333 17731
rect 10367 17697 10379 17731
rect 10321 17691 10379 17697
rect 10336 17660 10364 17691
rect 9600 17632 10364 17660
rect 3789 17595 3847 17601
rect 3789 17561 3801 17595
rect 3835 17592 3847 17595
rect 5537 17595 5595 17601
rect 3835 17564 4200 17592
rect 3835 17561 3847 17564
rect 3789 17555 3847 17561
rect 1854 17484 1860 17536
rect 1912 17524 1918 17536
rect 1949 17527 2007 17533
rect 1949 17524 1961 17527
rect 1912 17496 1961 17524
rect 1912 17484 1918 17496
rect 1949 17493 1961 17496
rect 1995 17493 2007 17527
rect 1949 17487 2007 17493
rect 2222 17484 2228 17536
rect 2280 17484 2286 17536
rect 3973 17527 4031 17533
rect 3973 17493 3985 17527
rect 4019 17524 4031 17527
rect 4062 17524 4068 17536
rect 4019 17496 4068 17524
rect 4019 17493 4031 17496
rect 3973 17487 4031 17493
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 4172 17524 4200 17564
rect 5537 17561 5549 17595
rect 5583 17561 5595 17595
rect 5537 17555 5595 17561
rect 6270 17552 6276 17604
rect 6328 17552 6334 17604
rect 6656 17564 7328 17592
rect 6656 17524 6684 17564
rect 4172 17496 6684 17524
rect 6730 17484 6736 17536
rect 6788 17484 6794 17536
rect 6822 17484 6828 17536
rect 6880 17484 6886 17536
rect 7300 17524 7328 17564
rect 9600 17524 9628 17632
rect 10318 17592 10324 17604
rect 9692 17564 10324 17592
rect 9692 17533 9720 17564
rect 10318 17552 10324 17564
rect 10376 17552 10382 17604
rect 7300 17496 9628 17524
rect 9677 17527 9735 17533
rect 9677 17493 9689 17527
rect 9723 17493 9735 17527
rect 9677 17487 9735 17493
rect 9766 17484 9772 17536
rect 9824 17484 9830 17536
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 10612 17524 10640 17768
rect 10980 17737 11008 17768
rect 10781 17731 10839 17737
rect 10781 17697 10793 17731
rect 10827 17697 10839 17731
rect 10781 17691 10839 17697
rect 10965 17731 11023 17737
rect 10965 17697 10977 17731
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 10796 17592 10824 17691
rect 11146 17688 11152 17740
rect 11204 17688 11210 17740
rect 11238 17688 11244 17740
rect 11296 17688 11302 17740
rect 11348 17737 11376 17768
rect 16485 17765 16497 17768
rect 16531 17765 16543 17799
rect 16485 17759 16543 17765
rect 18046 17756 18052 17808
rect 18104 17796 18110 17808
rect 18104 17768 18552 17796
rect 18104 17756 18110 17768
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17697 11391 17731
rect 11333 17691 11391 17697
rect 11609 17731 11667 17737
rect 11609 17697 11621 17731
rect 11655 17728 11667 17731
rect 11882 17728 11888 17740
rect 11655 17700 11888 17728
rect 11655 17697 11667 17700
rect 11609 17691 11667 17697
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 12526 17688 12532 17740
rect 12584 17728 12590 17740
rect 12998 17731 13056 17737
rect 12998 17728 13010 17731
rect 12584 17700 13010 17728
rect 12584 17688 12590 17700
rect 12998 17697 13010 17700
rect 13044 17697 13056 17731
rect 12998 17691 13056 17697
rect 13354 17688 13360 17740
rect 13412 17688 13418 17740
rect 13449 17731 13507 17737
rect 13449 17697 13461 17731
rect 13495 17728 13507 17731
rect 13722 17728 13728 17740
rect 13495 17700 13728 17728
rect 13495 17697 13507 17700
rect 13449 17691 13507 17697
rect 13722 17688 13728 17700
rect 13780 17688 13786 17740
rect 13998 17688 14004 17740
rect 14056 17688 14062 17740
rect 14274 17688 14280 17740
rect 14332 17688 14338 17740
rect 14366 17688 14372 17740
rect 14424 17728 14430 17740
rect 14809 17731 14867 17737
rect 14809 17728 14821 17731
rect 14424 17700 14821 17728
rect 14424 17688 14430 17700
rect 14809 17697 14821 17700
rect 14855 17728 14867 17731
rect 15102 17728 15108 17740
rect 14855 17700 15108 17728
rect 14855 17697 14867 17700
rect 14809 17691 14867 17697
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 16298 17688 16304 17740
rect 16356 17688 16362 17740
rect 16393 17731 16451 17737
rect 16393 17697 16405 17731
rect 16439 17697 16451 17731
rect 16393 17691 16451 17697
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17660 13323 17663
rect 14458 17660 14464 17672
rect 13311 17632 14464 17660
rect 13311 17629 13323 17632
rect 13265 17623 13323 17629
rect 14458 17620 14464 17632
rect 14516 17660 14522 17672
rect 14553 17663 14611 17669
rect 14553 17660 14565 17663
rect 14516 17632 14565 17660
rect 14516 17620 14522 17632
rect 14553 17629 14565 17632
rect 14599 17629 14611 17663
rect 16408 17660 16436 17691
rect 16574 17688 16580 17740
rect 16632 17728 16638 17740
rect 18524 17737 18552 17768
rect 18616 17737 18644 17836
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 16632 17700 16681 17728
rect 16632 17688 16638 17700
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 17037 17731 17095 17737
rect 17037 17697 17049 17731
rect 17083 17728 17095 17731
rect 18253 17731 18311 17737
rect 18253 17728 18265 17731
rect 17083 17700 18265 17728
rect 17083 17697 17095 17700
rect 17037 17691 17095 17697
rect 18253 17697 18265 17700
rect 18299 17728 18311 17731
rect 18509 17731 18567 17737
rect 18299 17700 18460 17728
rect 18299 17697 18311 17700
rect 18253 17691 18311 17697
rect 18432 17660 18460 17700
rect 18509 17697 18521 17731
rect 18555 17697 18567 17731
rect 18509 17691 18567 17697
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17697 18659 17731
rect 18601 17691 18659 17697
rect 18782 17688 18788 17740
rect 18840 17688 18846 17740
rect 18800 17660 18828 17688
rect 16408 17632 16712 17660
rect 18432 17632 18828 17660
rect 14553 17623 14611 17629
rect 16684 17604 16712 17632
rect 11422 17592 11428 17604
rect 10796 17564 11428 17592
rect 11422 17552 11428 17564
rect 11480 17592 11486 17604
rect 11701 17595 11759 17601
rect 11701 17592 11713 17595
rect 11480 17564 11713 17592
rect 11480 17552 11486 17564
rect 11701 17561 11713 17564
rect 11747 17561 11759 17595
rect 11701 17555 11759 17561
rect 14093 17595 14151 17601
rect 14093 17561 14105 17595
rect 14139 17592 14151 17595
rect 14182 17592 14188 17604
rect 14139 17564 14188 17592
rect 14139 17561 14151 17564
rect 14093 17555 14151 17561
rect 14182 17552 14188 17564
rect 14240 17552 14246 17604
rect 16298 17592 16304 17604
rect 15948 17564 16304 17592
rect 9916 17496 10640 17524
rect 9916 17484 9922 17496
rect 10686 17484 10692 17536
rect 10744 17484 10750 17536
rect 11514 17484 11520 17536
rect 11572 17484 11578 17536
rect 11885 17527 11943 17533
rect 11885 17493 11897 17527
rect 11931 17524 11943 17527
rect 12894 17524 12900 17536
rect 11931 17496 12900 17524
rect 11931 17493 11943 17496
rect 11885 17487 11943 17493
rect 12894 17484 12900 17496
rect 12952 17484 12958 17536
rect 13817 17527 13875 17533
rect 13817 17493 13829 17527
rect 13863 17524 13875 17527
rect 14550 17524 14556 17536
rect 13863 17496 14556 17524
rect 13863 17493 13875 17496
rect 13817 17487 13875 17493
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 15948 17533 15976 17564
rect 16298 17552 16304 17564
rect 16356 17552 16362 17604
rect 16666 17552 16672 17604
rect 16724 17552 16730 17604
rect 15933 17527 15991 17533
rect 15933 17493 15945 17527
rect 15979 17493 15991 17527
rect 15933 17487 15991 17493
rect 16114 17484 16120 17536
rect 16172 17484 16178 17536
rect 16758 17484 16764 17536
rect 16816 17524 16822 17536
rect 16945 17527 17003 17533
rect 16945 17524 16957 17527
rect 16816 17496 16957 17524
rect 16816 17484 16822 17496
rect 16945 17493 16957 17496
rect 16991 17493 17003 17527
rect 16945 17487 17003 17493
rect 17129 17527 17187 17533
rect 17129 17493 17141 17527
rect 17175 17524 17187 17527
rect 17218 17524 17224 17536
rect 17175 17496 17224 17524
rect 17175 17493 17187 17496
rect 17129 17487 17187 17493
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 18690 17484 18696 17536
rect 18748 17484 18754 17536
rect 552 17434 19412 17456
rect 552 17382 2755 17434
rect 2807 17382 2819 17434
rect 2871 17382 2883 17434
rect 2935 17382 2947 17434
rect 2999 17382 3011 17434
rect 3063 17382 7470 17434
rect 7522 17382 7534 17434
rect 7586 17382 7598 17434
rect 7650 17382 7662 17434
rect 7714 17382 7726 17434
rect 7778 17382 12185 17434
rect 12237 17382 12249 17434
rect 12301 17382 12313 17434
rect 12365 17382 12377 17434
rect 12429 17382 12441 17434
rect 12493 17382 16900 17434
rect 16952 17382 16964 17434
rect 17016 17382 17028 17434
rect 17080 17382 17092 17434
rect 17144 17382 17156 17434
rect 17208 17382 19412 17434
rect 552 17360 19412 17382
rect 1397 17323 1455 17329
rect 1397 17289 1409 17323
rect 1443 17320 1455 17323
rect 2222 17320 2228 17332
rect 1443 17292 2228 17320
rect 1443 17289 1455 17292
rect 1397 17283 1455 17289
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 2961 17323 3019 17329
rect 2961 17289 2973 17323
rect 3007 17320 3019 17323
rect 4338 17320 4344 17332
rect 3007 17292 4344 17320
rect 3007 17289 3019 17292
rect 2961 17283 3019 17289
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 4430 17280 4436 17332
rect 4488 17320 4494 17332
rect 4617 17323 4675 17329
rect 4617 17320 4629 17323
rect 4488 17292 4629 17320
rect 4488 17280 4494 17292
rect 4617 17289 4629 17292
rect 4663 17320 4675 17323
rect 4893 17323 4951 17329
rect 4893 17320 4905 17323
rect 4663 17292 4905 17320
rect 4663 17289 4675 17292
rect 4617 17283 4675 17289
rect 4893 17289 4905 17292
rect 4939 17289 4951 17323
rect 4893 17283 4951 17289
rect 6822 17280 6828 17332
rect 6880 17280 6886 17332
rect 8478 17280 8484 17332
rect 8536 17280 8542 17332
rect 9398 17280 9404 17332
rect 9456 17280 9462 17332
rect 9582 17280 9588 17332
rect 9640 17280 9646 17332
rect 10134 17280 10140 17332
rect 10192 17320 10198 17332
rect 11146 17320 11152 17332
rect 10192 17292 11152 17320
rect 10192 17280 10198 17292
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 11422 17280 11428 17332
rect 11480 17280 11486 17332
rect 11701 17323 11759 17329
rect 11701 17289 11713 17323
rect 11747 17320 11759 17323
rect 11790 17320 11796 17332
rect 11747 17292 11796 17320
rect 11747 17289 11759 17292
rect 11701 17283 11759 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 11974 17280 11980 17332
rect 12032 17280 12038 17332
rect 13633 17323 13691 17329
rect 13633 17289 13645 17323
rect 13679 17320 13691 17323
rect 13722 17320 13728 17332
rect 13679 17292 13728 17320
rect 13679 17289 13691 17292
rect 13633 17283 13691 17289
rect 13722 17280 13728 17292
rect 13780 17320 13786 17332
rect 14274 17320 14280 17332
rect 13780 17292 14280 17320
rect 13780 17280 13786 17292
rect 14274 17280 14280 17292
rect 14332 17280 14338 17332
rect 14550 17280 14556 17332
rect 14608 17280 14614 17332
rect 15102 17280 15108 17332
rect 15160 17320 15166 17332
rect 15473 17323 15531 17329
rect 15473 17320 15485 17323
rect 15160 17292 15485 17320
rect 15160 17280 15166 17292
rect 4448 17252 4476 17280
rect 3988 17224 4476 17252
rect 1578 17144 1584 17196
rect 1636 17144 1642 17196
rect 842 17076 848 17128
rect 900 17076 906 17128
rect 1486 17076 1492 17128
rect 1544 17076 1550 17128
rect 1854 17125 1860 17128
rect 1848 17116 1860 17125
rect 1815 17088 1860 17116
rect 1848 17079 1860 17088
rect 1854 17076 1860 17079
rect 1912 17076 1918 17128
rect 3513 17119 3571 17125
rect 3513 17085 3525 17119
rect 3559 17085 3571 17119
rect 3513 17079 3571 17085
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17116 3847 17119
rect 3988 17116 4016 17224
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 5537 17187 5595 17193
rect 5537 17184 5549 17187
rect 4212 17156 5549 17184
rect 4212 17144 4218 17156
rect 5537 17153 5549 17156
rect 5583 17153 5595 17187
rect 6840 17184 6868 17280
rect 6840 17156 7880 17184
rect 5537 17147 5595 17153
rect 3835 17088 4016 17116
rect 4065 17119 4123 17125
rect 3835 17085 3847 17088
rect 3789 17079 3847 17085
rect 4065 17085 4077 17119
rect 4111 17116 4123 17119
rect 4246 17116 4252 17128
rect 4111 17088 4252 17116
rect 4111 17085 4123 17088
rect 4065 17079 4123 17085
rect 3142 17048 3148 17060
rect 2746 17020 3148 17048
rect 2314 16940 2320 16992
rect 2372 16980 2378 16992
rect 2746 16980 2774 17020
rect 3142 17008 3148 17020
rect 3200 17048 3206 17060
rect 3421 17051 3479 17057
rect 3421 17048 3433 17051
rect 3200 17020 3433 17048
rect 3200 17008 3206 17020
rect 3421 17017 3433 17020
rect 3467 17017 3479 17051
rect 3528 17048 3556 17079
rect 4246 17076 4252 17088
rect 4304 17076 4310 17128
rect 4338 17076 4344 17128
rect 4396 17076 4402 17128
rect 4709 17119 4767 17125
rect 4709 17085 4721 17119
rect 4755 17085 4767 17119
rect 4709 17079 4767 17085
rect 3878 17048 3884 17060
rect 3528 17020 3884 17048
rect 3421 17011 3479 17017
rect 3878 17008 3884 17020
rect 3936 17008 3942 17060
rect 4724 17048 4752 17079
rect 4798 17076 4804 17128
rect 4856 17076 4862 17128
rect 7852 17125 7880 17156
rect 7944 17156 9260 17184
rect 7944 17128 7972 17156
rect 7561 17119 7619 17125
rect 7561 17116 7573 17119
rect 6932 17088 7573 17116
rect 4982 17048 4988 17060
rect 4724 17020 4988 17048
rect 4982 17008 4988 17020
rect 5040 17048 5046 17060
rect 5782 17051 5840 17057
rect 5782 17048 5794 17051
rect 5040 17020 5794 17048
rect 5040 17008 5046 17020
rect 5782 17017 5794 17020
rect 5828 17017 5840 17051
rect 5782 17011 5840 17017
rect 2372 16952 2774 16980
rect 2372 16940 2378 16952
rect 3694 16940 3700 16992
rect 3752 16940 3758 16992
rect 3786 16940 3792 16992
rect 3844 16980 3850 16992
rect 3973 16983 4031 16989
rect 3973 16980 3985 16983
rect 3844 16952 3985 16980
rect 3844 16940 3850 16952
rect 3973 16949 3985 16952
rect 4019 16949 4031 16983
rect 3973 16943 4031 16949
rect 4062 16940 4068 16992
rect 4120 16980 4126 16992
rect 6932 16989 6960 17088
rect 7561 17085 7573 17088
rect 7607 17085 7619 17119
rect 7561 17079 7619 17085
rect 7837 17119 7895 17125
rect 7837 17085 7849 17119
rect 7883 17085 7895 17119
rect 7837 17079 7895 17085
rect 7926 17076 7932 17128
rect 7984 17076 7990 17128
rect 8110 17076 8116 17128
rect 8168 17116 8174 17128
rect 9232 17125 9260 17156
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 10152 17184 10180 17280
rect 11808 17252 11836 17280
rect 13265 17255 13323 17261
rect 11808 17224 11928 17252
rect 11606 17184 11612 17196
rect 9364 17156 10180 17184
rect 11256 17156 11612 17184
rect 9364 17144 9370 17156
rect 8573 17119 8631 17125
rect 8573 17116 8585 17119
rect 8168 17088 8585 17116
rect 8168 17076 8174 17088
rect 8573 17085 8585 17088
rect 8619 17085 8631 17119
rect 8573 17079 8631 17085
rect 9217 17119 9275 17125
rect 9217 17085 9229 17119
rect 9263 17116 9275 17119
rect 9490 17116 9496 17128
rect 9263 17088 9496 17116
rect 9263 17085 9275 17088
rect 9217 17079 9275 17085
rect 7742 17008 7748 17060
rect 7800 17048 7806 17060
rect 8588 17048 8616 17079
rect 9490 17076 9496 17088
rect 9548 17076 9554 17128
rect 9582 17076 9588 17128
rect 9640 17116 9646 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 9640 17088 9689 17116
rect 9640 17076 9646 17088
rect 9677 17085 9689 17088
rect 9723 17116 9735 17119
rect 10686 17116 10692 17128
rect 9723 17088 10692 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 10686 17076 10692 17088
rect 10744 17076 10750 17128
rect 10781 17119 10839 17125
rect 10781 17085 10793 17119
rect 10827 17116 10839 17119
rect 10870 17116 10876 17128
rect 10827 17088 10876 17116
rect 10827 17085 10839 17088
rect 10781 17079 10839 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 11256 17125 11284 17156
rect 11606 17144 11612 17156
rect 11664 17184 11670 17196
rect 11664 17156 11836 17184
rect 11664 17144 11670 17156
rect 11149 17119 11207 17125
rect 11149 17085 11161 17119
rect 11195 17085 11207 17119
rect 11149 17079 11207 17085
rect 11241 17119 11299 17125
rect 11241 17085 11253 17119
rect 11287 17085 11299 17119
rect 11241 17079 11299 17085
rect 11054 17048 11060 17060
rect 7800 17020 8248 17048
rect 8588 17020 11060 17048
rect 7800 17008 7806 17020
rect 4249 16983 4307 16989
rect 4249 16980 4261 16983
rect 4120 16952 4261 16980
rect 4120 16940 4126 16952
rect 4249 16949 4261 16952
rect 4295 16949 4307 16983
rect 4249 16943 4307 16949
rect 6917 16983 6975 16989
rect 6917 16949 6929 16983
rect 6963 16949 6975 16983
rect 6917 16943 6975 16949
rect 8110 16940 8116 16992
rect 8168 16940 8174 16992
rect 8220 16980 8248 17020
rect 11054 17008 11060 17020
rect 11112 17048 11118 17060
rect 11164 17048 11192 17079
rect 11422 17076 11428 17128
rect 11480 17116 11486 17128
rect 11808 17125 11836 17156
rect 11900 17125 11928 17224
rect 13265 17221 13277 17255
rect 13311 17252 13323 17255
rect 14182 17252 14188 17264
rect 13311 17224 14188 17252
rect 13311 17221 13323 17224
rect 13265 17215 13323 17221
rect 14182 17212 14188 17224
rect 14240 17212 14246 17264
rect 13538 17144 13544 17196
rect 13596 17184 13602 17196
rect 13596 17156 13768 17184
rect 13596 17144 13602 17156
rect 13740 17125 13768 17156
rect 13906 17144 13912 17196
rect 13964 17144 13970 17196
rect 14200 17184 14228 17212
rect 14568 17184 14596 17280
rect 15102 17184 15108 17196
rect 14200 17156 14320 17184
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 11480 17088 11529 17116
rect 11480 17076 11486 17088
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 11793 17119 11851 17125
rect 11793 17085 11805 17119
rect 11839 17085 11851 17119
rect 11793 17079 11851 17085
rect 11885 17119 11943 17125
rect 11885 17085 11897 17119
rect 11931 17085 11943 17119
rect 11885 17079 11943 17085
rect 13357 17119 13415 17125
rect 13357 17085 13369 17119
rect 13403 17085 13415 17119
rect 13357 17079 13415 17085
rect 13725 17119 13783 17125
rect 13725 17085 13737 17119
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 13372 17048 13400 17079
rect 13924 17048 13952 17144
rect 14292 17125 14320 17156
rect 14568 17156 15108 17184
rect 14185 17119 14243 17125
rect 14185 17085 14197 17119
rect 14231 17085 14243 17119
rect 14185 17079 14243 17085
rect 14277 17119 14335 17125
rect 14277 17085 14289 17119
rect 14323 17085 14335 17119
rect 14568 17116 14596 17156
rect 15102 17144 15108 17156
rect 15160 17184 15166 17196
rect 15197 17187 15255 17193
rect 15197 17184 15209 17187
rect 15160 17156 15209 17184
rect 15160 17144 15166 17156
rect 15197 17153 15209 17156
rect 15243 17153 15255 17187
rect 15197 17147 15255 17153
rect 14737 17119 14795 17125
rect 14737 17116 14749 17119
rect 14568 17088 14749 17116
rect 14277 17079 14335 17085
rect 14737 17085 14749 17088
rect 14783 17085 14795 17119
rect 14737 17079 14795 17085
rect 14829 17119 14887 17125
rect 14829 17085 14841 17119
rect 14875 17116 14887 17119
rect 14918 17116 14924 17128
rect 14875 17088 14924 17116
rect 14875 17085 14887 17088
rect 14829 17079 14887 17085
rect 11112 17020 11928 17048
rect 13372 17020 13952 17048
rect 14200 17048 14228 17079
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 15304 17125 15332 17292
rect 15473 17289 15485 17292
rect 15519 17320 15531 17323
rect 15562 17320 15568 17332
rect 15519 17292 15568 17320
rect 15519 17289 15531 17292
rect 15473 17283 15531 17289
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 16577 17323 16635 17329
rect 16577 17289 16589 17323
rect 16623 17320 16635 17323
rect 16758 17320 16764 17332
rect 16623 17292 16764 17320
rect 16623 17289 16635 17292
rect 16577 17283 16635 17289
rect 16758 17280 16764 17292
rect 16816 17280 16822 17332
rect 16853 17323 16911 17329
rect 16853 17289 16865 17323
rect 16899 17320 16911 17323
rect 18690 17320 18696 17332
rect 16899 17292 18696 17320
rect 16899 17289 16911 17292
rect 16853 17283 16911 17289
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 18782 17280 18788 17332
rect 18840 17280 18846 17332
rect 17405 17255 17463 17261
rect 17405 17221 17417 17255
rect 17451 17252 17463 17255
rect 18800 17252 18828 17280
rect 17451 17224 18828 17252
rect 17451 17221 17463 17224
rect 17405 17215 17463 17221
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 16960 17156 17693 17184
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17085 15347 17119
rect 15289 17079 15347 17085
rect 15378 17076 15384 17128
rect 15436 17076 15442 17128
rect 16669 17119 16727 17125
rect 16669 17085 16681 17119
rect 16715 17085 16727 17119
rect 16669 17079 16727 17085
rect 16684 17048 16712 17079
rect 16758 17076 16764 17128
rect 16816 17076 16822 17128
rect 16960 17048 16988 17156
rect 17681 17153 17693 17156
rect 17727 17184 17739 17187
rect 17727 17156 18184 17184
rect 17727 17153 17739 17156
rect 17681 17147 17739 17153
rect 17037 17119 17095 17125
rect 17037 17085 17049 17119
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 17497 17119 17555 17125
rect 17497 17085 17509 17119
rect 17543 17116 17555 17119
rect 17543 17088 17724 17116
rect 17543 17085 17555 17088
rect 17497 17079 17555 17085
rect 14200 17020 14688 17048
rect 11112 17008 11118 17020
rect 11900 16992 11928 17020
rect 9306 16980 9312 16992
rect 8220 16952 9312 16980
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 11882 16940 11888 16992
rect 11940 16940 11946 16992
rect 14090 16940 14096 16992
rect 14148 16980 14154 16992
rect 14660 16989 14688 17020
rect 16684 17020 16988 17048
rect 16684 16992 16712 17020
rect 14369 16983 14427 16989
rect 14369 16980 14381 16983
rect 14148 16952 14381 16980
rect 14148 16940 14154 16952
rect 14369 16949 14381 16952
rect 14415 16949 14427 16983
rect 14369 16943 14427 16949
rect 14645 16983 14703 16989
rect 14645 16949 14657 16983
rect 14691 16980 14703 16983
rect 14921 16983 14979 16989
rect 14921 16980 14933 16983
rect 14691 16952 14933 16980
rect 14691 16949 14703 16952
rect 14645 16943 14703 16949
rect 14921 16949 14933 16952
rect 14967 16980 14979 16983
rect 15194 16980 15200 16992
rect 14967 16952 15200 16980
rect 14967 16949 14979 16952
rect 14921 16943 14979 16949
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 16666 16940 16672 16992
rect 16724 16940 16730 16992
rect 16942 16940 16948 16992
rect 17000 16980 17006 16992
rect 17052 16980 17080 17079
rect 17129 17051 17187 17057
rect 17129 17017 17141 17051
rect 17175 17048 17187 17051
rect 17310 17048 17316 17060
rect 17175 17020 17316 17048
rect 17175 17017 17187 17020
rect 17129 17011 17187 17017
rect 17310 17008 17316 17020
rect 17368 17008 17374 17060
rect 17696 17048 17724 17088
rect 17770 17076 17776 17128
rect 17828 17076 17834 17128
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18156 17125 18184 17156
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 18012 17088 18061 17116
rect 18012 17076 18018 17088
rect 18049 17085 18061 17088
rect 18095 17085 18107 17119
rect 18049 17079 18107 17085
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 18690 17076 18696 17128
rect 18748 17118 18754 17128
rect 18748 17090 18791 17118
rect 18748 17076 18754 17090
rect 17696 17020 17908 17048
rect 17880 16992 17908 17020
rect 17000 16952 17080 16980
rect 17000 16940 17006 16952
rect 17862 16940 17868 16992
rect 17920 16980 17926 16992
rect 17957 16983 18015 16989
rect 17957 16980 17969 16983
rect 17920 16952 17969 16980
rect 17920 16940 17926 16952
rect 17957 16949 17969 16952
rect 18003 16949 18015 16983
rect 17957 16943 18015 16949
rect 18230 16940 18236 16992
rect 18288 16940 18294 16992
rect 552 16890 19571 16912
rect 552 16838 5112 16890
rect 5164 16838 5176 16890
rect 5228 16838 5240 16890
rect 5292 16838 5304 16890
rect 5356 16838 5368 16890
rect 5420 16838 9827 16890
rect 9879 16838 9891 16890
rect 9943 16838 9955 16890
rect 10007 16838 10019 16890
rect 10071 16838 10083 16890
rect 10135 16838 14542 16890
rect 14594 16838 14606 16890
rect 14658 16838 14670 16890
rect 14722 16838 14734 16890
rect 14786 16838 14798 16890
rect 14850 16838 19257 16890
rect 19309 16838 19321 16890
rect 19373 16838 19385 16890
rect 19437 16838 19449 16890
rect 19501 16838 19513 16890
rect 19565 16838 19571 16890
rect 552 16816 19571 16838
rect 1305 16779 1363 16785
rect 1305 16745 1317 16779
rect 1351 16776 1363 16779
rect 1394 16776 1400 16788
rect 1351 16748 1400 16776
rect 1351 16745 1363 16748
rect 1305 16739 1363 16745
rect 1394 16736 1400 16748
rect 1452 16776 1458 16788
rect 1854 16776 1860 16788
rect 1452 16748 1860 16776
rect 1452 16736 1458 16748
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2222 16736 2228 16788
rect 2280 16736 2286 16788
rect 2314 16736 2320 16788
rect 2372 16776 2378 16788
rect 2409 16779 2467 16785
rect 2409 16776 2421 16779
rect 2372 16748 2421 16776
rect 2372 16736 2378 16748
rect 2409 16745 2421 16748
rect 2455 16745 2467 16779
rect 2409 16739 2467 16745
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 2961 16779 3019 16785
rect 2961 16776 2973 16779
rect 2832 16748 2973 16776
rect 2832 16736 2838 16748
rect 2961 16745 2973 16748
rect 3007 16745 3019 16779
rect 2961 16739 3019 16745
rect 3142 16736 3148 16788
rect 3200 16736 3206 16788
rect 3237 16779 3295 16785
rect 3237 16745 3249 16779
rect 3283 16776 3295 16779
rect 3694 16776 3700 16788
rect 3283 16748 3700 16776
rect 3283 16745 3295 16748
rect 3237 16739 3295 16745
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 1578 16640 1584 16652
rect 1443 16612 1584 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 1673 16643 1731 16649
rect 1673 16609 1685 16643
rect 1719 16640 1731 16643
rect 1949 16643 2007 16649
rect 1719 16612 1900 16640
rect 1719 16609 1731 16612
rect 1673 16603 1731 16609
rect 1872 16572 1900 16612
rect 1949 16609 1961 16643
rect 1995 16640 2007 16643
rect 2041 16643 2099 16649
rect 2041 16640 2053 16643
rect 1995 16612 2053 16640
rect 1995 16609 2007 16612
rect 1949 16603 2007 16609
rect 2041 16609 2053 16612
rect 2087 16640 2099 16643
rect 2240 16640 2268 16736
rect 2590 16708 2596 16720
rect 2087 16612 2268 16640
rect 2332 16680 2596 16708
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 2332 16572 2360 16680
rect 2590 16668 2596 16680
rect 2648 16668 2654 16720
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16609 2559 16643
rect 2608 16640 2636 16668
rect 3160 16649 3188 16736
rect 2685 16643 2743 16649
rect 2685 16640 2697 16643
rect 2608 16612 2697 16640
rect 2501 16603 2559 16609
rect 2685 16609 2697 16612
rect 2731 16609 2743 16643
rect 2685 16603 2743 16609
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 3053 16643 3111 16649
rect 2823 16612 3004 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 1872 16544 2360 16572
rect 1854 16396 1860 16448
rect 1912 16396 1918 16448
rect 2133 16439 2191 16445
rect 2133 16405 2145 16439
rect 2179 16436 2191 16439
rect 2406 16436 2412 16448
rect 2179 16408 2412 16436
rect 2179 16405 2191 16408
rect 2133 16399 2191 16405
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 2516 16436 2544 16603
rect 2976 16504 3004 16612
rect 3053 16609 3065 16643
rect 3099 16609 3111 16643
rect 3053 16603 3111 16609
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16609 3203 16643
rect 3145 16603 3203 16609
rect 3068 16572 3096 16603
rect 3252 16584 3280 16739
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 3878 16736 3884 16788
rect 3936 16776 3942 16788
rect 4065 16779 4123 16785
rect 4065 16776 4077 16779
rect 3936 16748 4077 16776
rect 3936 16736 3942 16748
rect 4065 16745 4077 16748
rect 4111 16776 4123 16779
rect 4617 16779 4675 16785
rect 4617 16776 4629 16779
rect 4111 16748 4629 16776
rect 4111 16745 4123 16748
rect 4065 16739 4123 16745
rect 4617 16745 4629 16748
rect 4663 16776 4675 16779
rect 4798 16776 4804 16788
rect 4663 16748 4804 16776
rect 4663 16745 4675 16748
rect 4617 16739 4675 16745
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 4982 16736 4988 16788
rect 5040 16776 5046 16788
rect 5537 16779 5595 16785
rect 5537 16776 5549 16779
rect 5040 16748 5549 16776
rect 5040 16736 5046 16748
rect 5537 16745 5549 16748
rect 5583 16745 5595 16779
rect 5537 16739 5595 16745
rect 6086 16736 6092 16788
rect 6144 16776 6150 16788
rect 6546 16776 6552 16788
rect 6144 16748 6408 16776
rect 6144 16736 6150 16748
rect 4338 16668 4344 16720
rect 4396 16708 4402 16720
rect 6380 16717 6408 16748
rect 6472 16748 6552 16776
rect 4893 16711 4951 16717
rect 4893 16708 4905 16711
rect 4396 16680 4905 16708
rect 4396 16668 4402 16680
rect 4893 16677 4905 16680
rect 4939 16708 4951 16711
rect 5261 16711 5319 16717
rect 5261 16708 5273 16711
rect 4939 16680 5273 16708
rect 4939 16677 4951 16680
rect 4893 16671 4951 16677
rect 5261 16677 5273 16680
rect 5307 16677 5319 16711
rect 6365 16711 6423 16717
rect 5261 16671 5319 16677
rect 5736 16680 6132 16708
rect 3697 16643 3755 16649
rect 3697 16640 3709 16643
rect 3344 16612 3709 16640
rect 3234 16572 3240 16584
rect 3068 16544 3240 16572
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 3344 16504 3372 16612
rect 3697 16609 3709 16612
rect 3743 16640 3755 16643
rect 4062 16640 4068 16652
rect 3743 16612 4068 16640
rect 3743 16609 3755 16612
rect 3697 16603 3755 16609
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16609 4215 16643
rect 4157 16603 4215 16609
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16640 4307 16643
rect 4356 16640 4384 16668
rect 5736 16652 5764 16680
rect 4295 16612 4384 16640
rect 4709 16643 4767 16649
rect 4295 16609 4307 16612
rect 4249 16603 4307 16609
rect 4709 16609 4721 16643
rect 4755 16640 4767 16643
rect 4755 16612 4936 16640
rect 4755 16609 4767 16612
rect 4709 16603 4767 16609
rect 4172 16572 4200 16603
rect 4908 16572 4936 16612
rect 4982 16600 4988 16652
rect 5040 16600 5046 16652
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16640 5411 16643
rect 5534 16640 5540 16652
rect 5399 16612 5540 16640
rect 5399 16609 5411 16612
rect 5353 16603 5411 16609
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16609 5687 16643
rect 5629 16603 5687 16609
rect 5644 16572 5672 16603
rect 5718 16600 5724 16652
rect 5776 16600 5782 16652
rect 5994 16640 6000 16652
rect 6052 16649 6058 16652
rect 6104 16649 6132 16680
rect 6365 16677 6377 16711
rect 6411 16677 6423 16711
rect 6365 16671 6423 16677
rect 5963 16612 6000 16640
rect 5994 16600 6000 16612
rect 6052 16603 6063 16649
rect 6104 16643 6167 16649
rect 6104 16612 6121 16643
rect 6109 16609 6121 16612
rect 6155 16609 6167 16643
rect 6109 16603 6167 16609
rect 6052 16600 6058 16603
rect 6270 16600 6276 16652
rect 6328 16600 6334 16652
rect 6472 16649 6500 16748
rect 6546 16736 6552 16748
rect 6604 16776 6610 16788
rect 7926 16776 7932 16788
rect 6604 16748 7932 16776
rect 6604 16736 6610 16748
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 9493 16779 9551 16785
rect 9493 16745 9505 16779
rect 9539 16776 9551 16779
rect 10778 16776 10784 16788
rect 9539 16748 10784 16776
rect 9539 16745 9551 16748
rect 9493 16739 9551 16745
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 10870 16736 10876 16788
rect 10928 16736 10934 16788
rect 11054 16736 11060 16788
rect 11112 16736 11118 16788
rect 11606 16736 11612 16788
rect 11664 16776 11670 16788
rect 11885 16779 11943 16785
rect 11885 16776 11897 16779
rect 11664 16748 11897 16776
rect 11664 16736 11670 16748
rect 11885 16745 11897 16748
rect 11931 16745 11943 16779
rect 14918 16776 14924 16788
rect 11885 16739 11943 16745
rect 14752 16748 14924 16776
rect 6932 16680 8248 16708
rect 6932 16649 6960 16680
rect 8220 16652 8248 16680
rect 6457 16643 6515 16649
rect 6457 16609 6469 16643
rect 6503 16609 6515 16643
rect 6457 16603 6515 16609
rect 6917 16643 6975 16649
rect 6917 16609 6929 16643
rect 6963 16609 6975 16643
rect 6917 16603 6975 16609
rect 7742 16600 7748 16652
rect 7800 16600 7806 16652
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16609 8171 16643
rect 8113 16603 8171 16609
rect 5902 16572 5908 16584
rect 4172 16544 4384 16572
rect 4908 16544 5908 16572
rect 2976 16476 3372 16504
rect 4246 16464 4252 16516
rect 4304 16504 4310 16516
rect 4356 16513 4384 16544
rect 5902 16532 5908 16544
rect 5960 16532 5966 16584
rect 6288 16572 6316 16600
rect 7760 16572 7788 16600
rect 6288 16544 7788 16572
rect 4341 16507 4399 16513
rect 4341 16504 4353 16507
rect 4304 16476 4353 16504
rect 4304 16464 4310 16476
rect 4341 16473 4353 16476
rect 4387 16504 4399 16507
rect 4387 16476 6868 16504
rect 4387 16473 4399 16476
rect 4341 16467 4399 16473
rect 6840 16448 6868 16476
rect 3605 16439 3663 16445
rect 3605 16436 3617 16439
rect 2516 16408 3617 16436
rect 3605 16405 3617 16408
rect 3651 16436 3663 16439
rect 3786 16436 3792 16448
rect 3651 16408 3792 16436
rect 3651 16405 3663 16408
rect 3605 16399 3663 16405
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 6638 16396 6644 16448
rect 6696 16396 6702 16448
rect 6822 16396 6828 16448
rect 6880 16396 6886 16448
rect 8128 16436 8156 16603
rect 8202 16600 8208 16652
rect 8260 16640 8266 16652
rect 8369 16643 8427 16649
rect 8369 16640 8381 16643
rect 8260 16612 8381 16640
rect 8260 16600 8266 16612
rect 8369 16609 8381 16612
rect 8415 16609 8427 16643
rect 10888 16640 10916 16736
rect 13906 16668 13912 16720
rect 13964 16708 13970 16720
rect 14642 16708 14648 16720
rect 13964 16680 14648 16708
rect 13964 16668 13970 16680
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 11149 16643 11207 16649
rect 10888 16612 11100 16640
rect 8369 16603 8427 16609
rect 11072 16516 11100 16612
rect 11149 16609 11161 16643
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 11164 16572 11192 16603
rect 11422 16600 11428 16652
rect 11480 16600 11486 16652
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16640 11575 16643
rect 11563 16612 11744 16640
rect 11563 16609 11575 16612
rect 11517 16603 11575 16609
rect 11606 16572 11612 16584
rect 11164 16544 11612 16572
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 11054 16464 11060 16516
rect 11112 16504 11118 16516
rect 11333 16507 11391 16513
rect 11333 16504 11345 16507
rect 11112 16476 11345 16504
rect 11112 16464 11118 16476
rect 11333 16473 11345 16476
rect 11379 16504 11391 16507
rect 11716 16504 11744 16612
rect 11974 16600 11980 16652
rect 12032 16600 12038 16652
rect 14090 16600 14096 16652
rect 14148 16640 14154 16652
rect 14752 16649 14780 16748
rect 14918 16736 14924 16748
rect 14976 16776 14982 16788
rect 15473 16779 15531 16785
rect 15473 16776 15485 16779
rect 14976 16748 15485 16776
rect 14976 16736 14982 16748
rect 15473 16745 15485 16748
rect 15519 16776 15531 16779
rect 15749 16779 15807 16785
rect 15749 16776 15761 16779
rect 15519 16748 15761 16776
rect 15519 16745 15531 16748
rect 15473 16739 15531 16745
rect 15749 16745 15761 16748
rect 15795 16745 15807 16779
rect 15749 16739 15807 16745
rect 16666 16736 16672 16788
rect 16724 16736 16730 16788
rect 16942 16736 16948 16788
rect 17000 16776 17006 16788
rect 18230 16776 18236 16788
rect 17000 16748 18236 16776
rect 17000 16736 17006 16748
rect 18230 16736 18236 16748
rect 18288 16736 18294 16788
rect 14826 16668 14832 16720
rect 14884 16708 14890 16720
rect 15197 16711 15255 16717
rect 15197 16708 15209 16711
rect 14884 16680 15209 16708
rect 14884 16668 14890 16680
rect 15197 16677 15209 16680
rect 15243 16677 15255 16711
rect 15197 16671 15255 16677
rect 15562 16668 15568 16720
rect 15620 16668 15626 16720
rect 16776 16680 17908 16708
rect 14461 16643 14519 16649
rect 14148 16612 14412 16640
rect 14148 16600 14154 16612
rect 14384 16572 14412 16612
rect 14461 16609 14473 16643
rect 14507 16640 14519 16643
rect 14737 16643 14795 16649
rect 14737 16640 14749 16643
rect 14507 16612 14749 16640
rect 14507 16609 14519 16612
rect 14461 16603 14519 16609
rect 14737 16609 14749 16612
rect 14783 16609 14795 16643
rect 14737 16603 14795 16609
rect 15010 16600 15016 16652
rect 15068 16600 15074 16652
rect 15102 16600 15108 16652
rect 15160 16600 15166 16652
rect 15381 16643 15439 16649
rect 15381 16609 15393 16643
rect 15427 16609 15439 16643
rect 15580 16640 15608 16668
rect 16776 16649 16804 16680
rect 17880 16652 17908 16680
rect 18046 16668 18052 16720
rect 18104 16708 18110 16720
rect 18104 16680 18552 16708
rect 18104 16668 18110 16680
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 15580 16612 15669 16640
rect 15381 16603 15439 16609
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 16761 16643 16819 16649
rect 16761 16609 16773 16643
rect 16807 16609 16819 16643
rect 16761 16603 16819 16609
rect 17037 16643 17095 16649
rect 17037 16609 17049 16643
rect 17083 16640 17095 16643
rect 17494 16640 17500 16652
rect 17083 16612 17500 16640
rect 17083 16609 17095 16612
rect 17037 16603 17095 16609
rect 15396 16572 15424 16603
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 17862 16600 17868 16652
rect 17920 16640 17926 16652
rect 18524 16649 18552 16680
rect 18242 16643 18300 16649
rect 18242 16640 18254 16643
rect 17920 16612 18254 16640
rect 17920 16600 17926 16612
rect 18242 16609 18254 16612
rect 18288 16609 18300 16643
rect 18242 16603 18300 16609
rect 18509 16643 18567 16649
rect 18509 16609 18521 16643
rect 18555 16609 18567 16643
rect 18509 16603 18567 16609
rect 18598 16600 18604 16652
rect 18656 16600 18662 16652
rect 19058 16600 19064 16652
rect 19116 16600 19122 16652
rect 14384 16544 15424 16572
rect 17218 16532 17224 16584
rect 17276 16532 17282 16584
rect 11379 16476 11744 16504
rect 11379 16473 11391 16476
rect 11333 16467 11391 16473
rect 13170 16464 13176 16516
rect 13228 16504 13234 16516
rect 17236 16504 17264 16532
rect 13228 16476 17264 16504
rect 13228 16464 13234 16476
rect 17310 16464 17316 16516
rect 17368 16464 17374 16516
rect 8386 16436 8392 16448
rect 8128 16408 8392 16436
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 11882 16436 11888 16448
rect 11204 16408 11888 16436
rect 11204 16396 11210 16408
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 13998 16396 14004 16448
rect 14056 16396 14062 16448
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 14369 16439 14427 16445
rect 14369 16436 14381 16439
rect 14332 16408 14381 16436
rect 14332 16396 14338 16408
rect 14369 16405 14381 16408
rect 14415 16405 14427 16439
rect 14369 16399 14427 16405
rect 14645 16439 14703 16445
rect 14645 16405 14657 16439
rect 14691 16436 14703 16439
rect 14826 16436 14832 16448
rect 14691 16408 14832 16436
rect 14691 16405 14703 16408
rect 14645 16399 14703 16405
rect 14826 16396 14832 16408
rect 14884 16396 14890 16448
rect 14921 16439 14979 16445
rect 14921 16405 14933 16439
rect 14967 16436 14979 16439
rect 15102 16436 15108 16448
rect 14967 16408 15108 16436
rect 14967 16405 14979 16408
rect 14921 16399 14979 16405
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 17129 16439 17187 16445
rect 17129 16405 17141 16439
rect 17175 16436 17187 16439
rect 17218 16436 17224 16448
rect 17175 16408 17224 16436
rect 17175 16405 17187 16408
rect 17129 16399 17187 16405
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 17328 16436 17356 16464
rect 18690 16436 18696 16448
rect 17328 16408 18696 16436
rect 18690 16396 18696 16408
rect 18748 16396 18754 16448
rect 552 16346 19412 16368
rect 552 16294 2755 16346
rect 2807 16294 2819 16346
rect 2871 16294 2883 16346
rect 2935 16294 2947 16346
rect 2999 16294 3011 16346
rect 3063 16294 7470 16346
rect 7522 16294 7534 16346
rect 7586 16294 7598 16346
rect 7650 16294 7662 16346
rect 7714 16294 7726 16346
rect 7778 16294 12185 16346
rect 12237 16294 12249 16346
rect 12301 16294 12313 16346
rect 12365 16294 12377 16346
rect 12429 16294 12441 16346
rect 12493 16294 16900 16346
rect 16952 16294 16964 16346
rect 17016 16294 17028 16346
rect 17080 16294 17092 16346
rect 17144 16294 17156 16346
rect 17208 16294 19412 16346
rect 552 16272 19412 16294
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5353 16235 5411 16241
rect 5353 16232 5365 16235
rect 5040 16204 5365 16232
rect 5040 16192 5046 16204
rect 5353 16201 5365 16204
rect 5399 16201 5411 16235
rect 5353 16195 5411 16201
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 5629 16235 5687 16241
rect 5629 16232 5641 16235
rect 5592 16204 5641 16232
rect 5592 16192 5598 16204
rect 5629 16201 5641 16204
rect 5675 16201 5687 16235
rect 5629 16195 5687 16201
rect 1578 16124 1584 16176
rect 1636 16164 1642 16176
rect 2593 16167 2651 16173
rect 2593 16164 2605 16167
rect 1636 16136 2605 16164
rect 1636 16124 1642 16136
rect 1412 16068 1992 16096
rect 1412 16040 1440 16068
rect 1394 15988 1400 16040
rect 1452 15988 1458 16040
rect 1854 15988 1860 16040
rect 1912 15988 1918 16040
rect 1964 16037 1992 16068
rect 2424 16037 2452 16136
rect 2593 16133 2605 16136
rect 2639 16133 2651 16167
rect 2593 16127 2651 16133
rect 2498 16056 2504 16108
rect 2556 16056 2562 16108
rect 5644 16096 5672 16195
rect 5902 16192 5908 16244
rect 5960 16232 5966 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5960 16204 6193 16232
rect 5960 16192 5966 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 6181 16195 6239 16201
rect 6288 16204 8033 16232
rect 5905 16099 5963 16105
rect 5644 16068 5856 16096
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 15997 2007 16031
rect 1949 15991 2007 15997
rect 2409 16031 2467 16037
rect 2409 15997 2421 16031
rect 2455 15997 2467 16031
rect 2516 16028 2544 16056
rect 2685 16031 2743 16037
rect 2685 16028 2697 16031
rect 2516 16000 2697 16028
rect 2409 15991 2467 15997
rect 2685 15997 2697 16000
rect 2731 15997 2743 16031
rect 2685 15991 2743 15997
rect 1489 15963 1547 15969
rect 1489 15929 1501 15963
rect 1535 15960 1547 15963
rect 1872 15960 1900 15988
rect 2700 15960 2728 15991
rect 3234 15988 3240 16040
rect 3292 16028 3298 16040
rect 3602 16028 3608 16040
rect 3292 16000 3608 16028
rect 3292 15988 3298 16000
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 5828 16037 5856 16068
rect 5905 16065 5917 16099
rect 5951 16096 5963 16099
rect 5994 16096 6000 16108
rect 5951 16068 6000 16096
rect 5951 16065 5963 16068
rect 5905 16059 5963 16065
rect 5994 16056 6000 16068
rect 6052 16096 6058 16108
rect 6288 16096 6316 16204
rect 8021 16201 8033 16204
rect 8067 16232 8079 16235
rect 8202 16232 8208 16244
rect 8067 16204 8208 16232
rect 8067 16201 8079 16204
rect 8021 16195 8079 16201
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 9306 16192 9312 16244
rect 9364 16232 9370 16244
rect 11146 16232 11152 16244
rect 9364 16204 11152 16232
rect 9364 16192 9370 16204
rect 9769 16167 9827 16173
rect 9769 16133 9781 16167
rect 9815 16133 9827 16167
rect 9769 16127 9827 16133
rect 6052 16068 6316 16096
rect 8036 16068 8432 16096
rect 6052 16056 6058 16068
rect 5445 16031 5503 16037
rect 5445 15997 5457 16031
rect 5491 16028 5503 16031
rect 5721 16031 5779 16037
rect 5721 16028 5733 16031
rect 5491 16000 5733 16028
rect 5491 15997 5503 16000
rect 5445 15991 5503 15997
rect 5721 15997 5733 16000
rect 5767 15997 5779 16031
rect 5721 15991 5779 15997
rect 5813 16031 5871 16037
rect 5813 15997 5825 16031
rect 5859 15997 5871 16031
rect 5813 15991 5871 15997
rect 6273 16031 6331 16037
rect 6273 15997 6285 16031
rect 6319 15997 6331 16031
rect 6273 15991 6331 15997
rect 6457 16031 6515 16037
rect 6457 15997 6469 16031
rect 6503 16028 6515 16031
rect 8036 16028 8064 16068
rect 8404 16040 8432 16068
rect 6503 16000 8064 16028
rect 8113 16031 8171 16037
rect 6503 15997 6515 16000
rect 6457 15991 6515 15997
rect 8113 15997 8125 16031
rect 8159 15997 8171 16031
rect 8113 15991 8171 15997
rect 3329 15963 3387 15969
rect 3329 15960 3341 15963
rect 1535 15932 2452 15960
rect 2700 15932 3341 15960
rect 1535 15929 1547 15932
rect 1489 15923 1547 15929
rect 2424 15904 2452 15932
rect 3329 15929 3341 15932
rect 3375 15960 3387 15963
rect 3510 15960 3516 15972
rect 3375 15932 3516 15960
rect 3375 15929 3387 15932
rect 3329 15923 3387 15929
rect 3510 15920 3516 15932
rect 3568 15920 3574 15972
rect 5460 15904 5488 15991
rect 6288 15904 6316 15991
rect 6724 15963 6782 15969
rect 6724 15929 6736 15963
rect 6770 15960 6782 15963
rect 6822 15960 6828 15972
rect 6770 15932 6828 15960
rect 6770 15929 6782 15932
rect 6724 15923 6782 15929
rect 6822 15920 6828 15932
rect 6880 15920 6886 15972
rect 7558 15920 7564 15972
rect 7616 15960 7622 15972
rect 8128 15960 8156 15991
rect 8386 15988 8392 16040
rect 8444 15988 8450 16040
rect 9784 16028 9812 16127
rect 10520 16037 10548 16204
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 13998 16192 14004 16244
rect 14056 16232 14062 16244
rect 14093 16235 14151 16241
rect 14093 16232 14105 16235
rect 14056 16204 14105 16232
rect 14056 16192 14062 16204
rect 14093 16201 14105 16204
rect 14139 16201 14151 16235
rect 14093 16195 14151 16201
rect 15286 16192 15292 16244
rect 15344 16232 15350 16244
rect 15344 16204 15700 16232
rect 15344 16192 15350 16204
rect 10689 16167 10747 16173
rect 10689 16133 10701 16167
rect 10735 16164 10747 16167
rect 11330 16164 11336 16176
rect 10735 16136 11336 16164
rect 10735 16133 10747 16136
rect 10689 16127 10747 16133
rect 11330 16124 11336 16136
rect 11388 16124 11394 16176
rect 11514 16124 11520 16176
rect 11572 16164 11578 16176
rect 14277 16167 14335 16173
rect 14277 16164 14289 16167
rect 11572 16136 14289 16164
rect 11572 16124 11578 16136
rect 14277 16133 14289 16136
rect 14323 16133 14335 16167
rect 14277 16127 14335 16133
rect 15672 16105 15700 16204
rect 17494 16192 17500 16244
rect 17552 16232 17558 16244
rect 17589 16235 17647 16241
rect 17589 16232 17601 16235
rect 17552 16204 17601 16232
rect 17552 16192 17558 16204
rect 17589 16201 17601 16204
rect 17635 16201 17647 16235
rect 17589 16195 17647 16201
rect 15657 16099 15715 16105
rect 10704 16068 14228 16096
rect 10137 16031 10195 16037
rect 10137 16028 10149 16031
rect 9784 16000 10149 16028
rect 10137 15997 10149 16000
rect 10183 15997 10195 16031
rect 10520 16031 10587 16037
rect 10520 16000 10541 16031
rect 10137 15991 10195 15997
rect 10529 15997 10541 16000
rect 10575 15997 10587 16031
rect 10529 15991 10587 15997
rect 8634 15963 8692 15969
rect 8634 15960 8646 15963
rect 7616 15932 8646 15960
rect 7616 15920 7622 15932
rect 8634 15929 8646 15932
rect 8680 15929 8692 15963
rect 8634 15923 8692 15929
rect 9122 15920 9128 15972
rect 9180 15960 9186 15972
rect 10321 15963 10379 15969
rect 10321 15960 10333 15963
rect 9180 15932 10333 15960
rect 9180 15920 9186 15932
rect 10321 15929 10333 15932
rect 10367 15929 10379 15963
rect 10321 15923 10379 15929
rect 10413 15963 10471 15969
rect 10413 15929 10425 15963
rect 10459 15960 10471 15963
rect 10704 15960 10732 16068
rect 10778 15988 10784 16040
rect 10836 15988 10842 16040
rect 11146 15988 11152 16040
rect 11204 15988 11210 16040
rect 11517 16031 11575 16037
rect 11517 15997 11529 16031
rect 11563 16028 11575 16031
rect 11606 16028 11612 16040
rect 11563 16000 11612 16028
rect 11563 15997 11575 16000
rect 11517 15991 11575 15997
rect 11606 15988 11612 16000
rect 11664 16028 11670 16040
rect 12342 16028 12348 16040
rect 11664 16000 12348 16028
rect 11664 15988 11670 16000
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 13170 15988 13176 16040
rect 13228 15988 13234 16040
rect 13357 16031 13415 16037
rect 13357 15997 13369 16031
rect 13403 16028 13415 16031
rect 13906 16028 13912 16040
rect 13403 16000 13912 16028
rect 13403 15997 13415 16000
rect 13357 15991 13415 15997
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 16028 14059 16031
rect 14200 16028 14228 16068
rect 15657 16065 15669 16099
rect 15703 16065 15715 16099
rect 17604 16096 17632 16195
rect 17862 16192 17868 16244
rect 17920 16192 17926 16244
rect 17770 16124 17776 16176
rect 17828 16164 17834 16176
rect 18414 16164 18420 16176
rect 17828 16136 18420 16164
rect 17828 16124 17834 16136
rect 18414 16124 18420 16136
rect 18472 16124 18478 16176
rect 17604 16068 18092 16096
rect 15657 16059 15715 16065
rect 17218 16028 17224 16040
rect 14047 16000 14136 16028
rect 14200 16000 17224 16028
rect 14047 15997 14059 16000
rect 14001 15991 14059 15997
rect 10459 15932 10732 15960
rect 10965 15963 11023 15969
rect 10459 15929 10471 15932
rect 10413 15923 10471 15929
rect 10965 15929 10977 15963
rect 11011 15929 11023 15963
rect 10965 15923 11023 15929
rect 11057 15963 11115 15969
rect 11057 15929 11069 15963
rect 11103 15960 11115 15963
rect 13188 15960 13216 15988
rect 11103 15932 13216 15960
rect 13265 15963 13323 15969
rect 11103 15929 11115 15932
rect 11057 15923 11115 15929
rect 13265 15929 13277 15963
rect 13311 15960 13323 15963
rect 14108 15960 14136 16000
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 17681 16031 17739 16037
rect 17681 15997 17693 16031
rect 17727 16028 17739 16031
rect 17770 16028 17776 16040
rect 17727 16000 17776 16028
rect 17727 15997 17739 16000
rect 17681 15991 17739 15997
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 18064 16037 18092 16068
rect 17957 16031 18015 16037
rect 17957 16028 17969 16031
rect 17920 16000 17969 16028
rect 17920 15988 17926 16000
rect 17957 15997 17969 16000
rect 18003 15997 18015 16031
rect 17957 15991 18015 15997
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 18325 16031 18383 16037
rect 18325 15997 18337 16031
rect 18371 15997 18383 16031
rect 18325 15991 18383 15997
rect 13311 15932 14136 15960
rect 13311 15929 13323 15932
rect 13265 15923 13323 15929
rect 1762 15852 1768 15904
rect 1820 15852 1826 15904
rect 2041 15895 2099 15901
rect 2041 15861 2053 15895
rect 2087 15892 2099 15895
rect 2222 15892 2228 15904
rect 2087 15864 2228 15892
rect 2087 15861 2099 15864
rect 2041 15855 2099 15861
rect 2222 15852 2228 15864
rect 2280 15852 2286 15904
rect 2314 15852 2320 15904
rect 2372 15852 2378 15904
rect 2406 15852 2412 15904
rect 2464 15852 2470 15904
rect 5442 15852 5448 15904
rect 5500 15852 5506 15904
rect 6270 15852 6276 15904
rect 6328 15852 6334 15904
rect 7834 15852 7840 15904
rect 7892 15852 7898 15904
rect 10336 15892 10364 15923
rect 10980 15892 11008 15923
rect 14108 15904 14136 15932
rect 15194 15920 15200 15972
rect 15252 15960 15258 15972
rect 15390 15963 15448 15969
rect 15390 15960 15402 15963
rect 15252 15932 15402 15960
rect 15252 15920 15258 15932
rect 15390 15929 15402 15932
rect 15436 15929 15448 15963
rect 17972 15960 18000 15991
rect 18340 15960 18368 15991
rect 17972 15932 18368 15960
rect 15390 15923 15448 15929
rect 10336 15864 11008 15892
rect 11146 15852 11152 15904
rect 11204 15892 11210 15904
rect 11333 15895 11391 15901
rect 11333 15892 11345 15895
rect 11204 15864 11345 15892
rect 11204 15852 11210 15864
rect 11333 15861 11345 15864
rect 11379 15861 11391 15895
rect 11333 15855 11391 15861
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 11609 15895 11667 15901
rect 11609 15892 11621 15895
rect 11480 15864 11621 15892
rect 11480 15852 11486 15864
rect 11609 15861 11621 15864
rect 11655 15892 11667 15895
rect 12066 15892 12072 15904
rect 11655 15864 12072 15892
rect 11655 15861 11667 15864
rect 11609 15855 11667 15861
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 12158 15852 12164 15904
rect 12216 15892 12222 15904
rect 13170 15892 13176 15904
rect 12216 15864 13176 15892
rect 12216 15852 12222 15864
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 13817 15895 13875 15901
rect 13817 15892 13829 15895
rect 13596 15864 13829 15892
rect 13596 15852 13602 15864
rect 13817 15861 13829 15864
rect 13863 15861 13875 15895
rect 13817 15855 13875 15861
rect 14090 15852 14096 15904
rect 14148 15852 14154 15904
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 17954 15892 17960 15904
rect 17368 15864 17960 15892
rect 17368 15852 17374 15864
rect 17954 15852 17960 15864
rect 18012 15892 18018 15904
rect 18141 15895 18199 15901
rect 18141 15892 18153 15895
rect 18012 15864 18153 15892
rect 18012 15852 18018 15864
rect 18141 15861 18153 15864
rect 18187 15892 18199 15895
rect 18598 15892 18604 15904
rect 18187 15864 18604 15892
rect 18187 15861 18199 15864
rect 18141 15855 18199 15861
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 552 15802 19571 15824
rect 552 15750 5112 15802
rect 5164 15750 5176 15802
rect 5228 15750 5240 15802
rect 5292 15750 5304 15802
rect 5356 15750 5368 15802
rect 5420 15750 9827 15802
rect 9879 15750 9891 15802
rect 9943 15750 9955 15802
rect 10007 15750 10019 15802
rect 10071 15750 10083 15802
rect 10135 15750 14542 15802
rect 14594 15750 14606 15802
rect 14658 15750 14670 15802
rect 14722 15750 14734 15802
rect 14786 15750 14798 15802
rect 14850 15750 19257 15802
rect 19309 15750 19321 15802
rect 19373 15750 19385 15802
rect 19437 15750 19449 15802
rect 19501 15750 19513 15802
rect 19565 15750 19571 15802
rect 552 15728 19571 15750
rect 1762 15648 1768 15700
rect 1820 15688 1826 15700
rect 2777 15691 2835 15697
rect 2777 15688 2789 15691
rect 1820 15660 2789 15688
rect 1820 15648 1826 15660
rect 2777 15657 2789 15660
rect 2823 15657 2835 15691
rect 2777 15651 2835 15657
rect 5534 15648 5540 15700
rect 5592 15648 5598 15700
rect 7009 15691 7067 15697
rect 7009 15688 7021 15691
rect 6380 15660 7021 15688
rect 1486 15512 1492 15564
rect 1544 15552 1550 15564
rect 1780 15561 1808 15648
rect 2222 15620 2228 15632
rect 2056 15592 2228 15620
rect 2056 15561 2084 15592
rect 2222 15580 2228 15592
rect 2280 15580 2286 15632
rect 2498 15580 2504 15632
rect 2556 15620 2562 15632
rect 2556 15592 2912 15620
rect 2556 15580 2562 15592
rect 1765 15555 1823 15561
rect 1765 15552 1777 15555
rect 1544 15524 1777 15552
rect 1544 15512 1550 15524
rect 1765 15521 1777 15524
rect 1811 15521 1823 15555
rect 1765 15515 1823 15521
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15552 2191 15555
rect 2179 15524 2360 15552
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 2332 15496 2360 15524
rect 2406 15512 2412 15564
rect 2464 15512 2470 15564
rect 2884 15561 2912 15592
rect 3528 15592 4200 15620
rect 2869 15555 2927 15561
rect 2869 15521 2881 15555
rect 2915 15521 2927 15555
rect 2869 15515 2927 15521
rect 3326 15512 3332 15564
rect 3384 15552 3390 15564
rect 3528 15561 3556 15592
rect 4172 15564 4200 15592
rect 3513 15555 3571 15561
rect 3513 15552 3525 15555
rect 3384 15524 3525 15552
rect 3384 15512 3390 15524
rect 3513 15521 3525 15524
rect 3559 15521 3571 15555
rect 3513 15515 3571 15521
rect 3602 15512 3608 15564
rect 3660 15552 3666 15564
rect 3769 15555 3827 15561
rect 3769 15552 3781 15555
rect 3660 15524 3781 15552
rect 3660 15512 3666 15524
rect 3769 15521 3781 15524
rect 3815 15521 3827 15555
rect 3769 15515 3827 15521
rect 4154 15512 4160 15564
rect 4212 15512 4218 15564
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15552 5411 15555
rect 5629 15555 5687 15561
rect 5399 15524 5580 15552
rect 5399 15521 5411 15524
rect 5353 15515 5411 15521
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15484 1455 15487
rect 2314 15484 2320 15496
rect 1443 15456 2320 15484
rect 1443 15453 1455 15456
rect 1397 15447 1455 15453
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 1949 15419 2007 15425
rect 1949 15385 1961 15419
rect 1995 15416 2007 15419
rect 2038 15416 2044 15428
rect 1995 15388 2044 15416
rect 1995 15385 2007 15388
rect 1949 15379 2007 15385
rect 2038 15376 2044 15388
rect 2096 15416 2102 15428
rect 2501 15419 2559 15425
rect 2501 15416 2513 15419
rect 2096 15388 2513 15416
rect 2096 15376 2102 15388
rect 2501 15385 2513 15388
rect 2547 15385 2559 15419
rect 5552 15416 5580 15524
rect 5629 15521 5641 15555
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 6181 15555 6239 15561
rect 6181 15521 6193 15555
rect 6227 15552 6239 15555
rect 6380 15552 6408 15660
rect 7009 15657 7021 15660
rect 7055 15688 7067 15691
rect 7558 15688 7564 15700
rect 7055 15660 7564 15688
rect 7055 15657 7067 15660
rect 7009 15651 7067 15657
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 7834 15648 7840 15700
rect 7892 15648 7898 15700
rect 11054 15648 11060 15700
rect 11112 15648 11118 15700
rect 11440 15660 11928 15688
rect 7852 15620 7880 15648
rect 11440 15629 11468 15660
rect 11425 15623 11483 15629
rect 6748 15592 7420 15620
rect 7852 15592 11284 15620
rect 6227 15524 6408 15552
rect 6227 15521 6239 15524
rect 6181 15515 6239 15521
rect 5644 15484 5672 15515
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 6748 15561 6776 15592
rect 7392 15564 7420 15592
rect 6641 15555 6699 15561
rect 6641 15552 6653 15555
rect 6512 15524 6653 15552
rect 6512 15512 6518 15524
rect 6641 15521 6653 15524
rect 6687 15521 6699 15555
rect 6641 15515 6699 15521
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15521 6791 15555
rect 6733 15515 6791 15521
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15521 6975 15555
rect 6917 15515 6975 15521
rect 6365 15487 6423 15493
rect 6365 15484 6377 15487
rect 5644 15456 6377 15484
rect 6365 15453 6377 15456
rect 6411 15484 6423 15487
rect 6546 15484 6552 15496
rect 6411 15456 6552 15484
rect 6411 15453 6423 15456
rect 6365 15447 6423 15453
rect 6546 15444 6552 15456
rect 6604 15484 6610 15496
rect 6932 15484 6960 15515
rect 7282 15512 7288 15564
rect 7340 15512 7346 15564
rect 7374 15512 7380 15564
rect 7432 15512 7438 15564
rect 11256 15561 11284 15592
rect 11425 15589 11437 15623
rect 11471 15589 11483 15623
rect 11425 15583 11483 15589
rect 11514 15580 11520 15632
rect 11572 15580 11578 15632
rect 11900 15564 11928 15660
rect 11974 15648 11980 15700
rect 12032 15648 12038 15700
rect 12066 15648 12072 15700
rect 12124 15648 12130 15700
rect 12342 15648 12348 15700
rect 12400 15648 12406 15700
rect 13170 15648 13176 15700
rect 13228 15688 13234 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 13228 15660 13461 15688
rect 13228 15648 13234 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 13449 15651 13507 15657
rect 11992 15620 12020 15648
rect 12621 15623 12679 15629
rect 12621 15620 12633 15623
rect 11992 15592 12633 15620
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15521 7711 15555
rect 7653 15515 7711 15521
rect 11149 15555 11207 15561
rect 11149 15521 11161 15555
rect 11195 15521 11207 15555
rect 11149 15515 11207 15521
rect 11241 15555 11299 15561
rect 11241 15521 11253 15555
rect 11287 15521 11299 15555
rect 11241 15515 11299 15521
rect 6604 15456 6960 15484
rect 7300 15484 7328 15512
rect 7668 15484 7696 15515
rect 7300 15456 7696 15484
rect 11164 15484 11192 15515
rect 11606 15512 11612 15564
rect 11664 15512 11670 15564
rect 11882 15512 11888 15564
rect 11940 15512 11946 15564
rect 12066 15512 12072 15564
rect 12124 15552 12130 15564
rect 12268 15561 12296 15592
rect 12621 15589 12633 15592
rect 12667 15620 12679 15623
rect 12897 15623 12955 15629
rect 12897 15620 12909 15623
rect 12667 15592 12909 15620
rect 12667 15589 12679 15592
rect 12621 15583 12679 15589
rect 12897 15589 12909 15592
rect 12943 15589 12955 15623
rect 12897 15583 12955 15589
rect 12161 15555 12219 15561
rect 12161 15552 12173 15555
rect 12124 15524 12173 15552
rect 12124 15512 12130 15524
rect 12161 15521 12173 15524
rect 12207 15521 12219 15555
rect 12161 15515 12219 15521
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15552 12311 15555
rect 12710 15552 12716 15564
rect 12299 15524 12333 15552
rect 12406 15524 12716 15552
rect 12299 15521 12311 15524
rect 12253 15515 12311 15521
rect 12406 15484 12434 15524
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 12986 15512 12992 15564
rect 13044 15512 13050 15564
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15521 13139 15555
rect 13081 15515 13139 15521
rect 11164 15456 12434 15484
rect 6604 15444 6610 15456
rect 12802 15444 12808 15496
rect 12860 15484 12866 15496
rect 13096 15484 13124 15515
rect 12860 15456 13124 15484
rect 13464 15484 13492 15651
rect 13998 15648 14004 15700
rect 14056 15648 14062 15700
rect 17310 15648 17316 15700
rect 17368 15648 17374 15700
rect 17494 15648 17500 15700
rect 17552 15688 17558 15700
rect 17589 15691 17647 15697
rect 17589 15688 17601 15691
rect 17552 15660 17601 15688
rect 17552 15648 17558 15660
rect 17589 15657 17601 15660
rect 17635 15657 17647 15691
rect 17589 15651 17647 15657
rect 18414 15648 18420 15700
rect 18472 15688 18478 15700
rect 18601 15691 18659 15697
rect 18601 15688 18613 15691
rect 18472 15660 18613 15688
rect 18472 15648 18478 15660
rect 18601 15657 18613 15660
rect 18647 15657 18659 15691
rect 18601 15651 18659 15657
rect 14016 15620 14044 15648
rect 14820 15623 14878 15629
rect 14016 15592 14228 15620
rect 13538 15512 13544 15564
rect 13596 15512 13602 15564
rect 13817 15555 13875 15561
rect 13817 15521 13829 15555
rect 13863 15552 13875 15555
rect 14016 15552 14044 15592
rect 13863 15524 14044 15552
rect 13863 15521 13875 15524
rect 13817 15515 13875 15521
rect 14090 15512 14096 15564
rect 14148 15512 14154 15564
rect 14200 15561 14228 15592
rect 14820 15589 14832 15623
rect 14866 15620 14878 15623
rect 14918 15620 14924 15632
rect 14866 15592 14924 15620
rect 14866 15589 14878 15592
rect 14820 15583 14878 15589
rect 14918 15580 14924 15592
rect 14976 15580 14982 15632
rect 18230 15620 18236 15632
rect 17696 15592 18236 15620
rect 14185 15555 14243 15561
rect 14185 15521 14197 15555
rect 14231 15521 14243 15555
rect 14185 15515 14243 15521
rect 14458 15512 14464 15564
rect 14516 15552 14522 15564
rect 14553 15555 14611 15561
rect 14553 15552 14565 15555
rect 14516 15524 14565 15552
rect 14516 15512 14522 15524
rect 14553 15521 14565 15524
rect 14599 15521 14611 15555
rect 15102 15552 15108 15564
rect 14553 15515 14611 15521
rect 14660 15524 15108 15552
rect 14001 15487 14059 15493
rect 14001 15484 14013 15487
rect 13464 15456 14013 15484
rect 12860 15444 12866 15456
rect 14001 15453 14013 15456
rect 14047 15453 14059 15487
rect 14108 15484 14136 15512
rect 14660 15484 14688 15524
rect 15102 15512 15108 15524
rect 15160 15512 15166 15564
rect 17696 15561 17724 15592
rect 18230 15580 18236 15592
rect 18288 15620 18294 15632
rect 18969 15623 19027 15629
rect 18969 15620 18981 15623
rect 18288 15592 18460 15620
rect 18288 15580 18294 15592
rect 18432 15561 18460 15592
rect 18708 15592 18981 15620
rect 18708 15564 18736 15592
rect 18969 15589 18981 15592
rect 19015 15589 19027 15623
rect 18969 15583 19027 15589
rect 17405 15555 17463 15561
rect 17405 15521 17417 15555
rect 17451 15521 17463 15555
rect 17405 15515 17463 15521
rect 17681 15555 17739 15561
rect 17681 15521 17693 15555
rect 17727 15521 17739 15555
rect 17681 15515 17739 15521
rect 17957 15555 18015 15561
rect 17957 15521 17969 15555
rect 18003 15552 18015 15555
rect 18417 15555 18475 15561
rect 18003 15524 18368 15552
rect 18003 15521 18015 15524
rect 17957 15515 18015 15521
rect 14108 15456 14688 15484
rect 17420 15484 17448 15515
rect 17972 15484 18000 15515
rect 17420 15456 18000 15484
rect 14001 15447 14059 15453
rect 6089 15419 6147 15425
rect 6089 15416 6101 15419
rect 2501 15379 2559 15385
rect 4908 15388 5488 15416
rect 5552 15388 6101 15416
rect 1670 15308 1676 15360
rect 1728 15308 1734 15360
rect 2222 15308 2228 15360
rect 2280 15308 2286 15360
rect 4908 15357 4936 15388
rect 4893 15351 4951 15357
rect 4893 15317 4905 15351
rect 4939 15317 4951 15351
rect 4893 15311 4951 15317
rect 5261 15351 5319 15357
rect 5261 15317 5273 15351
rect 5307 15348 5319 15351
rect 5350 15348 5356 15360
rect 5307 15320 5356 15348
rect 5307 15317 5319 15320
rect 5261 15311 5319 15317
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 5460 15348 5488 15388
rect 6089 15385 6101 15388
rect 6135 15416 6147 15419
rect 6270 15416 6276 15428
rect 6135 15388 6276 15416
rect 6135 15385 6147 15388
rect 6089 15379 6147 15385
rect 6270 15376 6276 15388
rect 6328 15416 6334 15428
rect 7285 15419 7343 15425
rect 7285 15416 7297 15419
rect 6328 15388 7297 15416
rect 6328 15376 6334 15388
rect 7285 15385 7297 15388
rect 7331 15385 7343 15419
rect 7285 15379 7343 15385
rect 10686 15376 10692 15428
rect 10744 15416 10750 15428
rect 10744 15388 13768 15416
rect 10744 15376 10750 15388
rect 8294 15348 8300 15360
rect 5460 15320 8300 15348
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 11790 15308 11796 15360
rect 11848 15308 11854 15360
rect 12526 15308 12532 15360
rect 12584 15348 12590 15360
rect 13173 15351 13231 15357
rect 13173 15348 13185 15351
rect 12584 15320 13185 15348
rect 12584 15308 12590 15320
rect 13173 15317 13185 15320
rect 13219 15348 13231 15351
rect 13538 15348 13544 15360
rect 13219 15320 13544 15348
rect 13219 15317 13231 15320
rect 13173 15311 13231 15317
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 13740 15357 13768 15388
rect 18340 15360 18368 15524
rect 18417 15521 18429 15555
rect 18463 15521 18475 15555
rect 18417 15515 18475 15521
rect 18690 15512 18696 15564
rect 18748 15512 18754 15564
rect 18874 15512 18880 15564
rect 18932 15512 18938 15564
rect 13725 15351 13783 15357
rect 13725 15317 13737 15351
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 15933 15351 15991 15357
rect 15933 15317 15945 15351
rect 15979 15348 15991 15351
rect 16574 15348 16580 15360
rect 15979 15320 16580 15348
rect 15979 15317 15991 15320
rect 15933 15311 15991 15317
rect 16574 15308 16580 15320
rect 16632 15308 16638 15360
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 17862 15348 17868 15360
rect 17460 15320 17868 15348
rect 17460 15308 17466 15320
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 18322 15308 18328 15360
rect 18380 15308 18386 15360
rect 552 15258 19412 15280
rect 552 15206 2755 15258
rect 2807 15206 2819 15258
rect 2871 15206 2883 15258
rect 2935 15206 2947 15258
rect 2999 15206 3011 15258
rect 3063 15206 7470 15258
rect 7522 15206 7534 15258
rect 7586 15206 7598 15258
rect 7650 15206 7662 15258
rect 7714 15206 7726 15258
rect 7778 15206 12185 15258
rect 12237 15206 12249 15258
rect 12301 15206 12313 15258
rect 12365 15206 12377 15258
rect 12429 15206 12441 15258
rect 12493 15206 16900 15258
rect 16952 15206 16964 15258
rect 17016 15206 17028 15258
rect 17080 15206 17092 15258
rect 17144 15206 17156 15258
rect 17208 15206 19412 15258
rect 552 15184 19412 15206
rect 6546 15104 6552 15156
rect 6604 15144 6610 15156
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 6604 15116 6653 15144
rect 6604 15104 6610 15116
rect 6641 15113 6653 15116
rect 6687 15113 6699 15147
rect 6641 15107 6699 15113
rect 6917 15147 6975 15153
rect 6917 15113 6929 15147
rect 6963 15144 6975 15147
rect 7374 15144 7380 15156
rect 6963 15116 7380 15144
rect 6963 15113 6975 15116
rect 6917 15107 6975 15113
rect 7374 15104 7380 15116
rect 7432 15144 7438 15156
rect 7745 15147 7803 15153
rect 7745 15144 7757 15147
rect 7432 15116 7757 15144
rect 7432 15104 7438 15116
rect 7745 15113 7757 15116
rect 7791 15113 7803 15147
rect 7745 15107 7803 15113
rect 9398 15104 9404 15156
rect 9456 15144 9462 15156
rect 9456 15116 9812 15144
rect 9456 15104 9462 15116
rect 2406 15036 2412 15088
rect 2464 15076 2470 15088
rect 2593 15079 2651 15085
rect 2593 15076 2605 15079
rect 2464 15048 2605 15076
rect 2464 15036 2470 15048
rect 2593 15045 2605 15048
rect 2639 15045 2651 15079
rect 2593 15039 2651 15045
rect 9125 15079 9183 15085
rect 9125 15045 9137 15079
rect 9171 15045 9183 15079
rect 9582 15076 9588 15088
rect 9125 15039 9183 15045
rect 9232 15048 9588 15076
rect 9140 15008 9168 15039
rect 6748 14980 7144 15008
rect 1486 14949 1492 14952
rect 1213 14943 1271 14949
rect 1213 14909 1225 14943
rect 1259 14909 1271 14943
rect 1480 14940 1492 14949
rect 1447 14912 1492 14940
rect 1213 14903 1271 14909
rect 1480 14903 1492 14912
rect 1228 14872 1256 14903
rect 1486 14900 1492 14903
rect 1544 14900 1550 14952
rect 2314 14900 2320 14952
rect 2372 14940 2378 14952
rect 2685 14943 2743 14949
rect 2685 14940 2697 14943
rect 2372 14912 2697 14940
rect 2372 14900 2378 14912
rect 2685 14909 2697 14912
rect 2731 14909 2743 14943
rect 2685 14903 2743 14909
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14940 3295 14943
rect 3326 14940 3332 14952
rect 3283 14912 3332 14940
rect 3283 14909 3295 14912
rect 3237 14903 3295 14909
rect 2866 14872 2872 14884
rect 1228 14844 2872 14872
rect 2866 14832 2872 14844
rect 2924 14872 2930 14884
rect 3252 14872 3280 14903
rect 3326 14900 3332 14912
rect 3384 14940 3390 14952
rect 6748 14949 6776 14980
rect 7116 14949 7144 14980
rect 8680 14980 9168 15008
rect 5077 14943 5135 14949
rect 5077 14940 5089 14943
rect 3384 14912 5089 14940
rect 3384 14900 3390 14912
rect 5077 14909 5089 14912
rect 5123 14909 5135 14943
rect 6733 14943 6791 14949
rect 6733 14940 6745 14943
rect 5077 14903 5135 14909
rect 6288 14912 6745 14940
rect 3510 14881 3516 14884
rect 3504 14872 3516 14881
rect 2924 14844 3280 14872
rect 3471 14844 3516 14872
rect 2924 14832 2930 14844
rect 3504 14835 3516 14844
rect 3510 14832 3516 14835
rect 3568 14832 3574 14884
rect 5350 14881 5356 14884
rect 5344 14835 5356 14881
rect 5408 14872 5414 14884
rect 5902 14872 5908 14884
rect 5408 14844 5908 14872
rect 5350 14832 5356 14835
rect 5408 14832 5414 14844
rect 5902 14832 5908 14844
rect 5960 14832 5966 14884
rect 6288 14816 6316 14912
rect 6733 14909 6745 14912
rect 6779 14909 6791 14943
rect 6733 14903 6791 14909
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14909 7067 14943
rect 7009 14903 7067 14909
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14940 7159 14943
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 7147 14912 7481 14940
rect 7147 14909 7159 14912
rect 7101 14903 7159 14909
rect 7469 14909 7481 14912
rect 7515 14909 7527 14943
rect 7469 14903 7527 14909
rect 7024 14872 7052 14903
rect 7558 14900 7564 14952
rect 7616 14940 7622 14952
rect 7616 14912 7788 14940
rect 7616 14900 7622 14912
rect 7760 14872 7788 14912
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 8113 14943 8171 14949
rect 8113 14909 8125 14943
rect 8159 14940 8171 14943
rect 8202 14940 8208 14952
rect 8159 14912 8208 14940
rect 8159 14909 8171 14912
rect 8113 14903 8171 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 8680 14949 8708 14980
rect 8665 14943 8723 14949
rect 8665 14940 8677 14943
rect 8628 14912 8677 14940
rect 8628 14900 8634 14912
rect 8665 14909 8677 14912
rect 8711 14909 8723 14943
rect 8665 14903 8723 14909
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14909 8999 14943
rect 8941 14903 8999 14909
rect 8021 14875 8079 14881
rect 8021 14872 8033 14875
rect 7024 14844 7236 14872
rect 7760 14844 8033 14872
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 2777 14807 2835 14813
rect 2777 14804 2789 14807
rect 2648 14776 2789 14804
rect 2648 14764 2654 14776
rect 2777 14773 2789 14776
rect 2823 14773 2835 14807
rect 2777 14767 2835 14773
rect 4614 14764 4620 14816
rect 4672 14764 4678 14816
rect 6270 14764 6276 14816
rect 6328 14764 6334 14816
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 7208 14813 7236 14844
rect 8021 14841 8033 14844
rect 8067 14872 8079 14875
rect 8849 14875 8907 14881
rect 8849 14872 8861 14875
rect 8067 14844 8861 14872
rect 8067 14841 8079 14844
rect 8021 14835 8079 14841
rect 8849 14841 8861 14844
rect 8895 14841 8907 14875
rect 8956 14872 8984 14903
rect 9030 14900 9036 14952
rect 9088 14940 9094 14952
rect 9232 14949 9260 15048
rect 9582 15036 9588 15048
rect 9640 15036 9646 15088
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 9088 14912 9229 14940
rect 9088 14900 9094 14912
rect 9217 14909 9229 14912
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 9398 14900 9404 14952
rect 9456 14942 9462 14952
rect 9493 14945 9551 14951
rect 9493 14942 9505 14945
rect 9456 14914 9505 14942
rect 9456 14900 9462 14914
rect 9493 14911 9505 14914
rect 9539 14911 9551 14945
rect 9493 14905 9551 14911
rect 9582 14900 9588 14952
rect 9640 14940 9646 14952
rect 9784 14949 9812 15116
rect 10410 15104 10416 15156
rect 10468 15144 10474 15156
rect 11606 15144 11612 15156
rect 10468 15116 11612 15144
rect 10468 15104 10474 15116
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 12529 15147 12587 15153
rect 12529 15144 12541 15147
rect 12308 15116 12541 15144
rect 12308 15104 12314 15116
rect 12529 15113 12541 15116
rect 12575 15144 12587 15147
rect 12618 15144 12624 15156
rect 12575 15116 12624 15144
rect 12575 15113 12587 15116
rect 12529 15107 12587 15113
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 12710 15104 12716 15156
rect 12768 15104 12774 15156
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 14274 15144 14280 15156
rect 12860 15116 14280 15144
rect 12860 15104 12866 15116
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 18417 15147 18475 15153
rect 18417 15113 18429 15147
rect 18463 15144 18475 15147
rect 18690 15144 18696 15156
rect 18463 15116 18696 15144
rect 18463 15113 18475 15116
rect 18417 15107 18475 15113
rect 12066 15076 12072 15088
rect 11348 15048 12072 15076
rect 11348 15008 11376 15048
rect 12066 15036 12072 15048
rect 12124 15036 12130 15088
rect 12728 15076 12756 15104
rect 13081 15079 13139 15085
rect 13081 15076 13093 15079
rect 12728 15048 13093 15076
rect 13081 15045 13093 15048
rect 13127 15045 13139 15079
rect 13081 15039 13139 15045
rect 12802 15008 12808 15020
rect 11256 14980 11376 15008
rect 11716 14980 12808 15008
rect 9677 14943 9735 14949
rect 9677 14940 9689 14943
rect 9640 14912 9689 14940
rect 9640 14900 9646 14912
rect 9677 14909 9689 14912
rect 9723 14909 9735 14943
rect 9677 14903 9735 14909
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 10686 14940 10692 14952
rect 9815 14912 10692 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 9692 14872 9720 14903
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 11054 14900 11060 14952
rect 11112 14949 11118 14952
rect 11112 14940 11124 14949
rect 11112 14912 11157 14940
rect 11112 14903 11124 14912
rect 11112 14900 11118 14903
rect 11256 14872 11284 14980
rect 11716 14949 11744 14980
rect 12802 14968 12808 14980
rect 12860 14968 12866 15020
rect 12912 14980 13952 15008
rect 11333 14943 11391 14949
rect 11333 14909 11345 14943
rect 11379 14909 11391 14943
rect 11333 14903 11391 14909
rect 11701 14943 11759 14949
rect 11701 14909 11713 14943
rect 11747 14909 11759 14943
rect 11701 14903 11759 14909
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 12526 14940 12532 14952
rect 12207 14912 12532 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 8956 14844 9628 14872
rect 9692 14844 11284 14872
rect 11348 14872 11376 14903
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 12912 14949 12940 14980
rect 12621 14943 12679 14949
rect 12621 14909 12633 14943
rect 12667 14934 12679 14943
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12728 14934 12909 14940
rect 12667 14912 12909 14934
rect 12667 14909 12756 14912
rect 12621 14906 12756 14909
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12621 14903 12679 14906
rect 12897 14903 12955 14909
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13219 14912 13308 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 11348 14844 12572 14872
rect 8849 14835 8907 14841
rect 9600 14816 9628 14844
rect 12544 14816 12572 14844
rect 13280 14816 13308 14912
rect 13924 14884 13952 14980
rect 14274 14900 14280 14952
rect 14332 14900 14338 14952
rect 14921 14943 14979 14949
rect 14921 14940 14933 14943
rect 14476 14912 14933 14940
rect 13906 14832 13912 14884
rect 13964 14832 13970 14884
rect 6457 14807 6515 14813
rect 6457 14804 6469 14807
rect 6420 14776 6469 14804
rect 6420 14764 6426 14776
rect 6457 14773 6469 14776
rect 6503 14773 6515 14807
rect 6457 14767 6515 14773
rect 7193 14807 7251 14813
rect 7193 14773 7205 14807
rect 7239 14804 7251 14807
rect 7374 14804 7380 14816
rect 7239 14776 7380 14804
rect 7239 14773 7251 14776
rect 7193 14767 7251 14773
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 8573 14807 8631 14813
rect 8573 14773 8585 14807
rect 8619 14804 8631 14807
rect 8938 14804 8944 14816
rect 8619 14776 8944 14804
rect 8619 14773 8631 14776
rect 8573 14767 8631 14773
rect 8938 14764 8944 14776
rect 8996 14804 9002 14816
rect 9401 14807 9459 14813
rect 9401 14804 9413 14807
rect 8996 14776 9413 14804
rect 8996 14764 9002 14776
rect 9401 14773 9413 14776
rect 9447 14773 9459 14807
rect 9401 14767 9459 14773
rect 9582 14764 9588 14816
rect 9640 14764 9646 14816
rect 9953 14807 10011 14813
rect 9953 14773 9965 14807
rect 9999 14804 10011 14807
rect 10594 14804 10600 14816
rect 9999 14776 10600 14804
rect 9999 14773 10011 14776
rect 9953 14767 10011 14773
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 11606 14764 11612 14816
rect 11664 14764 11670 14816
rect 12066 14764 12072 14816
rect 12124 14764 12130 14816
rect 12526 14764 12532 14816
rect 12584 14764 12590 14816
rect 12805 14807 12863 14813
rect 12805 14773 12817 14807
rect 12851 14804 12863 14807
rect 13262 14804 13268 14816
rect 12851 14776 13268 14804
rect 12851 14773 12863 14776
rect 12805 14767 12863 14773
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13541 14807 13599 14813
rect 13541 14773 13553 14807
rect 13587 14804 13599 14807
rect 13998 14804 14004 14816
rect 13587 14776 14004 14804
rect 13587 14773 13599 14776
rect 13541 14767 13599 14773
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 14292 14804 14320 14900
rect 14476 14884 14504 14912
rect 14921 14909 14933 14912
rect 14967 14940 14979 14943
rect 15013 14943 15071 14949
rect 15013 14940 15025 14943
rect 14967 14912 15025 14940
rect 14967 14909 14979 14912
rect 14921 14903 14979 14909
rect 15013 14909 15025 14912
rect 15059 14909 15071 14943
rect 15013 14903 15071 14909
rect 15102 14900 15108 14952
rect 15160 14940 15166 14952
rect 15269 14943 15327 14949
rect 15269 14940 15281 14943
rect 15160 14912 15281 14940
rect 15160 14900 15166 14912
rect 15269 14909 15281 14912
rect 15315 14909 15327 14943
rect 15269 14903 15327 14909
rect 17586 14900 17592 14952
rect 17644 14949 17650 14952
rect 17644 14903 17656 14949
rect 17644 14900 17650 14903
rect 17770 14900 17776 14952
rect 17828 14940 17834 14952
rect 17865 14943 17923 14949
rect 17865 14940 17877 14943
rect 17828 14912 17877 14940
rect 17828 14900 17834 14912
rect 17865 14909 17877 14912
rect 17911 14909 17923 14943
rect 17865 14903 17923 14909
rect 18141 14943 18199 14949
rect 18141 14909 18153 14943
rect 18187 14940 18199 14943
rect 18432 14940 18460 15107
rect 18690 15104 18696 15116
rect 18748 15104 18754 15156
rect 18874 15104 18880 15156
rect 18932 15144 18938 15156
rect 18969 15147 19027 15153
rect 18969 15144 18981 15147
rect 18932 15116 18981 15144
rect 18932 15104 18938 15116
rect 18969 15113 18981 15116
rect 19015 15113 19027 15147
rect 18969 15107 19027 15113
rect 18187 14912 18460 14940
rect 18509 14943 18567 14949
rect 18187 14909 18199 14912
rect 18141 14903 18199 14909
rect 18509 14909 18521 14943
rect 18555 14940 18567 14943
rect 18877 14943 18935 14949
rect 18555 14912 18644 14940
rect 18555 14909 18567 14912
rect 18509 14903 18567 14909
rect 18616 14884 18644 14912
rect 18877 14909 18889 14943
rect 18923 14940 18935 14943
rect 18966 14940 18972 14952
rect 18923 14912 18972 14940
rect 18923 14909 18935 14912
rect 18877 14903 18935 14909
rect 18966 14900 18972 14912
rect 19024 14900 19030 14952
rect 14458 14832 14464 14884
rect 14516 14832 14522 14884
rect 14654 14875 14712 14881
rect 14654 14872 14666 14875
rect 14568 14844 14666 14872
rect 14568 14804 14596 14844
rect 14654 14841 14666 14844
rect 14700 14841 14712 14875
rect 14654 14835 14712 14841
rect 18598 14832 18604 14884
rect 18656 14832 18662 14884
rect 14292 14776 14596 14804
rect 16390 14764 16396 14816
rect 16448 14764 16454 14816
rect 16482 14764 16488 14816
rect 16540 14764 16546 14816
rect 18049 14807 18107 14813
rect 18049 14773 18061 14807
rect 18095 14804 18107 14807
rect 18230 14804 18236 14816
rect 18095 14776 18236 14804
rect 18095 14773 18107 14776
rect 18049 14767 18107 14773
rect 18230 14764 18236 14776
rect 18288 14804 18294 14816
rect 18690 14804 18696 14816
rect 18288 14776 18696 14804
rect 18288 14764 18294 14776
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 552 14714 19571 14736
rect 552 14662 5112 14714
rect 5164 14662 5176 14714
rect 5228 14662 5240 14714
rect 5292 14662 5304 14714
rect 5356 14662 5368 14714
rect 5420 14662 9827 14714
rect 9879 14662 9891 14714
rect 9943 14662 9955 14714
rect 10007 14662 10019 14714
rect 10071 14662 10083 14714
rect 10135 14662 14542 14714
rect 14594 14662 14606 14714
rect 14658 14662 14670 14714
rect 14722 14662 14734 14714
rect 14786 14662 14798 14714
rect 14850 14662 19257 14714
rect 19309 14662 19321 14714
rect 19373 14662 19385 14714
rect 19437 14662 19449 14714
rect 19501 14662 19513 14714
rect 19565 14662 19571 14714
rect 552 14640 19571 14662
rect 1121 14603 1179 14609
rect 1121 14569 1133 14603
rect 1167 14600 1179 14603
rect 1578 14600 1584 14612
rect 1167 14572 1584 14600
rect 1167 14569 1179 14572
rect 1121 14563 1179 14569
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 1673 14603 1731 14609
rect 1673 14569 1685 14603
rect 1719 14600 1731 14603
rect 2590 14600 2596 14612
rect 1719 14572 2596 14600
rect 1719 14569 1731 14572
rect 1673 14563 1731 14569
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 5902 14560 5908 14612
rect 5960 14560 5966 14612
rect 6181 14603 6239 14609
rect 6181 14569 6193 14603
rect 6227 14600 6239 14603
rect 6454 14600 6460 14612
rect 6227 14572 6460 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 2038 14532 2044 14544
rect 1228 14504 2044 14532
rect 1228 14473 1256 14504
rect 2038 14492 2044 14504
rect 2096 14492 2102 14544
rect 2866 14532 2872 14544
rect 2148 14504 2872 14532
rect 1213 14467 1271 14473
rect 1213 14433 1225 14467
rect 1259 14433 1271 14467
rect 1213 14427 1271 14433
rect 1489 14467 1547 14473
rect 1489 14433 1501 14467
rect 1535 14433 1547 14467
rect 1489 14427 1547 14433
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 1670 14464 1676 14476
rect 1627 14436 1676 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 1504 14328 1532 14427
rect 1670 14424 1676 14436
rect 1728 14424 1734 14476
rect 2056 14463 2084 14492
rect 2148 14473 2176 14504
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 2133 14467 2191 14473
rect 2041 14457 2099 14463
rect 2041 14423 2053 14457
rect 2087 14423 2099 14457
rect 2133 14433 2145 14467
rect 2179 14433 2191 14467
rect 2133 14427 2191 14433
rect 2222 14424 2228 14476
rect 2280 14464 2286 14476
rect 2389 14467 2447 14473
rect 2389 14464 2401 14467
rect 2280 14436 2401 14464
rect 2280 14424 2286 14436
rect 2389 14433 2401 14436
rect 2435 14433 2447 14467
rect 2389 14427 2447 14433
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 5997 14467 6055 14473
rect 5997 14464 6009 14467
rect 5960 14436 6009 14464
rect 5960 14424 5966 14436
rect 5997 14433 6009 14436
rect 6043 14464 6055 14467
rect 6196 14464 6224 14563
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 7558 14560 7564 14612
rect 7616 14560 7622 14612
rect 9582 14600 9588 14612
rect 7760 14572 9588 14600
rect 6043 14436 6224 14464
rect 6273 14467 6331 14473
rect 6043 14433 6055 14436
rect 5997 14427 6055 14433
rect 6273 14433 6285 14467
rect 6319 14464 6331 14467
rect 6365 14467 6423 14473
rect 6365 14464 6377 14467
rect 6319 14436 6377 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 6365 14433 6377 14436
rect 6411 14464 6423 14467
rect 6825 14467 6883 14473
rect 6411 14436 6684 14464
rect 6411 14433 6423 14436
rect 6365 14427 6423 14433
rect 2041 14417 2099 14423
rect 2240 14396 2268 14424
rect 2148 14368 2268 14396
rect 2148 14328 2176 14368
rect 1504 14300 2176 14328
rect 6270 14288 6276 14340
rect 6328 14328 6334 14340
rect 6457 14331 6515 14337
rect 6457 14328 6469 14331
rect 6328 14300 6469 14328
rect 6328 14288 6334 14300
rect 6457 14297 6469 14300
rect 6503 14297 6515 14331
rect 6457 14291 6515 14297
rect 6656 14272 6684 14436
rect 6825 14433 6837 14467
rect 6871 14464 6883 14467
rect 7101 14467 7159 14473
rect 6871 14436 7052 14464
rect 6871 14433 6883 14436
rect 6825 14427 6883 14433
rect 7024 14337 7052 14436
rect 7101 14433 7113 14467
rect 7147 14433 7159 14467
rect 7101 14427 7159 14433
rect 7377 14467 7435 14473
rect 7377 14433 7389 14467
rect 7423 14464 7435 14467
rect 7576 14464 7604 14560
rect 7760 14532 7788 14572
rect 9582 14560 9588 14572
rect 9640 14600 9646 14612
rect 10689 14603 10747 14609
rect 10689 14600 10701 14603
rect 9640 14572 10701 14600
rect 9640 14560 9646 14572
rect 10689 14569 10701 14572
rect 10735 14600 10747 14603
rect 12066 14600 12072 14612
rect 10735 14572 12072 14600
rect 10735 14569 10747 14572
rect 10689 14563 10747 14569
rect 12066 14560 12072 14572
rect 12124 14560 12130 14612
rect 15194 14600 15200 14612
rect 13372 14572 15200 14600
rect 7668 14504 7788 14532
rect 7668 14473 7696 14504
rect 7926 14492 7932 14544
rect 7984 14532 7990 14544
rect 8665 14535 8723 14541
rect 8665 14532 8677 14535
rect 7984 14504 8677 14532
rect 7984 14492 7990 14504
rect 8665 14501 8677 14504
rect 8711 14532 8723 14535
rect 11054 14532 11060 14544
rect 8711 14504 11060 14532
rect 8711 14501 8723 14504
rect 8665 14495 8723 14501
rect 11054 14492 11060 14504
rect 11112 14532 11118 14544
rect 13372 14541 13400 14572
rect 15194 14560 15200 14572
rect 15252 14560 15258 14612
rect 17405 14603 17463 14609
rect 17405 14569 17417 14603
rect 17451 14569 17463 14603
rect 17405 14563 17463 14569
rect 13357 14535 13415 14541
rect 13357 14532 13369 14535
rect 11112 14504 13369 14532
rect 11112 14492 11118 14504
rect 13357 14501 13369 14504
rect 13403 14501 13415 14535
rect 16393 14535 16451 14541
rect 13357 14495 13415 14501
rect 13648 14504 14504 14532
rect 7423 14436 7604 14464
rect 7653 14467 7711 14473
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 7653 14433 7665 14467
rect 7699 14433 7711 14467
rect 8846 14464 8852 14476
rect 7653 14427 7711 14433
rect 7760 14436 8852 14464
rect 7116 14396 7144 14427
rect 7760 14396 7788 14436
rect 8846 14424 8852 14436
rect 8904 14424 8910 14476
rect 9030 14473 9036 14476
rect 9024 14464 9036 14473
rect 8991 14436 9036 14464
rect 9024 14427 9036 14436
rect 9030 14424 9036 14427
rect 9088 14424 9094 14476
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 10686 14464 10692 14476
rect 10551 14436 10692 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 10781 14467 10839 14473
rect 10781 14433 10793 14467
rect 10827 14464 10839 14467
rect 11606 14464 11612 14476
rect 10827 14436 11612 14464
rect 10827 14433 10839 14436
rect 10781 14427 10839 14433
rect 7116 14368 7788 14396
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14396 7987 14399
rect 8386 14396 8392 14408
rect 7975 14368 8392 14396
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 8386 14356 8392 14368
rect 8444 14396 8450 14408
rect 8757 14399 8815 14405
rect 8757 14396 8769 14399
rect 8444 14368 8769 14396
rect 8444 14356 8450 14368
rect 8680 14340 8708 14368
rect 8757 14365 8769 14368
rect 8803 14365 8815 14399
rect 8757 14359 8815 14365
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14396 10471 14399
rect 10796 14396 10824 14427
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 12089 14467 12147 14473
rect 12089 14433 12101 14467
rect 12135 14464 12147 14467
rect 12250 14464 12256 14476
rect 12135 14436 12256 14464
rect 12135 14433 12147 14436
rect 12089 14427 12147 14433
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 13648 14473 13676 14504
rect 14476 14476 14504 14504
rect 16393 14501 16405 14535
rect 16439 14532 16451 14535
rect 17420 14532 17448 14563
rect 16439 14504 17448 14532
rect 16439 14501 16451 14504
rect 16393 14495 16451 14501
rect 18414 14492 18420 14544
rect 18472 14532 18478 14544
rect 18966 14532 18972 14544
rect 18472 14504 18972 14532
rect 18472 14492 18478 14504
rect 18966 14492 18972 14504
rect 19024 14492 19030 14544
rect 13906 14473 13912 14476
rect 13633 14467 13691 14473
rect 13633 14433 13645 14467
rect 13679 14433 13691 14467
rect 13633 14427 13691 14433
rect 13900 14427 13912 14473
rect 13964 14464 13970 14476
rect 14274 14464 14280 14476
rect 13964 14436 14280 14464
rect 13906 14424 13912 14427
rect 13964 14424 13970 14436
rect 14274 14424 14280 14436
rect 14332 14424 14338 14476
rect 14458 14424 14464 14476
rect 14516 14424 14522 14476
rect 15654 14424 15660 14476
rect 15712 14464 15718 14476
rect 16206 14464 16212 14476
rect 15712 14436 16212 14464
rect 15712 14424 15718 14436
rect 16206 14424 16212 14436
rect 16264 14464 16270 14476
rect 16301 14467 16359 14473
rect 16301 14464 16313 14467
rect 16264 14436 16313 14464
rect 16264 14424 16270 14436
rect 16301 14433 16313 14436
rect 16347 14433 16359 14467
rect 16301 14427 16359 14433
rect 16485 14467 16543 14473
rect 16485 14433 16497 14467
rect 16531 14433 16543 14467
rect 16485 14427 16543 14433
rect 10459 14368 10824 14396
rect 12345 14399 12403 14405
rect 10459 14365 10471 14368
rect 10413 14359 10471 14365
rect 12345 14365 12357 14399
rect 12391 14396 12403 14399
rect 12526 14396 12532 14408
rect 12391 14368 12532 14396
rect 12391 14365 12403 14368
rect 12345 14359 12403 14365
rect 7009 14331 7067 14337
rect 7009 14297 7021 14331
rect 7055 14328 7067 14331
rect 7834 14328 7840 14340
rect 7055 14300 7840 14328
rect 7055 14297 7067 14300
rect 7009 14291 7067 14297
rect 7834 14288 7840 14300
rect 7892 14288 7898 14340
rect 8662 14288 8668 14340
rect 8720 14288 8726 14340
rect 10428 14328 10456 14359
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 15470 14356 15476 14408
rect 15528 14396 15534 14408
rect 16114 14396 16120 14408
rect 15528 14368 16120 14396
rect 15528 14356 15534 14368
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 10060 14300 10456 14328
rect 1394 14220 1400 14272
rect 1452 14220 1458 14272
rect 1946 14220 1952 14272
rect 2004 14220 2010 14272
rect 3513 14263 3571 14269
rect 3513 14229 3525 14263
rect 3559 14260 3571 14263
rect 4430 14260 4436 14272
rect 3559 14232 4436 14260
rect 3559 14229 3571 14232
rect 3513 14223 3571 14229
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 6638 14220 6644 14272
rect 6696 14260 6702 14272
rect 6733 14263 6791 14269
rect 6733 14260 6745 14263
rect 6696 14232 6745 14260
rect 6696 14220 6702 14232
rect 6733 14229 6745 14232
rect 6779 14229 6791 14263
rect 6733 14223 6791 14229
rect 7282 14220 7288 14272
rect 7340 14220 7346 14272
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 8570 14260 8576 14272
rect 7607 14232 8576 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 10060 14260 10088 14300
rect 15930 14288 15936 14340
rect 15988 14328 15994 14340
rect 16500 14328 16528 14427
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 16669 14467 16727 14473
rect 16669 14464 16681 14467
rect 16632 14436 16681 14464
rect 16632 14424 16638 14436
rect 16669 14433 16681 14436
rect 16715 14433 16727 14467
rect 16669 14427 16727 14433
rect 18529 14467 18587 14473
rect 18529 14433 18541 14467
rect 18575 14464 18587 14467
rect 18690 14464 18696 14476
rect 18575 14436 18696 14464
rect 18575 14433 18587 14436
rect 18529 14427 18587 14433
rect 18690 14424 18696 14436
rect 18748 14424 18754 14476
rect 18874 14424 18880 14476
rect 18932 14424 18938 14476
rect 18785 14399 18843 14405
rect 18785 14365 18797 14399
rect 18831 14365 18843 14399
rect 18785 14359 18843 14365
rect 15988 14300 16528 14328
rect 15988 14288 15994 14300
rect 9180 14232 10088 14260
rect 10137 14263 10195 14269
rect 9180 14220 9186 14232
rect 10137 14229 10149 14263
rect 10183 14260 10195 14263
rect 10226 14260 10232 14272
rect 10183 14232 10232 14260
rect 10183 14229 10195 14232
rect 10137 14223 10195 14229
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 10965 14263 11023 14269
rect 10965 14229 10977 14263
rect 11011 14260 11023 14263
rect 11330 14260 11336 14272
rect 11011 14232 11336 14260
rect 11011 14229 11023 14232
rect 10965 14223 11023 14229
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 15010 14220 15016 14272
rect 15068 14220 15074 14272
rect 16114 14220 16120 14272
rect 16172 14220 16178 14272
rect 18506 14220 18512 14272
rect 18564 14260 18570 14272
rect 18800 14260 18828 14359
rect 18564 14232 18828 14260
rect 18564 14220 18570 14232
rect 552 14170 19412 14192
rect 552 14118 2755 14170
rect 2807 14118 2819 14170
rect 2871 14118 2883 14170
rect 2935 14118 2947 14170
rect 2999 14118 3011 14170
rect 3063 14118 7470 14170
rect 7522 14118 7534 14170
rect 7586 14118 7598 14170
rect 7650 14118 7662 14170
rect 7714 14118 7726 14170
rect 7778 14118 12185 14170
rect 12237 14118 12249 14170
rect 12301 14118 12313 14170
rect 12365 14118 12377 14170
rect 12429 14118 12441 14170
rect 12493 14118 16900 14170
rect 16952 14118 16964 14170
rect 17016 14118 17028 14170
rect 17080 14118 17092 14170
rect 17144 14118 17156 14170
rect 17208 14118 19412 14170
rect 552 14096 19412 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 1581 14059 1639 14065
rect 1581 14056 1593 14059
rect 1452 14028 1593 14056
rect 1452 14016 1458 14028
rect 1581 14025 1593 14028
rect 1627 14056 1639 14059
rect 1762 14056 1768 14068
rect 1627 14028 1768 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 1857 14059 1915 14065
rect 1857 14025 1869 14059
rect 1903 14056 1915 14059
rect 1946 14056 1952 14068
rect 1903 14028 1952 14056
rect 1903 14025 1915 14028
rect 1857 14019 1915 14025
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2590 14016 2596 14068
rect 2648 14016 2654 14068
rect 5077 14059 5135 14065
rect 5077 14025 5089 14059
rect 5123 14056 5135 14059
rect 6546 14056 6552 14068
rect 5123 14028 6552 14056
rect 5123 14025 5135 14028
rect 5077 14019 5135 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 8021 14059 8079 14065
rect 8021 14056 8033 14059
rect 7892 14028 8033 14056
rect 7892 14016 7898 14028
rect 8021 14025 8033 14028
rect 8067 14025 8079 14059
rect 8021 14019 8079 14025
rect 12710 14016 12716 14068
rect 12768 14016 12774 14068
rect 12986 14016 12992 14068
rect 13044 14056 13050 14068
rect 13081 14059 13139 14065
rect 13081 14056 13093 14059
rect 13044 14028 13093 14056
rect 13044 14016 13050 14028
rect 13081 14025 13093 14028
rect 13127 14025 13139 14059
rect 13081 14019 13139 14025
rect 2608 13988 2636 14016
rect 1688 13960 2636 13988
rect 1578 13812 1584 13864
rect 1636 13812 1642 13864
rect 1688 13861 1716 13960
rect 2130 13880 2136 13932
rect 2188 13920 2194 13932
rect 2608 13920 2636 13960
rect 7742 13948 7748 14000
rect 7800 13988 7806 14000
rect 8202 13988 8208 14000
rect 7800 13960 8208 13988
rect 7800 13948 7806 13960
rect 8202 13948 8208 13960
rect 8260 13988 8266 14000
rect 8757 13991 8815 13997
rect 8757 13988 8769 13991
rect 8260 13960 8769 13988
rect 8260 13948 8266 13960
rect 8757 13957 8769 13960
rect 8803 13988 8815 13991
rect 9033 13991 9091 13997
rect 9033 13988 9045 13991
rect 8803 13960 9045 13988
rect 8803 13957 8815 13960
rect 8757 13951 8815 13957
rect 9033 13957 9045 13960
rect 9079 13957 9091 13991
rect 9033 13951 9091 13957
rect 2188 13892 2544 13920
rect 2608 13892 2820 13920
rect 2188 13880 2194 13892
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13821 1731 13855
rect 1673 13815 1731 13821
rect 1762 13812 1768 13864
rect 1820 13812 1826 13864
rect 2516 13861 2544 13892
rect 2792 13861 2820 13892
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 3697 13923 3755 13929
rect 3697 13920 3709 13923
rect 3384 13892 3709 13920
rect 3384 13880 3390 13892
rect 3697 13889 3709 13892
rect 3743 13889 3755 13923
rect 3697 13883 3755 13889
rect 7282 13880 7288 13932
rect 7340 13920 7346 13932
rect 8938 13920 8944 13932
rect 7340 13892 7880 13920
rect 7340 13880 7346 13892
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 2777 13855 2835 13861
rect 2547 13824 2728 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 1596 13784 1624 13812
rect 2056 13784 2084 13815
rect 1596 13756 2084 13784
rect 2700 13784 2728 13824
rect 2777 13821 2789 13855
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13821 2927 13855
rect 3421 13855 3479 13861
rect 3421 13852 3433 13855
rect 2869 13815 2927 13821
rect 3160 13824 3433 13852
rect 2884 13784 2912 13815
rect 2700 13756 2912 13784
rect 3160 13728 3188 13824
rect 3421 13821 3433 13824
rect 3467 13821 3479 13855
rect 3421 13815 3479 13821
rect 5626 13812 5632 13864
rect 5684 13812 5690 13864
rect 5902 13861 5908 13864
rect 5896 13852 5908 13861
rect 5863 13824 5908 13852
rect 5896 13815 5908 13824
rect 5902 13812 5908 13815
rect 5960 13812 5966 13864
rect 7374 13812 7380 13864
rect 7432 13852 7438 13864
rect 7852 13861 7880 13892
rect 8864 13892 8944 13920
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7432 13824 7757 13852
rect 7432 13812 7438 13824
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8018 13852 8024 13864
rect 7883 13824 8024 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 8018 13812 8024 13824
rect 8076 13852 8082 13864
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 8076 13824 8125 13852
rect 8076 13812 8082 13824
rect 8113 13821 8125 13824
rect 8159 13852 8171 13855
rect 8481 13855 8539 13861
rect 8481 13852 8493 13855
rect 8159 13824 8493 13852
rect 8159 13821 8171 13824
rect 8113 13815 8171 13821
rect 8481 13821 8493 13824
rect 8527 13821 8539 13855
rect 8481 13815 8539 13821
rect 8570 13812 8576 13864
rect 8628 13812 8634 13864
rect 8864 13861 8892 13892
rect 8938 13880 8944 13892
rect 8996 13880 9002 13932
rect 13096 13920 13124 14019
rect 13262 14016 13268 14068
rect 13320 14056 13326 14068
rect 13909 14059 13967 14065
rect 13909 14056 13921 14059
rect 13320 14028 13921 14056
rect 13320 14016 13326 14028
rect 13909 14025 13921 14028
rect 13955 14025 13967 14059
rect 13909 14019 13967 14025
rect 15010 14016 15016 14068
rect 15068 14016 15074 14068
rect 16945 14059 17003 14065
rect 16945 14025 16957 14059
rect 16991 14056 17003 14059
rect 17402 14056 17408 14068
rect 16991 14028 17408 14056
rect 16991 14025 17003 14028
rect 16945 14019 17003 14025
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 18785 14059 18843 14065
rect 18785 14025 18797 14059
rect 18831 14056 18843 14059
rect 18874 14056 18880 14068
rect 18831 14028 18880 14056
rect 18831 14025 18843 14028
rect 18785 14019 18843 14025
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 13633 13923 13691 13929
rect 13096 13892 13584 13920
rect 8849 13855 8907 13861
rect 8849 13821 8861 13855
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 9122 13812 9128 13864
rect 9180 13812 9186 13864
rect 13556 13861 13584 13892
rect 13633 13889 13645 13923
rect 13679 13920 13691 13923
rect 14274 13920 14280 13932
rect 13679 13892 14280 13920
rect 13679 13889 13691 13892
rect 13633 13883 13691 13889
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 14458 13880 14464 13932
rect 14516 13880 14522 13932
rect 15028 13920 15056 14016
rect 15166 13960 15608 13988
rect 15166 13920 15194 13960
rect 15028 13892 15194 13920
rect 12805 13855 12863 13861
rect 12805 13821 12817 13855
rect 12851 13852 12863 13855
rect 13173 13855 13231 13861
rect 13173 13852 13185 13855
rect 12851 13824 13185 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 13173 13821 13185 13824
rect 13219 13821 13231 13855
rect 13173 13815 13231 13821
rect 13541 13855 13599 13861
rect 13541 13821 13553 13855
rect 13587 13821 13599 13855
rect 13541 13815 13599 13821
rect 13817 13855 13875 13861
rect 13817 13821 13829 13855
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 3234 13744 3240 13796
rect 3292 13784 3298 13796
rect 3942 13787 4000 13793
rect 3942 13784 3954 13787
rect 3292 13756 3954 13784
rect 3292 13744 3298 13756
rect 3942 13753 3954 13756
rect 3988 13753 4000 13787
rect 3942 13747 4000 13753
rect 6270 13744 6276 13796
rect 6328 13784 6334 13796
rect 13188 13784 13216 13815
rect 6328 13756 7696 13784
rect 13188 13756 13768 13784
rect 6328 13744 6334 13756
rect 7668 13728 7696 13756
rect 13740 13728 13768 13756
rect 13832 13728 13860 13815
rect 15010 13812 15016 13864
rect 15068 13852 15074 13864
rect 15068 13824 15148 13852
rect 15068 13812 15074 13824
rect 15120 13784 15148 13824
rect 15194 13812 15200 13864
rect 15252 13812 15258 13864
rect 15580 13861 15608 13960
rect 15473 13855 15531 13861
rect 15473 13821 15485 13855
rect 15519 13821 15531 13855
rect 15473 13815 15531 13821
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 15488 13784 15516 13815
rect 15654 13812 15660 13864
rect 15712 13812 15718 13864
rect 15841 13855 15899 13861
rect 15841 13821 15853 13855
rect 15887 13852 15899 13855
rect 16482 13852 16488 13864
rect 15887 13824 16488 13852
rect 15887 13821 15899 13824
rect 15841 13815 15899 13821
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 16577 13855 16635 13861
rect 16577 13821 16589 13855
rect 16623 13821 16635 13855
rect 16577 13815 16635 13821
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13852 17095 13855
rect 17083 13824 17356 13852
rect 17083 13821 17095 13824
rect 17037 13815 17095 13821
rect 15120 13756 15516 13784
rect 16206 13744 16212 13796
rect 16264 13784 16270 13796
rect 16592 13784 16620 13815
rect 16264 13756 16620 13784
rect 16264 13744 16270 13756
rect 2133 13719 2191 13725
rect 2133 13685 2145 13719
rect 2179 13716 2191 13719
rect 2409 13719 2467 13725
rect 2409 13716 2421 13719
rect 2179 13688 2421 13716
rect 2179 13685 2191 13688
rect 2133 13679 2191 13685
rect 2409 13685 2421 13688
rect 2455 13716 2467 13719
rect 2498 13716 2504 13728
rect 2455 13688 2504 13716
rect 2455 13685 2467 13688
rect 2409 13679 2467 13685
rect 2498 13676 2504 13688
rect 2556 13676 2562 13728
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 2685 13719 2743 13725
rect 2685 13716 2697 13719
rect 2648 13688 2697 13716
rect 2648 13676 2654 13688
rect 2685 13685 2697 13688
rect 2731 13685 2743 13719
rect 2685 13679 2743 13685
rect 2961 13719 3019 13725
rect 2961 13685 2973 13719
rect 3007 13716 3019 13719
rect 3142 13716 3148 13728
rect 3007 13688 3148 13716
rect 3007 13685 3019 13688
rect 2961 13679 3019 13685
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 3513 13719 3571 13725
rect 3513 13685 3525 13719
rect 3559 13716 3571 13719
rect 4522 13716 4528 13728
rect 3559 13688 4528 13716
rect 3559 13685 3571 13688
rect 3513 13679 3571 13685
rect 4522 13676 4528 13688
rect 4580 13676 4586 13728
rect 7006 13676 7012 13728
rect 7064 13676 7070 13728
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 9030 13716 9036 13728
rect 7708 13688 9036 13716
rect 7708 13676 7714 13688
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 13722 13676 13728 13728
rect 13780 13676 13786 13728
rect 13814 13676 13820 13728
rect 13872 13676 13878 13728
rect 15286 13676 15292 13728
rect 15344 13676 15350 13728
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 16485 13719 16543 13725
rect 16485 13716 16497 13719
rect 16080 13688 16497 13716
rect 16080 13676 16086 13688
rect 16485 13685 16497 13688
rect 16531 13685 16543 13719
rect 16485 13679 16543 13685
rect 16574 13676 16580 13728
rect 16632 13716 16638 13728
rect 17129 13719 17187 13725
rect 17129 13716 17141 13719
rect 16632 13688 17141 13716
rect 16632 13676 16638 13688
rect 17129 13685 17141 13688
rect 17175 13685 17187 13719
rect 17328 13716 17356 13824
rect 17420 13784 17448 14016
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 18506 13852 18512 13864
rect 17828 13824 18512 13852
rect 17828 13812 17834 13824
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 18598 13812 18604 13864
rect 18656 13852 18662 13864
rect 18693 13855 18751 13861
rect 18693 13852 18705 13855
rect 18656 13824 18705 13852
rect 18656 13812 18662 13824
rect 18693 13821 18705 13824
rect 18739 13852 18751 13855
rect 18739 13824 19012 13852
rect 18739 13821 18751 13824
rect 18693 13815 18751 13821
rect 18242 13787 18300 13793
rect 18242 13784 18254 13787
rect 17420 13756 18254 13784
rect 18242 13753 18254 13756
rect 18288 13753 18300 13787
rect 18242 13747 18300 13753
rect 18782 13744 18788 13796
rect 18840 13744 18846 13796
rect 18138 13716 18144 13728
rect 17328 13688 18144 13716
rect 17129 13679 17187 13685
rect 18138 13676 18144 13688
rect 18196 13716 18202 13728
rect 18800 13716 18828 13744
rect 18984 13728 19012 13824
rect 18196 13688 18828 13716
rect 18196 13676 18202 13688
rect 18966 13676 18972 13728
rect 19024 13676 19030 13728
rect 552 13626 19571 13648
rect 552 13574 5112 13626
rect 5164 13574 5176 13626
rect 5228 13574 5240 13626
rect 5292 13574 5304 13626
rect 5356 13574 5368 13626
rect 5420 13574 9827 13626
rect 9879 13574 9891 13626
rect 9943 13574 9955 13626
rect 10007 13574 10019 13626
rect 10071 13574 10083 13626
rect 10135 13574 14542 13626
rect 14594 13574 14606 13626
rect 14658 13574 14670 13626
rect 14722 13574 14734 13626
rect 14786 13574 14798 13626
rect 14850 13574 19257 13626
rect 19309 13574 19321 13626
rect 19373 13574 19385 13626
rect 19437 13574 19449 13626
rect 19501 13574 19513 13626
rect 19565 13574 19571 13626
rect 552 13552 19571 13574
rect 5629 13515 5687 13521
rect 5629 13481 5641 13515
rect 5675 13512 5687 13515
rect 6086 13512 6092 13524
rect 5675 13484 6092 13512
rect 5675 13481 5687 13484
rect 5629 13475 5687 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 13814 13512 13820 13524
rect 7432 13484 12848 13512
rect 7432 13472 7438 13484
rect 1388 13447 1446 13453
rect 1388 13413 1400 13447
rect 1434 13444 1446 13447
rect 1578 13444 1584 13456
rect 1434 13416 1584 13444
rect 1434 13413 1446 13416
rect 1388 13407 1446 13413
rect 1578 13404 1584 13416
rect 1636 13404 1642 13456
rect 3234 13404 3240 13456
rect 3292 13404 3298 13456
rect 3326 13404 3332 13456
rect 3384 13404 3390 13456
rect 4154 13404 4160 13456
rect 4212 13444 4218 13456
rect 6457 13447 6515 13453
rect 6457 13444 6469 13447
rect 4212 13416 6469 13444
rect 4212 13404 4218 13416
rect 6457 13413 6469 13416
rect 6503 13444 6515 13447
rect 7926 13444 7932 13456
rect 6503 13416 7932 13444
rect 6503 13413 6515 13416
rect 6457 13407 6515 13413
rect 7926 13404 7932 13416
rect 7984 13404 7990 13456
rect 8570 13404 8576 13456
rect 8628 13444 8634 13456
rect 8910 13447 8968 13453
rect 8910 13444 8922 13447
rect 8628 13416 8922 13444
rect 8628 13404 8634 13416
rect 8910 13413 8922 13416
rect 8956 13413 8968 13447
rect 8910 13407 8968 13413
rect 12100 13447 12158 13453
rect 12100 13413 12112 13447
rect 12146 13444 12158 13447
rect 12710 13444 12716 13456
rect 12146 13416 12716 13444
rect 12146 13413 12158 13416
rect 12100 13407 12158 13413
rect 12710 13404 12716 13416
rect 12768 13404 12774 13456
rect 1121 13379 1179 13385
rect 1121 13345 1133 13379
rect 1167 13376 1179 13379
rect 1210 13376 1216 13388
rect 1167 13348 1216 13376
rect 1167 13345 1179 13348
rect 1121 13339 1179 13345
rect 1210 13336 1216 13348
rect 1268 13336 1274 13388
rect 2498 13336 2504 13388
rect 2556 13376 2562 13388
rect 2869 13379 2927 13385
rect 2869 13376 2881 13379
rect 2556 13348 2881 13376
rect 2556 13336 2562 13348
rect 2869 13345 2881 13348
rect 2915 13376 2927 13379
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 2915 13348 3157 13376
rect 2915 13345 2927 13348
rect 2869 13339 2927 13345
rect 3145 13345 3157 13348
rect 3191 13376 3203 13379
rect 3252 13376 3280 13404
rect 4522 13385 4528 13388
rect 4516 13376 4528 13385
rect 3191 13348 3280 13376
rect 3344 13348 4528 13376
rect 3191 13345 3203 13348
rect 3145 13339 3203 13345
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 3234 13308 3240 13320
rect 3099 13280 3240 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 3234 13268 3240 13280
rect 3292 13308 3298 13320
rect 3344 13308 3372 13348
rect 4516 13339 4528 13348
rect 4522 13336 4528 13339
rect 4580 13336 4586 13388
rect 4890 13336 4896 13388
rect 4948 13376 4954 13388
rect 5997 13379 6055 13385
rect 5997 13376 6009 13379
rect 4948 13348 6009 13376
rect 4948 13336 4954 13348
rect 5997 13345 6009 13348
rect 6043 13345 6055 13379
rect 5997 13339 6055 13345
rect 3292 13280 3372 13308
rect 3292 13268 3298 13280
rect 4246 13268 4252 13320
rect 4304 13268 4310 13320
rect 6012 13308 6040 13339
rect 6086 13336 6092 13388
rect 6144 13336 6150 13388
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13376 6239 13379
rect 6270 13376 6276 13388
rect 6227 13348 6276 13376
rect 6227 13345 6239 13348
rect 6181 13339 6239 13345
rect 6270 13336 6276 13348
rect 6328 13336 6334 13388
rect 6362 13336 6368 13388
rect 6420 13336 6426 13388
rect 6546 13336 6552 13388
rect 6604 13336 6610 13388
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7064 13348 7481 13376
rect 7064 13336 7070 13348
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 7650 13336 7656 13388
rect 7708 13336 7714 13388
rect 7745 13379 7803 13385
rect 7745 13345 7757 13379
rect 7791 13345 7803 13379
rect 7745 13339 7803 13345
rect 7837 13379 7895 13385
rect 7837 13345 7849 13379
rect 7883 13345 7895 13379
rect 7837 13339 7895 13345
rect 6012 13280 6500 13308
rect 2501 13243 2559 13249
rect 2501 13209 2513 13243
rect 2547 13240 2559 13243
rect 3510 13240 3516 13252
rect 2547 13212 3516 13240
rect 2547 13209 2559 13212
rect 2501 13203 2559 13209
rect 3510 13200 3516 13212
rect 3568 13200 3574 13252
rect 2590 13132 2596 13184
rect 2648 13172 2654 13184
rect 2777 13175 2835 13181
rect 2777 13172 2789 13175
rect 2648 13144 2789 13172
rect 2648 13132 2654 13144
rect 2777 13141 2789 13144
rect 2823 13141 2835 13175
rect 2777 13135 2835 13141
rect 5813 13175 5871 13181
rect 5813 13141 5825 13175
rect 5859 13172 5871 13175
rect 6362 13172 6368 13184
rect 5859 13144 6368 13172
rect 5859 13141 5871 13144
rect 5813 13135 5871 13141
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 6472 13172 6500 13280
rect 6564 13240 6592 13336
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 6788 13280 7205 13308
rect 6788 13268 6794 13280
rect 7193 13277 7205 13280
rect 7239 13277 7251 13311
rect 7193 13271 7251 13277
rect 7760 13240 7788 13339
rect 6564 13212 7788 13240
rect 7852 13308 7880 13339
rect 8662 13336 8668 13388
rect 8720 13336 8726 13388
rect 10594 13376 10600 13388
rect 8772 13348 10600 13376
rect 8772 13308 8800 13348
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 7852 13280 8800 13308
rect 12345 13311 12403 13317
rect 7852 13172 7880 13280
rect 12345 13277 12357 13311
rect 12391 13308 12403 13311
rect 12526 13308 12532 13320
rect 12391 13280 12532 13308
rect 12391 13277 12403 13280
rect 12345 13271 12403 13277
rect 12526 13268 12532 13280
rect 12584 13268 12590 13320
rect 6472 13144 7880 13172
rect 8021 13175 8079 13181
rect 8021 13141 8033 13175
rect 8067 13172 8079 13175
rect 8570 13172 8576 13184
rect 8067 13144 8576 13172
rect 8067 13141 8079 13144
rect 8021 13135 8079 13141
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 10042 13132 10048 13184
rect 10100 13132 10106 13184
rect 10962 13132 10968 13184
rect 11020 13132 11026 13184
rect 12820 13172 12848 13484
rect 13188 13484 13820 13512
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13376 13047 13379
rect 13078 13376 13084 13388
rect 13035 13348 13084 13376
rect 13035 13345 13047 13348
rect 12989 13339 13047 13345
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13308 12955 13311
rect 13188 13308 13216 13484
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 14274 13472 14280 13524
rect 14332 13472 14338 13524
rect 16114 13512 16120 13524
rect 14384 13484 16120 13512
rect 13832 13444 13860 13472
rect 14384 13444 14412 13484
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 16206 13472 16212 13524
rect 16264 13512 16270 13524
rect 16264 13484 17540 13512
rect 16264 13472 16270 13484
rect 13280 13416 13768 13444
rect 13832 13416 13952 13444
rect 13280 13385 13308 13416
rect 13265 13379 13323 13385
rect 13265 13345 13277 13379
rect 13311 13345 13323 13379
rect 13265 13339 13323 13345
rect 13538 13336 13544 13388
rect 13596 13336 13602 13388
rect 13740 13376 13768 13416
rect 13814 13376 13820 13388
rect 13740 13348 13820 13376
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 13924 13385 13952 13416
rect 14016 13416 14412 13444
rect 13909 13379 13967 13385
rect 13909 13345 13921 13379
rect 13955 13345 13967 13379
rect 13909 13339 13967 13345
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 12943 13280 13461 13308
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 13449 13277 13461 13280
rect 13495 13277 13507 13311
rect 14016 13308 14044 13416
rect 15194 13404 15200 13456
rect 15252 13444 15258 13456
rect 16485 13447 16543 13453
rect 16485 13444 16497 13447
rect 15252 13416 16497 13444
rect 15252 13404 15258 13416
rect 16485 13413 16497 13416
rect 16531 13444 16543 13447
rect 17218 13444 17224 13456
rect 16531 13416 17224 13444
rect 16531 13413 16543 13416
rect 16485 13407 16543 13413
rect 17218 13404 17224 13416
rect 17276 13404 17282 13456
rect 17512 13453 17540 13484
rect 17497 13447 17555 13453
rect 17497 13413 17509 13447
rect 17543 13413 17555 13447
rect 17497 13407 17555 13413
rect 14369 13379 14427 13385
rect 14369 13345 14381 13379
rect 14415 13345 14427 13379
rect 14369 13339 14427 13345
rect 15677 13379 15735 13385
rect 15677 13345 15689 13379
rect 15723 13376 15735 13379
rect 16022 13376 16028 13388
rect 15723 13348 16028 13376
rect 15723 13345 15735 13348
rect 15677 13339 15735 13345
rect 13449 13271 13507 13277
rect 13556 13280 14044 13308
rect 12986 13200 12992 13252
rect 13044 13240 13050 13252
rect 13173 13243 13231 13249
rect 13173 13240 13185 13243
rect 13044 13212 13185 13240
rect 13044 13200 13050 13212
rect 13173 13209 13185 13212
rect 13219 13209 13231 13243
rect 13556 13240 13584 13280
rect 14384 13240 14412 13339
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13376 16359 13379
rect 18141 13379 18199 13385
rect 18141 13376 18153 13379
rect 16347 13348 18153 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 18141 13345 18153 13348
rect 18187 13376 18199 13379
rect 18325 13379 18383 13385
rect 18325 13376 18337 13379
rect 18187 13348 18337 13376
rect 18187 13345 18199 13348
rect 18141 13339 18199 13345
rect 18325 13345 18337 13348
rect 18371 13345 18383 13379
rect 18325 13339 18383 13345
rect 18598 13336 18604 13388
rect 18656 13336 18662 13388
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13308 15991 13311
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 15979 13280 17233 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 17221 13277 17233 13280
rect 17267 13308 17279 13311
rect 17770 13308 17776 13320
rect 17267 13280 17776 13308
rect 17267 13277 17279 13280
rect 17221 13271 17279 13277
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 13173 13203 13231 13209
rect 13280 13212 13584 13240
rect 13740 13212 14412 13240
rect 13280 13172 13308 13212
rect 12820 13144 13308 13172
rect 13354 13132 13360 13184
rect 13412 13172 13418 13184
rect 13740 13181 13768 13212
rect 13725 13175 13783 13181
rect 13725 13172 13737 13175
rect 13412 13144 13737 13172
rect 13412 13132 13418 13144
rect 13725 13141 13737 13144
rect 13771 13141 13783 13175
rect 13725 13135 13783 13141
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 14001 13175 14059 13181
rect 14001 13172 14013 13175
rect 13872 13144 14013 13172
rect 13872 13132 13878 13144
rect 14001 13141 14013 13144
rect 14047 13172 14059 13175
rect 14182 13172 14188 13184
rect 14047 13144 14188 13172
rect 14047 13141 14059 13144
rect 14001 13135 14059 13141
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 14550 13132 14556 13184
rect 14608 13132 14614 13184
rect 16209 13175 16267 13181
rect 16209 13141 16221 13175
rect 16255 13172 16267 13175
rect 16482 13172 16488 13184
rect 16255 13144 16488 13172
rect 16255 13141 16267 13144
rect 16209 13135 16267 13141
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 552 13082 19412 13104
rect 552 13030 2755 13082
rect 2807 13030 2819 13082
rect 2871 13030 2883 13082
rect 2935 13030 2947 13082
rect 2999 13030 3011 13082
rect 3063 13030 7470 13082
rect 7522 13030 7534 13082
rect 7586 13030 7598 13082
rect 7650 13030 7662 13082
rect 7714 13030 7726 13082
rect 7778 13030 12185 13082
rect 12237 13030 12249 13082
rect 12301 13030 12313 13082
rect 12365 13030 12377 13082
rect 12429 13030 12441 13082
rect 12493 13030 16900 13082
rect 16952 13030 16964 13082
rect 17016 13030 17028 13082
rect 17080 13030 17092 13082
rect 17144 13030 17156 13082
rect 17208 13030 19412 13082
rect 552 13008 19412 13030
rect 2961 12971 3019 12977
rect 2961 12937 2973 12971
rect 3007 12968 3019 12971
rect 3970 12968 3976 12980
rect 3007 12940 3976 12968
rect 3007 12937 3019 12940
rect 2961 12931 3019 12937
rect 3970 12928 3976 12940
rect 4028 12968 4034 12980
rect 4985 12971 5043 12977
rect 4985 12968 4997 12971
rect 4028 12940 4997 12968
rect 4028 12928 4034 12940
rect 4985 12937 4997 12940
rect 5031 12937 5043 12971
rect 5626 12968 5632 12980
rect 4985 12931 5043 12937
rect 5368 12940 5632 12968
rect 2590 12900 2596 12912
rect 2516 12872 2596 12900
rect 2516 12773 2544 12872
rect 2590 12860 2596 12872
rect 2648 12900 2654 12912
rect 2648 12872 3556 12900
rect 2648 12860 2654 12872
rect 3234 12832 3240 12844
rect 3068 12804 3240 12832
rect 3068 12773 3096 12804
rect 3234 12792 3240 12804
rect 3292 12792 3298 12844
rect 2501 12767 2559 12773
rect 2501 12733 2513 12767
rect 2547 12733 2559 12767
rect 2501 12727 2559 12733
rect 2593 12767 2651 12773
rect 2593 12733 2605 12767
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12733 3111 12767
rect 3053 12727 3111 12733
rect 3329 12767 3387 12773
rect 3329 12733 3341 12767
rect 3375 12733 3387 12767
rect 3329 12727 3387 12733
rect 2608 12696 2636 12727
rect 2516 12668 2636 12696
rect 2685 12699 2743 12705
rect 2516 12640 2544 12668
rect 2685 12665 2697 12699
rect 2731 12696 2743 12699
rect 3142 12696 3148 12708
rect 2731 12668 3148 12696
rect 2731 12665 2743 12668
rect 2685 12659 2743 12665
rect 3142 12656 3148 12668
rect 3200 12696 3206 12708
rect 3344 12696 3372 12727
rect 3200 12668 3372 12696
rect 3528 12696 3556 12872
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 4304 12804 4353 12832
rect 4304 12792 4310 12804
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 4706 12792 4712 12844
rect 4764 12832 4770 12844
rect 5368 12841 5396 12940
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 6917 12971 6975 12977
rect 6917 12968 6929 12971
rect 6880 12940 6929 12968
rect 6880 12928 6886 12940
rect 6917 12937 6929 12940
rect 6963 12937 6975 12971
rect 6917 12931 6975 12937
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 8021 12971 8079 12977
rect 7331 12940 7972 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 6733 12903 6791 12909
rect 6733 12869 6745 12903
rect 6779 12900 6791 12903
rect 7944 12900 7972 12940
rect 8021 12937 8033 12971
rect 8067 12968 8079 12971
rect 8110 12968 8116 12980
rect 8067 12940 8116 12968
rect 8067 12937 8079 12940
rect 8021 12931 8079 12937
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 10689 12971 10747 12977
rect 8864 12940 10180 12968
rect 8864 12900 8892 12940
rect 10152 12912 10180 12940
rect 10689 12937 10701 12971
rect 10735 12937 10747 12971
rect 10689 12931 10747 12937
rect 13265 12971 13323 12977
rect 13265 12937 13277 12971
rect 13311 12968 13323 12971
rect 13814 12968 13820 12980
rect 13311 12940 13820 12968
rect 13311 12937 13323 12940
rect 13265 12931 13323 12937
rect 6779 12872 7604 12900
rect 7944 12872 8892 12900
rect 8941 12903 8999 12909
rect 6779 12869 6791 12872
rect 6733 12863 6791 12869
rect 5353 12835 5411 12841
rect 4764 12804 5028 12832
rect 4764 12792 4770 12804
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12764 3663 12767
rect 4154 12764 4160 12776
rect 3651 12736 4160 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 4154 12724 4160 12736
rect 4212 12724 4218 12776
rect 4522 12724 4528 12776
rect 4580 12764 4586 12776
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4580 12736 4629 12764
rect 4580 12724 4586 12736
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4617 12727 4675 12733
rect 4724 12736 4905 12764
rect 4724 12696 4752 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 5000 12764 5028 12804
rect 5353 12801 5365 12835
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12832 7067 12835
rect 7374 12832 7380 12844
rect 7055 12804 7380 12832
rect 7055 12801 7067 12804
rect 7009 12795 7067 12801
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 5609 12767 5667 12773
rect 5609 12764 5621 12767
rect 5000 12736 5621 12764
rect 4893 12727 4951 12733
rect 5609 12733 5621 12736
rect 5655 12733 5667 12767
rect 5609 12727 5667 12733
rect 7098 12724 7104 12776
rect 7156 12724 7162 12776
rect 7576 12764 7604 12872
rect 8941 12869 8953 12903
rect 8987 12869 8999 12903
rect 8941 12863 8999 12869
rect 7929 12835 7987 12841
rect 7929 12801 7941 12835
rect 7975 12832 7987 12835
rect 8956 12832 8984 12863
rect 10042 12860 10048 12912
rect 10100 12860 10106 12912
rect 10134 12860 10140 12912
rect 10192 12860 10198 12912
rect 9306 12832 9312 12844
rect 7975 12804 8984 12832
rect 9131 12804 9312 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 7576 12736 7972 12764
rect 3528 12668 4752 12696
rect 4908 12668 5120 12696
rect 3200 12656 3206 12668
rect 2409 12631 2467 12637
rect 2409 12597 2421 12631
rect 2455 12628 2467 12631
rect 2498 12628 2504 12640
rect 2455 12600 2504 12628
rect 2455 12597 2467 12600
rect 2409 12591 2467 12597
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 3421 12631 3479 12637
rect 3421 12597 3433 12631
rect 3467 12628 3479 12631
rect 3878 12628 3884 12640
rect 3467 12600 3884 12628
rect 3467 12597 3479 12600
rect 3421 12591 3479 12597
rect 3878 12588 3884 12600
rect 3936 12588 3942 12640
rect 4246 12588 4252 12640
rect 4304 12628 4310 12640
rect 4908 12628 4936 12668
rect 4304 12600 4936 12628
rect 5092 12628 5120 12668
rect 5442 12656 5448 12708
rect 5500 12696 5506 12708
rect 6825 12699 6883 12705
rect 6825 12696 6837 12699
rect 5500 12668 6837 12696
rect 5500 12656 5506 12668
rect 6825 12665 6837 12668
rect 6871 12665 6883 12699
rect 7745 12699 7803 12705
rect 7745 12696 7757 12699
rect 6825 12659 6883 12665
rect 6932 12668 7757 12696
rect 6932 12628 6960 12668
rect 7745 12665 7757 12668
rect 7791 12665 7803 12699
rect 7944 12696 7972 12736
rect 8018 12724 8024 12776
rect 8076 12724 8082 12776
rect 8389 12767 8447 12773
rect 8389 12733 8401 12767
rect 8435 12733 8447 12767
rect 8389 12727 8447 12733
rect 8404 12696 8432 12727
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 9131 12764 9159 12804
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 10060 12832 10088 12860
rect 10410 12832 10416 12844
rect 9692 12804 10088 12832
rect 10152 12804 10416 12832
rect 8812 12736 9159 12764
rect 8812 12724 8818 12736
rect 9214 12724 9220 12776
rect 9272 12764 9278 12776
rect 9692 12773 9720 12804
rect 9401 12767 9459 12773
rect 9401 12764 9413 12767
rect 9272 12736 9413 12764
rect 9272 12724 9278 12736
rect 9401 12733 9413 12736
rect 9447 12733 9459 12767
rect 9401 12727 9459 12733
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12733 9735 12767
rect 9677 12727 9735 12733
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 10152 12764 10180 12804
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10704 12764 10732 12931
rect 12894 12860 12900 12912
rect 12952 12900 12958 12912
rect 13354 12900 13360 12912
rect 12952 12872 13360 12900
rect 12952 12860 12958 12872
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12832 10839 12835
rect 11146 12832 11152 12844
rect 10827 12804 11152 12832
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 13464 12832 13492 12940
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 13906 12928 13912 12980
rect 13964 12968 13970 12980
rect 14185 12971 14243 12977
rect 14185 12968 14197 12971
rect 13964 12940 14197 12968
rect 13964 12928 13970 12940
rect 14185 12937 14197 12940
rect 14231 12937 14243 12971
rect 14185 12931 14243 12937
rect 15381 12971 15439 12977
rect 15381 12937 15393 12971
rect 15427 12968 15439 12971
rect 17586 12968 17592 12980
rect 15427 12940 17592 12968
rect 15427 12937 15439 12940
rect 15381 12931 15439 12937
rect 17586 12928 17592 12940
rect 17644 12928 17650 12980
rect 18322 12928 18328 12980
rect 18380 12928 18386 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 18785 12971 18843 12977
rect 18785 12968 18797 12971
rect 18748 12940 18797 12968
rect 18748 12928 18754 12940
rect 18785 12937 18797 12940
rect 18831 12937 18843 12971
rect 18785 12931 18843 12937
rect 12912 12804 13492 12832
rect 13648 12872 14412 12900
rect 12912 12776 12940 12804
rect 9815 12736 10180 12764
rect 10244 12736 10732 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 7944 12668 8432 12696
rect 8573 12699 8631 12705
rect 7745 12659 7803 12665
rect 8573 12665 8585 12699
rect 8619 12665 8631 12699
rect 8573 12659 8631 12665
rect 5092 12600 6960 12628
rect 4304 12588 4310 12600
rect 8202 12588 8208 12640
rect 8260 12588 8266 12640
rect 8588 12628 8616 12659
rect 8662 12656 8668 12708
rect 8720 12656 8726 12708
rect 9585 12699 9643 12705
rect 9585 12665 9597 12699
rect 9631 12665 9643 12699
rect 9585 12659 9643 12665
rect 9490 12628 9496 12640
rect 8588 12600 9496 12628
rect 9490 12588 9496 12600
rect 9548 12628 9554 12640
rect 9600 12628 9628 12659
rect 9548 12600 9628 12628
rect 9953 12631 10011 12637
rect 9548 12588 9554 12600
rect 9953 12597 9965 12631
rect 9999 12628 10011 12631
rect 10244 12628 10272 12736
rect 10870 12724 10876 12776
rect 10928 12724 10934 12776
rect 12894 12724 12900 12776
rect 12952 12724 12958 12776
rect 13357 12767 13415 12773
rect 13357 12733 13369 12767
rect 13403 12764 13415 12767
rect 13538 12766 13544 12776
rect 13464 12764 13544 12766
rect 13403 12738 13544 12764
rect 13403 12736 13492 12738
rect 13403 12733 13415 12736
rect 13357 12727 13415 12733
rect 10321 12699 10379 12705
rect 10321 12665 10333 12699
rect 10367 12696 10379 12699
rect 10597 12699 10655 12705
rect 10597 12696 10609 12699
rect 10367 12668 10609 12696
rect 10367 12665 10379 12668
rect 10321 12659 10379 12665
rect 10597 12665 10609 12668
rect 10643 12696 10655 12699
rect 10686 12696 10692 12708
rect 10643 12668 10692 12696
rect 10643 12665 10655 12668
rect 10597 12659 10655 12665
rect 10686 12656 10692 12668
rect 10744 12656 10750 12708
rect 9999 12600 10272 12628
rect 11057 12631 11115 12637
rect 9999 12597 10011 12600
rect 9953 12591 10011 12597
rect 11057 12597 11069 12631
rect 11103 12628 11115 12631
rect 11606 12628 11612 12640
rect 11103 12600 11612 12628
rect 11103 12597 11115 12600
rect 11057 12591 11115 12597
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12066 12628 12072 12640
rect 11848 12600 12072 12628
rect 11848 12588 11854 12600
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 12986 12588 12992 12640
rect 13044 12588 13050 12640
rect 13464 12628 13492 12736
rect 13538 12724 13544 12738
rect 13596 12724 13602 12776
rect 13648 12764 13676 12872
rect 14384 12844 14412 12872
rect 14550 12860 14556 12912
rect 14608 12860 14614 12912
rect 14366 12792 14372 12844
rect 14424 12792 14430 12844
rect 14568 12832 14596 12860
rect 14737 12835 14795 12841
rect 14737 12832 14749 12835
rect 14568 12804 14749 12832
rect 14737 12801 14749 12804
rect 14783 12801 14795 12835
rect 14737 12795 14795 12801
rect 14918 12792 14924 12844
rect 14976 12792 14982 12844
rect 13725 12767 13783 12773
rect 13725 12764 13737 12767
rect 13648 12736 13737 12764
rect 13725 12733 13737 12736
rect 13771 12733 13783 12767
rect 13725 12727 13783 12733
rect 13814 12724 13820 12776
rect 13872 12724 13878 12776
rect 14274 12724 14280 12776
rect 14332 12724 14338 12776
rect 14458 12724 14464 12776
rect 14516 12764 14522 12776
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 14516 12736 14657 12764
rect 14516 12724 14522 12736
rect 14645 12733 14657 12736
rect 14691 12733 14703 12767
rect 14645 12727 14703 12733
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 14884 12736 15025 12764
rect 14884 12724 14890 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12733 17187 12767
rect 17129 12727 17187 12733
rect 16206 12656 16212 12708
rect 16264 12696 16270 12708
rect 16862 12699 16920 12705
rect 16862 12696 16874 12699
rect 16264 12668 16874 12696
rect 16264 12656 16270 12668
rect 16862 12665 16874 12668
rect 16908 12665 16920 12699
rect 17144 12696 17172 12727
rect 17218 12724 17224 12776
rect 17276 12724 17282 12776
rect 18414 12724 18420 12776
rect 18472 12724 18478 12776
rect 18874 12724 18880 12776
rect 18932 12724 18938 12776
rect 18049 12699 18107 12705
rect 18049 12696 18061 12699
rect 17144 12668 18061 12696
rect 16862 12659 16920 12665
rect 18049 12665 18061 12668
rect 18095 12696 18107 12699
rect 18095 12668 18920 12696
rect 18095 12665 18107 12668
rect 18049 12659 18107 12665
rect 18892 12640 18920 12668
rect 13633 12631 13691 12637
rect 13633 12628 13645 12631
rect 13464 12600 13645 12628
rect 13633 12597 13645 12600
rect 13679 12628 13691 12631
rect 13906 12628 13912 12640
rect 13679 12600 13912 12628
rect 13679 12597 13691 12600
rect 13633 12591 13691 12597
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 15746 12588 15752 12640
rect 15804 12588 15810 12640
rect 18874 12588 18880 12640
rect 18932 12588 18938 12640
rect 552 12538 19571 12560
rect 552 12486 5112 12538
rect 5164 12486 5176 12538
rect 5228 12486 5240 12538
rect 5292 12486 5304 12538
rect 5356 12486 5368 12538
rect 5420 12486 9827 12538
rect 9879 12486 9891 12538
rect 9943 12486 9955 12538
rect 10007 12486 10019 12538
rect 10071 12486 10083 12538
rect 10135 12486 14542 12538
rect 14594 12486 14606 12538
rect 14658 12486 14670 12538
rect 14722 12486 14734 12538
rect 14786 12486 14798 12538
rect 14850 12486 19257 12538
rect 19309 12486 19321 12538
rect 19373 12486 19385 12538
rect 19437 12486 19449 12538
rect 19501 12486 19513 12538
rect 19565 12486 19571 12538
rect 552 12464 19571 12486
rect 2317 12427 2375 12433
rect 2317 12393 2329 12427
rect 2363 12424 2375 12427
rect 3602 12424 3608 12436
rect 2363 12396 3188 12424
rect 2363 12393 2375 12396
rect 2317 12387 2375 12393
rect 1204 12359 1262 12365
rect 1204 12325 1216 12359
rect 1250 12356 1262 12359
rect 1302 12356 1308 12368
rect 1250 12328 1308 12356
rect 1250 12325 1262 12328
rect 1204 12319 1262 12325
rect 1302 12316 1308 12328
rect 1360 12316 1366 12368
rect 2406 12316 2412 12368
rect 2464 12356 2470 12368
rect 2869 12359 2927 12365
rect 2869 12356 2881 12359
rect 2464 12328 2881 12356
rect 2464 12316 2470 12328
rect 2869 12325 2881 12328
rect 2915 12325 2927 12359
rect 2869 12319 2927 12325
rect 2590 12248 2596 12300
rect 2648 12248 2654 12300
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 2961 12291 3019 12297
rect 2823 12260 2912 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 937 12223 995 12229
rect 937 12189 949 12223
rect 983 12189 995 12223
rect 937 12183 995 12189
rect 952 12084 980 12183
rect 1210 12084 1216 12096
rect 952 12056 1216 12084
rect 1210 12044 1216 12056
rect 1268 12044 1274 12096
rect 2406 12044 2412 12096
rect 2464 12084 2470 12096
rect 2884 12084 2912 12260
rect 2961 12257 2973 12291
rect 3007 12288 3019 12291
rect 3160 12288 3188 12396
rect 3436 12396 3608 12424
rect 3436 12297 3464 12396
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 3789 12427 3847 12433
rect 3789 12393 3801 12427
rect 3835 12424 3847 12427
rect 5442 12424 5448 12436
rect 3835 12396 5448 12424
rect 3835 12393 3847 12396
rect 3789 12387 3847 12393
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 7193 12427 7251 12433
rect 7193 12393 7205 12427
rect 7239 12424 7251 12427
rect 7239 12396 8340 12424
rect 7239 12393 7251 12396
rect 7193 12387 7251 12393
rect 3510 12316 3516 12368
rect 3568 12316 3574 12368
rect 3896 12328 4660 12356
rect 3896 12300 3924 12328
rect 3237 12291 3295 12297
rect 3237 12288 3249 12291
rect 3007 12260 3096 12288
rect 3160 12260 3249 12288
rect 3007 12257 3019 12260
rect 2961 12251 3019 12257
rect 3068 12220 3096 12260
rect 3237 12257 3249 12260
rect 3283 12257 3295 12291
rect 3237 12251 3295 12257
rect 3421 12291 3479 12297
rect 3421 12257 3433 12291
rect 3467 12257 3479 12291
rect 3421 12251 3479 12257
rect 3605 12291 3663 12297
rect 3605 12257 3617 12291
rect 3651 12257 3663 12291
rect 3605 12251 3663 12257
rect 3510 12220 3516 12232
rect 3068 12192 3516 12220
rect 3510 12180 3516 12192
rect 3568 12220 3574 12232
rect 3620 12220 3648 12251
rect 3878 12248 3884 12300
rect 3936 12248 3942 12300
rect 3970 12248 3976 12300
rect 4028 12288 4034 12300
rect 4632 12297 4660 12328
rect 4706 12316 4712 12368
rect 4764 12356 4770 12368
rect 5261 12359 5319 12365
rect 5261 12356 5273 12359
rect 4764 12328 5273 12356
rect 4764 12316 4770 12328
rect 5092 12300 5120 12328
rect 5261 12325 5273 12328
rect 5307 12325 5319 12359
rect 6730 12356 6736 12368
rect 5261 12319 5319 12325
rect 5828 12328 6736 12356
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 4028 12260 4077 12288
rect 4028 12248 4034 12260
rect 4065 12257 4077 12260
rect 4111 12288 4123 12291
rect 4249 12291 4307 12297
rect 4249 12288 4261 12291
rect 4111 12260 4261 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4249 12257 4261 12260
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 4617 12291 4675 12297
rect 4617 12257 4629 12291
rect 4663 12288 4675 12291
rect 4663 12260 5028 12288
rect 4663 12257 4675 12260
rect 4617 12251 4675 12257
rect 4890 12220 4896 12232
rect 3568 12192 4896 12220
rect 3568 12180 3574 12192
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 5000 12220 5028 12260
rect 5074 12248 5080 12300
rect 5132 12248 5138 12300
rect 5169 12291 5227 12297
rect 5169 12257 5181 12291
rect 5215 12257 5227 12291
rect 5169 12251 5227 12257
rect 5184 12220 5212 12251
rect 5626 12248 5632 12300
rect 5684 12288 5690 12300
rect 5828 12297 5856 12328
rect 6730 12316 6736 12328
rect 6788 12356 6794 12368
rect 6788 12328 7880 12356
rect 6788 12316 6794 12328
rect 7852 12300 7880 12328
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5684 12260 5825 12288
rect 5684 12248 5690 12260
rect 5813 12257 5825 12260
rect 5859 12257 5871 12291
rect 6069 12291 6127 12297
rect 6069 12288 6081 12291
rect 5813 12251 5871 12257
rect 5920 12260 6081 12288
rect 5920 12220 5948 12260
rect 6069 12257 6081 12260
rect 6115 12257 6127 12291
rect 6069 12251 6127 12257
rect 7834 12248 7840 12300
rect 7892 12248 7898 12300
rect 8093 12291 8151 12297
rect 8093 12288 8105 12291
rect 7944 12260 8105 12288
rect 5000 12192 5212 12220
rect 5644 12192 5948 12220
rect 3145 12155 3203 12161
rect 3145 12121 3157 12155
rect 3191 12152 3203 12155
rect 4246 12152 4252 12164
rect 3191 12124 4252 12152
rect 3191 12121 3203 12124
rect 3145 12115 3203 12121
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 4341 12155 4399 12161
rect 4341 12121 4353 12155
rect 4387 12152 4399 12155
rect 4430 12152 4436 12164
rect 4387 12124 4436 12152
rect 4387 12121 4399 12124
rect 4341 12115 4399 12121
rect 4430 12112 4436 12124
rect 4488 12152 4494 12164
rect 4985 12155 5043 12161
rect 4985 12152 4997 12155
rect 4488 12124 4997 12152
rect 4488 12112 4494 12124
rect 4985 12121 4997 12124
rect 5031 12121 5043 12155
rect 4985 12115 5043 12121
rect 3602 12084 3608 12096
rect 2464 12056 3608 12084
rect 2464 12044 2470 12056
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 3970 12044 3976 12096
rect 4028 12044 4034 12096
rect 4706 12044 4712 12096
rect 4764 12044 4770 12096
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5644 12084 5672 12192
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7944 12220 7972 12260
rect 8093 12257 8105 12260
rect 8139 12257 8151 12291
rect 8312 12288 8340 12396
rect 9214 12384 9220 12436
rect 9272 12384 9278 12436
rect 10781 12427 10839 12433
rect 10781 12393 10793 12427
rect 10827 12424 10839 12427
rect 10870 12424 10876 12436
rect 10827 12396 10876 12424
rect 10827 12393 10839 12396
rect 10781 12387 10839 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11624 12396 16712 12424
rect 9581 12359 9639 12365
rect 9581 12325 9593 12359
rect 9627 12356 9639 12359
rect 10318 12356 10324 12368
rect 9627 12328 10324 12356
rect 9627 12325 9639 12328
rect 9581 12319 9639 12325
rect 10318 12316 10324 12328
rect 10376 12316 10382 12368
rect 10502 12316 10508 12368
rect 10560 12316 10566 12368
rect 9490 12297 9496 12300
rect 9309 12291 9367 12297
rect 9447 12294 9496 12297
rect 9309 12288 9321 12291
rect 8312 12260 9321 12288
rect 8093 12251 8151 12257
rect 9309 12257 9321 12260
rect 9355 12257 9367 12291
rect 9416 12291 9496 12294
rect 9416 12260 9459 12291
rect 9309 12251 9367 12257
rect 9447 12257 9459 12260
rect 9493 12257 9496 12291
rect 9447 12251 9496 12257
rect 9490 12248 9496 12251
rect 9548 12248 9554 12300
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 7248 12192 7972 12220
rect 7248 12180 7254 12192
rect 9578 12180 9584 12232
rect 9636 12220 9642 12232
rect 9692 12220 9720 12251
rect 9766 12248 9772 12300
rect 9824 12288 9830 12300
rect 10229 12291 10287 12297
rect 10229 12288 10241 12291
rect 9824 12260 10241 12288
rect 9824 12248 9830 12260
rect 10229 12257 10241 12260
rect 10275 12257 10287 12291
rect 10413 12291 10471 12297
rect 10413 12288 10425 12291
rect 10229 12251 10287 12257
rect 10336 12260 10425 12288
rect 10336 12232 10364 12260
rect 10413 12257 10425 12260
rect 10459 12257 10471 12291
rect 10413 12251 10471 12257
rect 10597 12291 10655 12297
rect 10597 12257 10609 12291
rect 10643 12257 10655 12291
rect 11624 12288 11652 12396
rect 12526 12356 12532 12368
rect 12360 12328 12532 12356
rect 12360 12297 12388 12328
rect 12526 12316 12532 12328
rect 12584 12356 12590 12368
rect 12584 12328 13860 12356
rect 12584 12316 12590 12328
rect 10597 12251 10655 12257
rect 11348 12260 11652 12288
rect 12089 12291 12147 12297
rect 10042 12220 10048 12232
rect 9636 12192 10048 12220
rect 9636 12180 9642 12192
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10318 12180 10324 12232
rect 10376 12180 10382 12232
rect 10612 12220 10640 12251
rect 10778 12220 10784 12232
rect 10612 12192 10784 12220
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 11348 12152 11376 12260
rect 12089 12257 12101 12291
rect 12135 12288 12147 12291
rect 12345 12291 12403 12297
rect 12135 12260 12296 12288
rect 12135 12257 12147 12260
rect 12089 12251 12147 12257
rect 12268 12220 12296 12260
rect 12345 12257 12357 12291
rect 12391 12257 12403 12291
rect 12345 12251 12403 12257
rect 12802 12248 12808 12300
rect 12860 12248 12866 12300
rect 13832 12297 13860 12328
rect 14274 12316 14280 12368
rect 14332 12356 14338 12368
rect 16022 12356 16028 12368
rect 14332 12328 15056 12356
rect 14332 12316 14338 12328
rect 13561 12291 13619 12297
rect 13561 12257 13573 12291
rect 13607 12288 13619 12291
rect 13817 12291 13875 12297
rect 13607 12260 13768 12288
rect 13607 12257 13619 12260
rect 13561 12251 13619 12257
rect 12820 12220 12848 12248
rect 12268 12192 12848 12220
rect 13740 12220 13768 12260
rect 13817 12257 13829 12291
rect 13863 12257 13875 12291
rect 13817 12251 13875 12257
rect 14090 12248 14096 12300
rect 14148 12248 14154 12300
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 15028 12286 15056 12328
rect 15672 12328 16028 12356
rect 15672 12297 15700 12328
rect 16022 12316 16028 12328
rect 16080 12316 16086 12368
rect 15105 12291 15163 12297
rect 15105 12286 15117 12291
rect 15028 12258 15117 12286
rect 14921 12251 14979 12257
rect 15105 12257 15117 12258
rect 15151 12257 15163 12291
rect 15105 12251 15163 12257
rect 15565 12291 15623 12297
rect 15565 12257 15577 12291
rect 15611 12288 15623 12291
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15611 12260 15669 12288
rect 15611 12257 15623 12260
rect 15565 12251 15623 12257
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 14200 12220 14228 12251
rect 13740 12192 14228 12220
rect 14936 12220 14964 12251
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 16684 12297 16712 12396
rect 17586 12384 17592 12436
rect 17644 12384 17650 12436
rect 16117 12291 16175 12297
rect 16117 12288 16129 12291
rect 15804 12260 16129 12288
rect 15804 12248 15810 12260
rect 16117 12257 16129 12260
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 16301 12291 16359 12297
rect 16301 12257 16313 12291
rect 16347 12257 16359 12291
rect 16301 12251 16359 12257
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 16206 12220 16212 12232
rect 14936 12192 16212 12220
rect 8925 12124 11376 12152
rect 5718 12084 5724 12096
rect 4856 12056 5724 12084
rect 4856 12044 4862 12056
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8925 12084 8953 12124
rect 8260 12056 8953 12084
rect 9861 12087 9919 12093
rect 8260 12044 8266 12056
rect 9861 12053 9873 12087
rect 9907 12084 9919 12087
rect 10134 12084 10140 12096
rect 9907 12056 10140 12084
rect 9907 12053 9919 12056
rect 9861 12047 9919 12053
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 10965 12087 11023 12093
rect 10965 12053 10977 12087
rect 11011 12084 11023 12087
rect 11146 12084 11152 12096
rect 11011 12056 11152 12084
rect 11011 12053 11023 12056
rect 10965 12047 11023 12053
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 12437 12087 12495 12093
rect 12437 12053 12449 12087
rect 12483 12084 12495 12087
rect 12526 12084 12532 12096
rect 12483 12056 12532 12084
rect 12483 12053 12495 12056
rect 12437 12047 12495 12053
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 13630 12044 13636 12096
rect 13688 12084 13694 12096
rect 14016 12093 14044 12192
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 14366 12112 14372 12164
rect 14424 12152 14430 12164
rect 15197 12155 15255 12161
rect 15197 12152 15209 12155
rect 14424 12124 15209 12152
rect 14424 12112 14430 12124
rect 15197 12121 15209 12124
rect 15243 12121 15255 12155
rect 16316 12152 16344 12251
rect 17310 12248 17316 12300
rect 17368 12248 17374 12300
rect 18690 12288 18696 12300
rect 18748 12297 18754 12300
rect 18660 12260 18696 12288
rect 18690 12248 18696 12260
rect 18748 12251 18760 12297
rect 18748 12248 18754 12251
rect 18874 12248 18880 12300
rect 18932 12288 18938 12300
rect 18969 12291 19027 12297
rect 18969 12288 18981 12291
rect 18932 12260 18981 12288
rect 18932 12248 18938 12260
rect 18969 12257 18981 12260
rect 19015 12257 19027 12291
rect 18969 12251 19027 12257
rect 16574 12180 16580 12232
rect 16632 12180 16638 12232
rect 15197 12115 15255 12121
rect 15856 12124 16344 12152
rect 15856 12096 15884 12124
rect 14001 12087 14059 12093
rect 14001 12084 14013 12087
rect 13688 12056 14013 12084
rect 13688 12044 13694 12056
rect 14001 12053 14013 12056
rect 14047 12053 14059 12087
rect 14001 12047 14059 12053
rect 14921 12087 14979 12093
rect 14921 12053 14933 12087
rect 14967 12084 14979 12087
rect 15102 12084 15108 12096
rect 14967 12056 15108 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 15102 12044 15108 12056
rect 15160 12044 15166 12096
rect 15473 12087 15531 12093
rect 15473 12053 15485 12087
rect 15519 12084 15531 12087
rect 15654 12084 15660 12096
rect 15519 12056 15660 12084
rect 15519 12053 15531 12056
rect 15473 12047 15531 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 15746 12044 15752 12096
rect 15804 12044 15810 12096
rect 15838 12044 15844 12096
rect 15896 12044 15902 12096
rect 552 11994 19412 12016
rect 552 11942 2755 11994
rect 2807 11942 2819 11994
rect 2871 11942 2883 11994
rect 2935 11942 2947 11994
rect 2999 11942 3011 11994
rect 3063 11942 7470 11994
rect 7522 11942 7534 11994
rect 7586 11942 7598 11994
rect 7650 11942 7662 11994
rect 7714 11942 7726 11994
rect 7778 11942 12185 11994
rect 12237 11942 12249 11994
rect 12301 11942 12313 11994
rect 12365 11942 12377 11994
rect 12429 11942 12441 11994
rect 12493 11942 16900 11994
rect 16952 11942 16964 11994
rect 17016 11942 17028 11994
rect 17080 11942 17092 11994
rect 17144 11942 17156 11994
rect 17208 11942 19412 11994
rect 552 11920 19412 11942
rect 2409 11883 2467 11889
rect 2409 11849 2421 11883
rect 2455 11880 2467 11883
rect 2590 11880 2596 11892
rect 2455 11852 2596 11880
rect 2455 11849 2467 11852
rect 2409 11843 2467 11849
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 3878 11840 3884 11892
rect 3936 11840 3942 11892
rect 10965 11883 11023 11889
rect 10965 11849 10977 11883
rect 11011 11880 11023 11883
rect 11238 11880 11244 11892
rect 11011 11852 11244 11880
rect 11011 11849 11023 11852
rect 10965 11843 11023 11849
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 11698 11840 11704 11892
rect 11756 11840 11762 11892
rect 12526 11840 12532 11892
rect 12584 11840 12590 11892
rect 12805 11883 12863 11889
rect 12805 11849 12817 11883
rect 12851 11880 12863 11883
rect 12894 11880 12900 11892
rect 12851 11852 12900 11880
rect 12851 11849 12863 11852
rect 12805 11843 12863 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 13906 11840 13912 11892
rect 13964 11840 13970 11892
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 14553 11883 14611 11889
rect 14553 11880 14565 11883
rect 14332 11852 14565 11880
rect 14332 11840 14338 11852
rect 14553 11849 14565 11852
rect 14599 11849 14611 11883
rect 14553 11843 14611 11849
rect 16022 11840 16028 11892
rect 16080 11880 16086 11892
rect 16485 11883 16543 11889
rect 16485 11880 16497 11883
rect 16080 11852 16497 11880
rect 16080 11840 16086 11852
rect 16485 11849 16497 11852
rect 16531 11849 16543 11883
rect 16485 11843 16543 11849
rect 18414 11840 18420 11892
rect 18472 11840 18478 11892
rect 18782 11840 18788 11892
rect 18840 11840 18846 11892
rect 2498 11772 2504 11824
rect 2556 11772 2562 11824
rect 4706 11772 4712 11824
rect 4764 11812 4770 11824
rect 11333 11815 11391 11821
rect 4764 11784 6040 11812
rect 4764 11772 4770 11784
rect 2516 11744 2544 11772
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 2516 11716 2605 11744
rect 2593 11713 2605 11716
rect 2639 11744 2651 11747
rect 2639 11716 2774 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 1029 11679 1087 11685
rect 1029 11645 1041 11679
rect 1075 11676 1087 11679
rect 1075 11648 1256 11676
rect 1075 11645 1087 11648
rect 1029 11639 1087 11645
rect 1228 11552 1256 11648
rect 1762 11636 1768 11688
rect 1820 11676 1826 11688
rect 2501 11679 2559 11685
rect 2501 11676 2513 11679
rect 1820 11648 2513 11676
rect 1820 11636 1826 11648
rect 2501 11645 2513 11648
rect 2547 11645 2559 11679
rect 2746 11676 2774 11716
rect 4430 11704 4436 11756
rect 4488 11744 4494 11756
rect 4488 11716 4936 11744
rect 4488 11704 4494 11716
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 2746 11648 3341 11676
rect 2501 11639 2559 11645
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 3329 11639 3387 11645
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 3970 11676 3976 11688
rect 3467 11648 3976 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 1296 11611 1354 11617
rect 1296 11577 1308 11611
rect 1342 11608 1354 11611
rect 1394 11608 1400 11620
rect 1342 11580 1400 11608
rect 1342 11577 1354 11580
rect 1296 11571 1354 11577
rect 1394 11568 1400 11580
rect 1452 11568 1458 11620
rect 3344 11552 3372 11639
rect 3970 11636 3976 11648
rect 4028 11676 4034 11688
rect 4540 11685 4568 11716
rect 4065 11679 4123 11685
rect 4065 11676 4077 11679
rect 4028 11648 4077 11676
rect 4028 11636 4034 11648
rect 4065 11645 4077 11648
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11645 4583 11679
rect 4525 11639 4583 11645
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11676 4675 11679
rect 4798 11676 4804 11688
rect 4663 11648 4804 11676
rect 4663 11645 4675 11648
rect 4617 11639 4675 11645
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4433 11611 4491 11617
rect 4433 11608 4445 11611
rect 4203 11580 4445 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 4433 11577 4445 11580
rect 4479 11608 4491 11611
rect 4632 11608 4660 11639
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 4908 11685 4936 11716
rect 5718 11704 5724 11756
rect 5776 11704 5782 11756
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 5074 11636 5080 11688
rect 5132 11676 5138 11688
rect 5169 11679 5227 11685
rect 5169 11676 5181 11679
rect 5132 11648 5181 11676
rect 5132 11636 5138 11648
rect 5169 11645 5181 11648
rect 5215 11645 5227 11679
rect 5169 11639 5227 11645
rect 5261 11679 5319 11685
rect 5261 11645 5273 11679
rect 5307 11676 5319 11679
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 5307 11648 5641 11676
rect 5307 11645 5319 11648
rect 5261 11639 5319 11645
rect 5629 11645 5641 11648
rect 5675 11645 5687 11679
rect 5736 11676 5764 11704
rect 6012 11685 6040 11784
rect 11333 11781 11345 11815
rect 11379 11812 11391 11815
rect 11379 11784 11928 11812
rect 11379 11781 11391 11784
rect 11333 11775 11391 11781
rect 8588 11716 9260 11744
rect 5905 11679 5963 11685
rect 5905 11676 5917 11679
rect 5736 11648 5917 11676
rect 5629 11639 5687 11645
rect 5905 11645 5917 11648
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 5997 11679 6055 11685
rect 5997 11645 6009 11679
rect 6043 11645 6055 11679
rect 5997 11639 6055 11645
rect 4479 11580 4660 11608
rect 4479 11577 4491 11580
rect 4433 11571 4491 11577
rect 4706 11568 4712 11620
rect 4764 11568 4770 11620
rect 4982 11568 4988 11620
rect 5040 11608 5046 11620
rect 5537 11611 5595 11617
rect 5537 11608 5549 11611
rect 5040 11580 5549 11608
rect 5040 11568 5046 11580
rect 5537 11577 5549 11580
rect 5583 11577 5595 11611
rect 5644 11608 5672 11639
rect 7558 11636 7564 11688
rect 7616 11676 7622 11688
rect 8588 11685 8616 11716
rect 9232 11688 9260 11716
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 11900 11753 11928 11784
rect 11885 11747 11943 11753
rect 10100 11716 11284 11744
rect 10100 11704 10106 11716
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 7616 11648 8401 11676
rect 7616 11636 7622 11648
rect 8389 11645 8401 11648
rect 8435 11645 8447 11679
rect 8389 11639 8447 11645
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 8662 11636 8668 11688
rect 8720 11636 8726 11688
rect 8754 11636 8760 11688
rect 8812 11636 8818 11688
rect 9214 11636 9220 11688
rect 9272 11676 9278 11688
rect 9272 11648 9444 11676
rect 9272 11636 9278 11648
rect 8772 11608 8800 11636
rect 9416 11608 9444 11648
rect 9582 11636 9588 11688
rect 9640 11685 9646 11688
rect 9640 11679 9663 11685
rect 9651 11645 9663 11679
rect 9640 11639 9663 11645
rect 9640 11636 9646 11639
rect 9858 11636 9864 11688
rect 9916 11636 9922 11688
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11670 10011 11679
rect 10410 11676 10416 11688
rect 10060 11670 10416 11676
rect 9999 11648 10416 11670
rect 9999 11645 10088 11648
rect 9953 11642 10088 11645
rect 9953 11639 10011 11642
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 10502 11636 10508 11688
rect 10560 11676 10566 11688
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 10560 11648 11069 11676
rect 10560 11636 10566 11648
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 11149 11679 11207 11685
rect 11149 11645 11161 11679
rect 11195 11645 11207 11679
rect 11149 11639 11207 11645
rect 9490 11608 9496 11620
rect 5644 11580 6132 11608
rect 8772 11580 9332 11608
rect 9416 11580 9496 11608
rect 5537 11571 5595 11577
rect 6104 11552 6132 11580
rect 9304 11552 9332 11580
rect 9490 11568 9496 11580
rect 9548 11608 9554 11620
rect 9769 11611 9827 11617
rect 9769 11608 9781 11611
rect 9548 11580 9781 11608
rect 9548 11568 9554 11580
rect 9769 11577 9781 11580
rect 9815 11577 9827 11611
rect 9769 11571 9827 11577
rect 10870 11568 10876 11620
rect 10928 11568 10934 11620
rect 1210 11500 1216 11552
rect 1268 11500 1274 11552
rect 3326 11500 3332 11552
rect 3384 11500 3390 11552
rect 5810 11500 5816 11552
rect 5868 11500 5874 11552
rect 6086 11500 6092 11552
rect 6144 11500 6150 11552
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 8941 11543 8999 11549
rect 8941 11540 8953 11543
rect 8076 11512 8953 11540
rect 8076 11500 8082 11512
rect 8941 11509 8953 11512
rect 8987 11509 8999 11543
rect 9304 11512 9312 11552
rect 8941 11503 8999 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 10137 11543 10195 11549
rect 10137 11540 10149 11543
rect 9456 11512 10149 11540
rect 9456 11500 9462 11512
rect 10137 11509 10149 11512
rect 10183 11509 10195 11543
rect 11164 11540 11192 11639
rect 11256 11608 11284 11716
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11744 12403 11747
rect 12544 11744 12572 11840
rect 14829 11815 14887 11821
rect 14829 11812 14841 11815
rect 14108 11784 14841 11812
rect 14108 11756 14136 11784
rect 14829 11781 14841 11784
rect 14875 11781 14887 11815
rect 17129 11815 17187 11821
rect 17129 11812 17141 11815
rect 14829 11775 14887 11781
rect 15488 11784 17141 11812
rect 13630 11744 13636 11756
rect 12391 11716 12572 11744
rect 12912 11716 13636 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 11606 11636 11612 11688
rect 11664 11676 11670 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11664 11648 12081 11676
rect 11664 11636 11670 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11676 12495 11679
rect 12526 11676 12532 11688
rect 12483 11648 12532 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 12526 11636 12532 11648
rect 12584 11636 12590 11688
rect 12912 11685 12940 11716
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 14090 11744 14096 11756
rect 14016 11716 14096 11744
rect 14016 11685 14044 11716
rect 14090 11704 14096 11716
rect 14148 11704 14154 11756
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 14844 11716 15393 11744
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 13541 11679 13599 11685
rect 13541 11645 13553 11679
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11645 14059 11679
rect 14001 11639 14059 11645
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11645 14243 11679
rect 14185 11639 14243 11645
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11676 14335 11679
rect 14458 11676 14464 11688
rect 14323 11648 14464 11676
rect 14323 11645 14335 11648
rect 14277 11639 14335 11645
rect 12802 11608 12808 11620
rect 11256 11580 12808 11608
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 13556 11608 13584 11639
rect 13814 11608 13820 11620
rect 13556 11580 13820 11608
rect 13814 11568 13820 11580
rect 13872 11608 13878 11620
rect 14200 11608 14228 11639
rect 14458 11636 14464 11648
rect 14516 11676 14522 11688
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 14516 11648 14657 11676
rect 14516 11636 14522 11648
rect 14645 11645 14657 11648
rect 14691 11676 14703 11679
rect 14844 11676 14872 11716
rect 15381 11713 15393 11716
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15488 11688 15516 11784
rect 17129 11781 17141 11784
rect 17175 11781 17187 11815
rect 17129 11775 17187 11781
rect 15654 11704 15660 11756
rect 15712 11704 15718 11756
rect 15746 11704 15752 11756
rect 15804 11744 15810 11756
rect 15804 11716 16068 11744
rect 15804 11704 15810 11716
rect 14691 11648 14872 11676
rect 14921 11679 14979 11685
rect 14691 11645 14703 11648
rect 14645 11639 14703 11645
rect 14921 11645 14933 11679
rect 14967 11676 14979 11679
rect 15197 11679 15255 11685
rect 15197 11676 15209 11679
rect 14967 11648 15209 11676
rect 14967 11645 14979 11648
rect 14921 11639 14979 11645
rect 15197 11645 15209 11648
rect 15243 11676 15255 11679
rect 15243 11648 15297 11676
rect 15243 11645 15255 11648
rect 15197 11639 15255 11645
rect 15212 11608 15240 11639
rect 15470 11636 15476 11688
rect 15528 11636 15534 11688
rect 15565 11679 15623 11685
rect 15565 11645 15577 11679
rect 15611 11676 15623 11679
rect 15672 11676 15700 11704
rect 16040 11685 16068 11716
rect 16960 11716 18644 11744
rect 15611 11648 15700 11676
rect 16025 11679 16083 11685
rect 15611 11645 15623 11648
rect 15565 11639 15623 11645
rect 16025 11645 16037 11679
rect 16071 11676 16083 11679
rect 16298 11676 16304 11688
rect 16071 11648 16304 11676
rect 16071 11645 16083 11648
rect 16025 11639 16083 11645
rect 16298 11636 16304 11648
rect 16356 11636 16362 11688
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 16960 11685 16988 11716
rect 17788 11685 17816 11716
rect 18616 11688 18644 11716
rect 16577 11679 16635 11685
rect 16577 11676 16589 11679
rect 16540 11648 16589 11676
rect 16540 11636 16546 11648
rect 16577 11645 16589 11648
rect 16623 11645 16635 11679
rect 16577 11639 16635 11645
rect 16945 11679 17003 11685
rect 16945 11645 16957 11679
rect 16991 11645 17003 11679
rect 16945 11639 17003 11645
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11676 17279 11679
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 17267 11648 17417 11676
rect 17267 11645 17279 11648
rect 17221 11639 17279 11645
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 17497 11679 17555 11685
rect 17497 11645 17509 11679
rect 17543 11676 17555 11679
rect 17773 11679 17831 11685
rect 17543 11648 17724 11676
rect 17543 11645 17555 11648
rect 17497 11639 17555 11645
rect 15657 11611 15715 11617
rect 15657 11608 15669 11611
rect 13872 11580 15148 11608
rect 15212 11580 15669 11608
rect 13872 11568 13878 11580
rect 13722 11540 13728 11552
rect 11164 11512 13728 11540
rect 10137 11503 10195 11509
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14918 11540 14924 11552
rect 14424 11512 14924 11540
rect 14424 11500 14430 11512
rect 14918 11500 14924 11512
rect 14976 11500 14982 11552
rect 15120 11549 15148 11580
rect 15657 11577 15669 11580
rect 15703 11608 15715 11611
rect 15933 11611 15991 11617
rect 15933 11608 15945 11611
rect 15703 11580 15945 11608
rect 15703 11577 15715 11580
rect 15657 11571 15715 11577
rect 15933 11577 15945 11580
rect 15979 11577 15991 11611
rect 16592 11608 16620 11639
rect 17236 11608 17264 11639
rect 16592 11580 17264 11608
rect 15933 11571 15991 11577
rect 17696 11552 17724 11648
rect 17773 11645 17785 11679
rect 17819 11645 17831 11679
rect 17773 11639 17831 11645
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11676 18291 11679
rect 18414 11676 18420 11688
rect 18279 11648 18420 11676
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 18509 11679 18567 11685
rect 18509 11645 18521 11679
rect 18555 11645 18567 11679
rect 18509 11639 18567 11645
rect 18524 11608 18552 11639
rect 18598 11636 18604 11688
rect 18656 11636 18662 11688
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 18156 11580 18552 11608
rect 18156 11552 18184 11580
rect 15105 11543 15163 11549
rect 15105 11509 15117 11543
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 16206 11500 16212 11552
rect 16264 11500 16270 11552
rect 17678 11500 17684 11552
rect 17736 11500 17742 11552
rect 18138 11500 18144 11552
rect 18196 11500 18202 11552
rect 18506 11500 18512 11552
rect 18564 11540 18570 11552
rect 18892 11540 18920 11639
rect 18564 11512 18920 11540
rect 18564 11500 18570 11512
rect 552 11450 19571 11472
rect 552 11398 5112 11450
rect 5164 11398 5176 11450
rect 5228 11398 5240 11450
rect 5292 11398 5304 11450
rect 5356 11398 5368 11450
rect 5420 11398 9827 11450
rect 9879 11398 9891 11450
rect 9943 11398 9955 11450
rect 10007 11398 10019 11450
rect 10071 11398 10083 11450
rect 10135 11398 14542 11450
rect 14594 11398 14606 11450
rect 14658 11398 14670 11450
rect 14722 11398 14734 11450
rect 14786 11398 14798 11450
rect 14850 11398 19257 11450
rect 19309 11398 19321 11450
rect 19373 11398 19385 11450
rect 19437 11398 19449 11450
rect 19501 11398 19513 11450
rect 19565 11398 19571 11450
rect 552 11376 19571 11398
rect 1302 11296 1308 11348
rect 1360 11296 1366 11348
rect 4801 11339 4859 11345
rect 4801 11305 4813 11339
rect 4847 11336 4859 11339
rect 4847 11308 7512 11336
rect 4847 11305 4859 11308
rect 4801 11299 4859 11305
rect 1394 11228 1400 11280
rect 1452 11228 1458 11280
rect 3234 11268 3240 11280
rect 1504 11240 3240 11268
rect 1412 11199 1440 11228
rect 1397 11193 1455 11199
rect 1397 11159 1409 11193
rect 1443 11159 1455 11193
rect 1397 11153 1455 11159
rect 1210 11092 1216 11144
rect 1268 11092 1274 11144
rect 1504 11141 1532 11240
rect 3234 11228 3240 11240
rect 3292 11268 3298 11280
rect 4338 11268 4344 11280
rect 3292 11240 4344 11268
rect 3292 11228 3298 11240
rect 1762 11209 1768 11212
rect 1756 11200 1768 11209
rect 1723 11172 1768 11200
rect 1756 11163 1768 11172
rect 1762 11160 1768 11163
rect 1820 11160 1826 11212
rect 3436 11209 3464 11240
rect 4338 11228 4344 11240
rect 4396 11268 4402 11280
rect 7484 11268 7512 11308
rect 7558 11296 7564 11348
rect 7616 11296 7622 11348
rect 9033 11339 9091 11345
rect 7760 11308 8248 11336
rect 7760 11268 7788 11308
rect 4396 11240 6224 11268
rect 7484 11240 7788 11268
rect 7920 11271 7978 11277
rect 4396 11228 4402 11240
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11169 3479 11203
rect 3421 11163 3479 11169
rect 3688 11203 3746 11209
rect 3688 11169 3700 11203
rect 3734 11200 3746 11203
rect 3970 11200 3976 11212
rect 3734 11172 3976 11200
rect 3734 11169 3746 11172
rect 3688 11163 3746 11169
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 4893 11203 4951 11209
rect 4893 11200 4905 11203
rect 4764 11172 4905 11200
rect 4764 11160 4770 11172
rect 4893 11169 4905 11172
rect 4939 11169 4951 11203
rect 4893 11163 4951 11169
rect 4982 11160 4988 11212
rect 5040 11200 5046 11212
rect 5169 11203 5227 11209
rect 5169 11200 5181 11203
rect 5040 11172 5181 11200
rect 5040 11160 5046 11172
rect 5169 11169 5181 11172
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 5261 11203 5319 11209
rect 5261 11169 5273 11203
rect 5307 11200 5319 11203
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 5307 11172 5641 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 5629 11169 5641 11172
rect 5675 11200 5687 11203
rect 5810 11200 5816 11212
rect 5675 11172 5816 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 5810 11160 5816 11172
rect 5868 11200 5874 11212
rect 6196 11209 6224 11240
rect 7920 11237 7932 11271
rect 7966 11268 7978 11271
rect 8110 11268 8116 11280
rect 7966 11240 8116 11268
rect 7966 11237 7978 11240
rect 7920 11231 7978 11237
rect 8110 11228 8116 11240
rect 8168 11228 8174 11280
rect 8220 11268 8248 11308
rect 9033 11305 9045 11339
rect 9079 11336 9091 11339
rect 9582 11336 9588 11348
rect 9079 11308 9588 11336
rect 9079 11305 9091 11308
rect 9033 11299 9091 11305
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 9953 11339 10011 11345
rect 9953 11305 9965 11339
rect 9999 11305 10011 11339
rect 9953 11299 10011 11305
rect 9968 11268 9996 11299
rect 10502 11296 10508 11348
rect 10560 11296 10566 11348
rect 14090 11296 14096 11348
rect 14148 11336 14154 11348
rect 14277 11339 14335 11345
rect 14277 11336 14289 11339
rect 14148 11308 14289 11336
rect 14148 11296 14154 11308
rect 14277 11305 14289 11308
rect 14323 11305 14335 11339
rect 14277 11299 14335 11305
rect 15194 11296 15200 11348
rect 15252 11336 15258 11348
rect 15252 11308 16252 11336
rect 15252 11296 15258 11308
rect 8220 11240 9904 11268
rect 9968 11240 11744 11268
rect 5905 11203 5963 11209
rect 5905 11200 5917 11203
rect 5868 11172 5917 11200
rect 5868 11160 5874 11172
rect 5905 11169 5917 11172
rect 5951 11169 5963 11203
rect 5905 11163 5963 11169
rect 6181 11203 6239 11209
rect 6181 11169 6193 11203
rect 6227 11169 6239 11203
rect 6437 11203 6495 11209
rect 6437 11200 6449 11203
rect 6181 11163 6239 11169
rect 6288 11172 6449 11200
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11101 1547 11135
rect 5920 11132 5948 11163
rect 6288 11132 6316 11172
rect 6437 11169 6449 11172
rect 6483 11169 6495 11203
rect 6437 11163 6495 11169
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 7742 11200 7748 11212
rect 7699 11172 7748 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 9490 11160 9496 11212
rect 9548 11160 9554 11212
rect 9766 11160 9772 11212
rect 9824 11160 9830 11212
rect 5920 11104 6316 11132
rect 1489 11095 1547 11101
rect 1228 11064 1256 11092
rect 1504 11064 1532 11095
rect 9674 11092 9680 11144
rect 9732 11092 9738 11144
rect 9876 11132 9904 11240
rect 10042 11160 10048 11212
rect 10100 11160 10106 11212
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11200 11483 11203
rect 11606 11200 11612 11212
rect 11471 11172 11612 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 10152 11132 10180 11163
rect 9876 11104 10180 11132
rect 1228 11036 1532 11064
rect 9324 11036 9628 11064
rect 2869 10999 2927 11005
rect 2869 10965 2881 10999
rect 2915 10996 2927 10999
rect 3142 10996 3148 11008
rect 2915 10968 3148 10996
rect 2915 10965 2927 10968
rect 2869 10959 2927 10965
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 4985 10999 5043 11005
rect 4985 10965 4997 10999
rect 5031 10996 5043 10999
rect 5442 10996 5448 11008
rect 5031 10968 5448 10996
rect 5031 10965 5043 10968
rect 4985 10959 5043 10965
rect 5442 10956 5448 10968
rect 5500 10996 5506 11008
rect 5537 10999 5595 11005
rect 5537 10996 5549 10999
rect 5500 10968 5549 10996
rect 5500 10956 5506 10968
rect 5537 10965 5549 10968
rect 5583 10965 5595 10999
rect 5537 10959 5595 10965
rect 5994 10956 6000 11008
rect 6052 10956 6058 11008
rect 6362 10956 6368 11008
rect 6420 10996 6426 11008
rect 9324 10996 9352 11036
rect 6420 10968 9352 10996
rect 6420 10956 6426 10968
rect 9398 10956 9404 11008
rect 9456 10996 9462 11008
rect 9493 10999 9551 11005
rect 9493 10996 9505 10999
rect 9456 10968 9505 10996
rect 9456 10956 9462 10968
rect 9493 10965 9505 10968
rect 9539 10965 9551 10999
rect 9600 10996 9628 11036
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 10336 11064 10364 11163
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 11716 11141 11744 11240
rect 14458 11228 14464 11280
rect 14516 11268 14522 11280
rect 15562 11268 15568 11280
rect 14516 11240 14688 11268
rect 14516 11228 14522 11240
rect 11790 11160 11796 11212
rect 11848 11160 11854 11212
rect 13814 11160 13820 11212
rect 13872 11209 13878 11212
rect 13872 11200 13884 11209
rect 14369 11203 14427 11209
rect 13872 11172 14320 11200
rect 13872 11163 13884 11172
rect 13872 11160 13878 11163
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11132 12495 11135
rect 13078 11132 13084 11144
rect 12483 11104 13084 11132
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 9916 11036 10364 11064
rect 11532 11064 11560 11095
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 14090 11092 14096 11144
rect 14148 11092 14154 11144
rect 12713 11067 12771 11073
rect 12713 11064 12725 11067
rect 11532 11036 12725 11064
rect 9916 11024 9922 11036
rect 12713 11033 12725 11036
rect 12759 11033 12771 11067
rect 14292 11064 14320 11172
rect 14369 11169 14381 11203
rect 14415 11200 14427 11203
rect 14550 11200 14556 11212
rect 14415 11172 14556 11200
rect 14415 11169 14427 11172
rect 14369 11163 14427 11169
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 14660 11209 14688 11240
rect 15120 11240 15568 11268
rect 15120 11209 15148 11240
rect 15562 11228 15568 11240
rect 15620 11268 15626 11280
rect 16224 11268 16252 11308
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 16356 11308 16497 11336
rect 16356 11296 16362 11308
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 16485 11299 16543 11305
rect 15620 11240 15700 11268
rect 16224 11240 16620 11268
rect 15620 11228 15626 11240
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 15105 11203 15163 11209
rect 15105 11169 15117 11203
rect 15151 11169 15163 11203
rect 15105 11163 15163 11169
rect 15381 11203 15439 11209
rect 15381 11169 15393 11203
rect 15427 11200 15439 11203
rect 15470 11200 15476 11212
rect 15427 11172 15476 11200
rect 15427 11169 15439 11172
rect 15381 11163 15439 11169
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 15672 11209 15700 11240
rect 15657 11203 15715 11209
rect 15657 11169 15669 11203
rect 15703 11200 15715 11203
rect 16206 11200 16212 11212
rect 15703 11172 16212 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 16592 11209 16620 11240
rect 16301 11203 16359 11209
rect 16301 11169 16313 11203
rect 16347 11169 16359 11203
rect 16301 11163 16359 11169
rect 16577 11203 16635 11209
rect 16577 11169 16589 11203
rect 16623 11200 16635 11203
rect 16669 11203 16727 11209
rect 16669 11200 16681 11203
rect 16623 11172 16681 11200
rect 16623 11169 16635 11172
rect 16577 11163 16635 11169
rect 16669 11169 16681 11172
rect 16715 11169 16727 11203
rect 16669 11163 16727 11169
rect 16761 11203 16819 11209
rect 16761 11169 16773 11203
rect 16807 11200 16819 11203
rect 17678 11200 17684 11212
rect 16807 11172 17684 11200
rect 16807 11169 16819 11172
rect 16761 11163 16819 11169
rect 15488 11132 15516 11160
rect 15565 11135 15623 11141
rect 15565 11132 15577 11135
rect 15488 11104 15577 11132
rect 15565 11101 15577 11104
rect 15611 11101 15623 11135
rect 16316 11132 16344 11163
rect 16776 11132 16804 11163
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 17954 11160 17960 11212
rect 18012 11160 18018 11212
rect 19058 11160 19064 11212
rect 19116 11160 19122 11212
rect 16316 11104 16804 11132
rect 15565 11095 15623 11101
rect 18598 11092 18604 11144
rect 18656 11092 18662 11144
rect 15013 11067 15071 11073
rect 15013 11064 15025 11067
rect 14292 11036 15025 11064
rect 12713 11027 12771 11033
rect 15013 11033 15025 11036
rect 15059 11033 15071 11067
rect 15013 11027 15071 11033
rect 12066 10996 12072 11008
rect 9600 10968 12072 10996
rect 9493 10959 9551 10965
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 14918 10996 14924 11008
rect 13412 10968 14924 10996
rect 13412 10956 13418 10968
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 15654 10996 15660 11008
rect 15344 10968 15660 10996
rect 15344 10956 15350 10968
rect 15654 10956 15660 10968
rect 15712 10956 15718 11008
rect 17865 10999 17923 11005
rect 17865 10965 17877 10999
rect 17911 10996 17923 10999
rect 18138 10996 18144 11008
rect 17911 10968 18144 10996
rect 17911 10965 17923 10968
rect 17865 10959 17923 10965
rect 18138 10956 18144 10968
rect 18196 10996 18202 11008
rect 18690 10996 18696 11008
rect 18196 10968 18696 10996
rect 18196 10956 18202 10968
rect 18690 10956 18696 10968
rect 18748 10956 18754 11008
rect 552 10906 19412 10928
rect 552 10854 2755 10906
rect 2807 10854 2819 10906
rect 2871 10854 2883 10906
rect 2935 10854 2947 10906
rect 2999 10854 3011 10906
rect 3063 10854 7470 10906
rect 7522 10854 7534 10906
rect 7586 10854 7598 10906
rect 7650 10854 7662 10906
rect 7714 10854 7726 10906
rect 7778 10854 12185 10906
rect 12237 10854 12249 10906
rect 12301 10854 12313 10906
rect 12365 10854 12377 10906
rect 12429 10854 12441 10906
rect 12493 10854 16900 10906
rect 16952 10854 16964 10906
rect 17016 10854 17028 10906
rect 17080 10854 17092 10906
rect 17144 10854 17156 10906
rect 17208 10854 19412 10906
rect 552 10832 19412 10854
rect 3510 10792 3516 10804
rect 2884 10764 3516 10792
rect 2406 10548 2412 10600
rect 2464 10548 2470 10600
rect 2498 10548 2504 10600
rect 2556 10548 2562 10600
rect 2884 10597 2912 10764
rect 3510 10752 3516 10764
rect 3568 10752 3574 10804
rect 6454 10752 6460 10804
rect 6512 10752 6518 10804
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 7248 10764 7389 10792
rect 7248 10752 7254 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 7377 10755 7435 10761
rect 9674 10752 9680 10804
rect 9732 10752 9738 10804
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10100 10764 10180 10792
rect 10100 10752 10106 10764
rect 4617 10727 4675 10733
rect 4617 10693 4629 10727
rect 4663 10724 4675 10727
rect 10152 10724 10180 10764
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11425 10795 11483 10801
rect 11425 10792 11437 10795
rect 11296 10764 11437 10792
rect 11296 10752 11302 10764
rect 11425 10761 11437 10764
rect 11471 10761 11483 10795
rect 11425 10755 11483 10761
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 11848 10764 11897 10792
rect 11848 10752 11854 10764
rect 11885 10761 11897 10764
rect 11931 10761 11943 10795
rect 11885 10755 11943 10761
rect 11977 10795 12035 10801
rect 11977 10761 11989 10795
rect 12023 10761 12035 10795
rect 11977 10755 12035 10761
rect 10502 10724 10508 10736
rect 4663 10696 10088 10724
rect 4663 10693 4675 10696
rect 4617 10687 4675 10693
rect 3234 10616 3240 10668
rect 3292 10616 3298 10668
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 6641 10659 6699 10665
rect 5040 10628 5488 10656
rect 5040 10616 5046 10628
rect 2869 10591 2927 10597
rect 2869 10557 2881 10591
rect 2915 10588 2927 10591
rect 3050 10588 3056 10600
rect 2915 10560 3056 10588
rect 2915 10557 2927 10560
rect 2869 10551 2927 10557
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 3142 10548 3148 10600
rect 3200 10548 3206 10600
rect 3326 10548 3332 10600
rect 3384 10588 3390 10600
rect 5460 10597 5488 10628
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 8018 10656 8024 10668
rect 6687 10628 8024 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 8110 10616 8116 10668
rect 8168 10616 8174 10668
rect 3493 10591 3551 10597
rect 3493 10588 3505 10591
rect 3384 10560 3505 10588
rect 3384 10548 3390 10560
rect 3493 10557 3505 10560
rect 3539 10557 3551 10591
rect 3493 10551 3551 10557
rect 5445 10591 5503 10597
rect 5445 10557 5457 10591
rect 5491 10557 5503 10591
rect 5445 10551 5503 10557
rect 5626 10548 5632 10600
rect 5684 10588 5690 10600
rect 5813 10591 5871 10597
rect 5813 10588 5825 10591
rect 5684 10560 5825 10588
rect 5684 10548 5690 10560
rect 5813 10557 5825 10560
rect 5859 10557 5871 10591
rect 5813 10551 5871 10557
rect 6362 10548 6368 10600
rect 6420 10588 6426 10600
rect 6733 10591 6791 10597
rect 6733 10588 6745 10591
rect 6420 10560 6745 10588
rect 6420 10548 6426 10560
rect 6733 10557 6745 10560
rect 6779 10557 6791 10591
rect 7285 10591 7343 10597
rect 7285 10588 7297 10591
rect 6733 10551 6791 10557
rect 6840 10560 7297 10588
rect 2424 10520 2452 10548
rect 2685 10523 2743 10529
rect 2685 10520 2697 10523
rect 2424 10492 2697 10520
rect 2685 10489 2697 10492
rect 2731 10489 2743 10523
rect 2685 10483 2743 10489
rect 2777 10523 2835 10529
rect 2777 10489 2789 10523
rect 2823 10520 2835 10523
rect 3160 10520 3188 10548
rect 6457 10523 6515 10529
rect 6457 10520 6469 10523
rect 2823 10492 3188 10520
rect 4540 10492 6469 10520
rect 2823 10489 2835 10492
rect 2777 10483 2835 10489
rect 3053 10455 3111 10461
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 4540 10452 4568 10492
rect 6457 10489 6469 10492
rect 6503 10489 6515 10523
rect 6457 10483 6515 10489
rect 3099 10424 4568 10452
rect 5537 10455 5595 10461
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 5537 10421 5549 10455
rect 5583 10452 5595 10455
rect 5626 10452 5632 10464
rect 5583 10424 5632 10452
rect 5583 10421 5595 10424
rect 5537 10415 5595 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5905 10455 5963 10461
rect 5905 10421 5917 10455
rect 5951 10452 5963 10455
rect 5994 10452 6000 10464
rect 5951 10424 6000 10452
rect 5951 10421 5963 10424
rect 5905 10415 5963 10421
rect 5994 10412 6000 10424
rect 6052 10452 6058 10464
rect 6840 10452 6868 10560
rect 7285 10557 7297 10560
rect 7331 10588 7343 10591
rect 8128 10588 8156 10616
rect 7331 10560 8156 10588
rect 7331 10557 7343 10560
rect 7285 10551 7343 10557
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 9858 10588 9864 10600
rect 9732 10560 9864 10588
rect 9732 10548 9738 10560
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 10060 10597 10088 10696
rect 10152 10696 10508 10724
rect 10152 10597 10180 10696
rect 10502 10684 10508 10696
rect 10560 10684 10566 10736
rect 10781 10727 10839 10733
rect 10781 10693 10793 10727
rect 10827 10724 10839 10727
rect 10827 10696 11744 10724
rect 10827 10693 10839 10696
rect 10781 10687 10839 10693
rect 10962 10656 10968 10668
rect 10520 10628 10968 10656
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 10137 10591 10195 10597
rect 10137 10557 10149 10591
rect 10183 10557 10195 10591
rect 10137 10551 10195 10557
rect 10229 10591 10287 10597
rect 10229 10557 10241 10591
rect 10275 10557 10287 10591
rect 10229 10551 10287 10557
rect 9766 10520 9772 10532
rect 6932 10492 9772 10520
rect 6932 10461 6960 10492
rect 9766 10480 9772 10492
rect 9824 10480 9830 10532
rect 6052 10424 6868 10452
rect 6917 10455 6975 10461
rect 6052 10412 6058 10424
rect 6917 10421 6929 10455
rect 6963 10421 6975 10455
rect 6917 10415 6975 10421
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 10244 10452 10272 10551
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 10520 10597 10548 10628
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 10413 10591 10471 10597
rect 10413 10588 10425 10591
rect 10376 10560 10425 10588
rect 10376 10548 10382 10560
rect 10413 10557 10425 10560
rect 10459 10557 10471 10591
rect 10413 10551 10471 10557
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10557 10563 10591
rect 10505 10551 10563 10557
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10588 10655 10591
rect 10778 10588 10784 10600
rect 10643 10560 10784 10588
rect 10643 10557 10655 10560
rect 10597 10551 10655 10557
rect 10428 10520 10456 10551
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 11422 10548 11428 10600
rect 11480 10548 11486 10600
rect 11716 10597 11744 10696
rect 11790 10616 11796 10668
rect 11848 10656 11854 10668
rect 11992 10656 12020 10755
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14274 10792 14280 10804
rect 13964 10764 14280 10792
rect 13964 10752 13970 10764
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 14550 10752 14556 10804
rect 14608 10752 14614 10804
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 18325 10795 18383 10801
rect 18325 10792 18337 10795
rect 18288 10764 18337 10792
rect 18288 10752 18294 10764
rect 18325 10761 18337 10764
rect 18371 10761 18383 10795
rect 18325 10755 18383 10761
rect 11848 10628 12020 10656
rect 11848 10616 11854 10628
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 12124 10628 12296 10656
rect 12124 10616 12130 10628
rect 11609 10591 11667 10597
rect 11609 10557 11621 10591
rect 11655 10557 11667 10591
rect 11609 10551 11667 10557
rect 11701 10591 11759 10597
rect 11701 10557 11713 10591
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 10962 10520 10968 10532
rect 10428 10492 10968 10520
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 7800 10424 10272 10452
rect 11149 10455 11207 10461
rect 7800 10412 7806 10424
rect 11149 10421 11161 10455
rect 11195 10452 11207 10455
rect 11238 10452 11244 10464
rect 11195 10424 11244 10452
rect 11195 10421 11207 10424
rect 11149 10415 11207 10421
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 11624 10452 11652 10551
rect 12158 10548 12164 10600
rect 12216 10548 12222 10600
rect 12268 10597 12296 10628
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10588 13875 10591
rect 14568 10588 14596 10752
rect 15286 10724 15292 10736
rect 15166 10696 15292 10724
rect 15166 10656 15194 10696
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 14660 10628 15194 10656
rect 18141 10659 18199 10665
rect 14660 10597 14688 10628
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 18187 10628 18920 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 13863 10560 14596 10588
rect 14645 10591 14703 10597
rect 13863 10557 13875 10560
rect 13817 10551 13875 10557
rect 14645 10557 14657 10591
rect 14691 10557 14703 10591
rect 14645 10551 14703 10557
rect 15102 10548 15108 10600
rect 15160 10588 15166 10600
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 15160 10560 15301 10588
rect 15160 10548 15166 10560
rect 15289 10557 15301 10560
rect 15335 10588 15347 10591
rect 18156 10588 18184 10619
rect 18892 10600 18920 10628
rect 15335 10560 18184 10588
rect 18233 10591 18291 10597
rect 15335 10557 15347 10560
rect 15289 10551 15347 10557
rect 18233 10557 18245 10591
rect 18279 10557 18291 10591
rect 18233 10551 18291 10557
rect 11974 10480 11980 10532
rect 12032 10480 12038 10532
rect 15562 10529 15568 10532
rect 15556 10520 15568 10529
rect 12084 10492 15194 10520
rect 15523 10492 15568 10520
rect 12084 10452 12112 10492
rect 11624 10424 12112 10452
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12618 10452 12624 10464
rect 12483 10424 12624 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 15166 10452 15194 10492
rect 15556 10483 15568 10492
rect 15562 10480 15568 10483
rect 15620 10480 15626 10532
rect 17678 10480 17684 10532
rect 17736 10520 17742 10532
rect 17874 10523 17932 10529
rect 17874 10520 17886 10523
rect 17736 10492 17886 10520
rect 17736 10480 17742 10492
rect 17874 10489 17886 10492
rect 17920 10489 17932 10523
rect 18248 10520 18276 10551
rect 18690 10548 18696 10600
rect 18748 10548 18754 10600
rect 18874 10548 18880 10600
rect 18932 10548 18938 10600
rect 18782 10520 18788 10532
rect 18248 10492 18788 10520
rect 17874 10483 17932 10489
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 16206 10452 16212 10464
rect 15166 10424 16212 10452
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16390 10412 16396 10464
rect 16448 10452 16454 10464
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 16448 10424 16681 10452
rect 16448 10412 16454 10424
rect 16669 10421 16681 10424
rect 16715 10421 16727 10455
rect 16669 10415 16727 10421
rect 16758 10412 16764 10464
rect 16816 10412 16822 10464
rect 552 10362 19571 10384
rect 552 10310 5112 10362
rect 5164 10310 5176 10362
rect 5228 10310 5240 10362
rect 5292 10310 5304 10362
rect 5356 10310 5368 10362
rect 5420 10310 9827 10362
rect 9879 10310 9891 10362
rect 9943 10310 9955 10362
rect 10007 10310 10019 10362
rect 10071 10310 10083 10362
rect 10135 10310 14542 10362
rect 14594 10310 14606 10362
rect 14658 10310 14670 10362
rect 14722 10310 14734 10362
rect 14786 10310 14798 10362
rect 14850 10310 19257 10362
rect 19309 10310 19321 10362
rect 19373 10310 19385 10362
rect 19437 10310 19449 10362
rect 19501 10310 19513 10362
rect 19565 10310 19571 10362
rect 552 10288 19571 10310
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 6457 10251 6515 10257
rect 6457 10248 6469 10251
rect 5684 10220 6469 10248
rect 5684 10208 5690 10220
rect 6457 10217 6469 10220
rect 6503 10217 6515 10251
rect 9309 10251 9367 10257
rect 6457 10211 6515 10217
rect 7024 10220 7236 10248
rect 1480 10183 1538 10189
rect 1480 10149 1492 10183
rect 1526 10180 1538 10183
rect 1578 10180 1584 10192
rect 1526 10152 1584 10180
rect 1526 10149 1538 10152
rect 1480 10143 1538 10149
rect 1578 10140 1584 10152
rect 1636 10140 1642 10192
rect 3418 10140 3424 10192
rect 3476 10180 3482 10192
rect 7024 10180 7052 10220
rect 3476 10152 7052 10180
rect 7208 10180 7236 10220
rect 9309 10217 9321 10251
rect 9355 10248 9367 10251
rect 10686 10248 10692 10260
rect 9355 10220 10692 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 12066 10248 12072 10260
rect 11112 10220 12072 10248
rect 11112 10208 11118 10220
rect 12066 10208 12072 10220
rect 12124 10248 12130 10260
rect 12253 10251 12311 10257
rect 12253 10248 12265 10251
rect 12124 10220 12265 10248
rect 12124 10208 12130 10220
rect 12253 10217 12265 10220
rect 12299 10217 12311 10251
rect 12253 10211 12311 10217
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 14148 10220 14780 10248
rect 14148 10208 14154 10220
rect 10953 10183 11011 10189
rect 10953 10180 10965 10183
rect 7208 10152 10965 10180
rect 3476 10140 3482 10152
rect 10953 10149 10965 10152
rect 10999 10149 11011 10183
rect 10953 10143 11011 10149
rect 1210 10072 1216 10124
rect 1268 10072 1274 10124
rect 5442 10072 5448 10124
rect 5500 10072 5506 10124
rect 5994 10072 6000 10124
rect 6052 10072 6058 10124
rect 6089 10115 6147 10121
rect 6089 10081 6101 10115
rect 6135 10081 6147 10115
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 6089 10075 6147 10081
rect 6196 10084 6561 10112
rect 5460 10044 5488 10072
rect 6104 10044 6132 10075
rect 6196 10056 6224 10084
rect 6549 10081 6561 10084
rect 6595 10081 6607 10115
rect 6549 10075 6607 10081
rect 6730 10072 6736 10124
rect 6788 10072 6794 10124
rect 6822 10072 6828 10124
rect 6880 10112 6886 10124
rect 6989 10115 7047 10121
rect 6989 10112 7001 10115
rect 6880 10084 7001 10112
rect 6880 10072 6886 10084
rect 6989 10081 7001 10084
rect 7035 10081 7047 10115
rect 6989 10075 7047 10081
rect 7558 10072 7564 10124
rect 7616 10112 7622 10124
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 7616 10084 9505 10112
rect 7616 10072 7622 10084
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10081 9827 10115
rect 9769 10075 9827 10081
rect 5460 10016 6132 10044
rect 6178 10004 6184 10056
rect 6236 10004 6242 10056
rect 7742 10004 7748 10056
rect 7800 10004 7806 10056
rect 9582 10004 9588 10056
rect 9640 10004 9646 10056
rect 9784 10044 9812 10075
rect 14458 10072 14464 10124
rect 14516 10121 14522 10124
rect 14752 10121 14780 10220
rect 18230 10140 18236 10192
rect 18288 10180 18294 10192
rect 18610 10183 18668 10189
rect 18610 10180 18622 10183
rect 18288 10152 18622 10180
rect 18288 10140 18294 10152
rect 18610 10149 18622 10152
rect 18656 10149 18668 10183
rect 18610 10143 18668 10149
rect 14516 10112 14528 10121
rect 14737 10115 14795 10121
rect 14516 10084 14561 10112
rect 14516 10075 14528 10084
rect 14737 10081 14749 10115
rect 14783 10112 14795 10115
rect 15102 10112 15108 10124
rect 14783 10084 15108 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 14516 10072 14522 10075
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15838 10072 15844 10124
rect 15896 10112 15902 10124
rect 16301 10115 16359 10121
rect 16301 10112 16313 10115
rect 15896 10084 16313 10112
rect 15896 10072 15902 10084
rect 16301 10081 16313 10084
rect 16347 10081 16359 10115
rect 16301 10075 16359 10081
rect 16666 10072 16672 10124
rect 16724 10072 16730 10124
rect 18874 10072 18880 10124
rect 18932 10072 18938 10124
rect 10594 10044 10600 10056
rect 9784 10016 10600 10044
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12032 10016 12434 10044
rect 12032 10004 12038 10016
rect 2593 9979 2651 9985
rect 2593 9945 2605 9979
rect 2639 9976 2651 9979
rect 2639 9948 6500 9976
rect 2639 9945 2651 9948
rect 2593 9939 2651 9945
rect 5537 9911 5595 9917
rect 5537 9877 5549 9911
rect 5583 9908 5595 9911
rect 5902 9908 5908 9920
rect 5583 9880 5908 9908
rect 5583 9877 5595 9880
rect 5537 9871 5595 9877
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 6178 9868 6184 9920
rect 6236 9868 6242 9920
rect 6472 9908 6500 9948
rect 7760 9908 7788 10004
rect 8113 9979 8171 9985
rect 8113 9945 8125 9979
rect 8159 9976 8171 9979
rect 11054 9976 11060 9988
rect 8159 9948 11060 9976
rect 8159 9945 8171 9948
rect 8113 9939 8171 9945
rect 11054 9936 11060 9948
rect 11112 9936 11118 9988
rect 12406 9976 12434 10016
rect 16390 10004 16396 10056
rect 16448 10004 16454 10056
rect 16574 10004 16580 10056
rect 16632 10004 16638 10056
rect 17221 10047 17279 10053
rect 17221 10013 17233 10047
rect 17267 10044 17279 10047
rect 17310 10044 17316 10056
rect 17267 10016 17316 10044
rect 17267 10013 17279 10016
rect 17221 10007 17279 10013
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 12406 9948 13860 9976
rect 6472 9880 7788 9908
rect 9769 9911 9827 9917
rect 9769 9877 9781 9911
rect 9815 9908 9827 9911
rect 10226 9908 10232 9920
rect 9815 9880 10232 9908
rect 9815 9877 9827 9880
rect 9769 9871 9827 9877
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 12158 9908 12164 9920
rect 12032 9880 12164 9908
rect 12032 9868 12038 9880
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 13357 9911 13415 9917
rect 13357 9908 13369 9911
rect 12584 9880 13369 9908
rect 12584 9868 12590 9880
rect 13357 9877 13369 9880
rect 13403 9877 13415 9911
rect 13832 9908 13860 9948
rect 15102 9908 15108 9920
rect 13832 9880 15108 9908
rect 13357 9871 13415 9877
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 17494 9868 17500 9920
rect 17552 9868 17558 9920
rect 552 9818 19412 9840
rect 552 9766 2755 9818
rect 2807 9766 2819 9818
rect 2871 9766 2883 9818
rect 2935 9766 2947 9818
rect 2999 9766 3011 9818
rect 3063 9766 7470 9818
rect 7522 9766 7534 9818
rect 7586 9766 7598 9818
rect 7650 9766 7662 9818
rect 7714 9766 7726 9818
rect 7778 9766 12185 9818
rect 12237 9766 12249 9818
rect 12301 9766 12313 9818
rect 12365 9766 12377 9818
rect 12429 9766 12441 9818
rect 12493 9766 16900 9818
rect 16952 9766 16964 9818
rect 17016 9766 17028 9818
rect 17080 9766 17092 9818
rect 17144 9766 17156 9818
rect 17208 9766 19412 9818
rect 552 9744 19412 9766
rect 2409 9707 2467 9713
rect 2409 9673 2421 9707
rect 2455 9704 2467 9707
rect 2498 9704 2504 9716
rect 2455 9676 2504 9704
rect 2455 9673 2467 9676
rect 2409 9667 2467 9673
rect 2498 9664 2504 9676
rect 2556 9664 2562 9716
rect 6822 9704 6828 9716
rect 6288 9676 6828 9704
rect 5994 9636 6000 9648
rect 5000 9608 6000 9636
rect 1026 9460 1032 9512
rect 1084 9460 1090 9512
rect 4614 9460 4620 9512
rect 4672 9460 4678 9512
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 4798 9500 4804 9512
rect 4755 9472 4804 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 4798 9460 4804 9472
rect 4856 9500 4862 9512
rect 5000 9509 5028 9608
rect 5994 9596 6000 9608
rect 6052 9636 6058 9648
rect 6288 9645 6316 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 9214 9664 9220 9716
rect 9272 9704 9278 9716
rect 11609 9707 11667 9713
rect 9272 9676 11376 9704
rect 9272 9664 9278 9676
rect 6273 9639 6331 9645
rect 6273 9636 6285 9639
rect 6052 9608 6285 9636
rect 6052 9596 6058 9608
rect 6273 9605 6285 9608
rect 6319 9636 6331 9639
rect 11348 9636 11376 9676
rect 11609 9673 11621 9707
rect 11655 9704 11667 9707
rect 11790 9704 11796 9716
rect 11655 9676 11796 9704
rect 11655 9673 11667 9676
rect 11609 9667 11667 9673
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 13722 9664 13728 9716
rect 13780 9704 13786 9716
rect 17770 9704 17776 9716
rect 13780 9676 17776 9704
rect 13780 9664 13786 9676
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 18785 9707 18843 9713
rect 18785 9673 18797 9707
rect 18831 9704 18843 9707
rect 18966 9704 18972 9716
rect 18831 9676 18972 9704
rect 18831 9673 18843 9676
rect 18785 9667 18843 9673
rect 18966 9664 18972 9676
rect 19024 9664 19030 9716
rect 13814 9636 13820 9648
rect 6319 9608 6353 9636
rect 11348 9608 13820 9636
rect 6319 9605 6331 9608
rect 6273 9599 6331 9605
rect 6546 9568 6552 9580
rect 5460 9540 6552 9568
rect 5460 9509 5488 9540
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 11348 9568 11376 9608
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 11256 9540 11376 9568
rect 12345 9571 12403 9577
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 4856 9472 4905 9500
rect 4856 9460 4862 9472
rect 4893 9469 4905 9472
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 4985 9503 5043 9509
rect 4985 9469 4997 9503
rect 5031 9469 5043 9503
rect 4985 9463 5043 9469
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 5445 9503 5503 9509
rect 5445 9469 5457 9503
rect 5491 9469 5503 9503
rect 5445 9463 5503 9469
rect 1118 9392 1124 9444
rect 1176 9432 1182 9444
rect 1274 9435 1332 9441
rect 1274 9432 1286 9435
rect 1176 9404 1286 9432
rect 1176 9392 1182 9404
rect 1274 9401 1286 9404
rect 1320 9401 1332 9435
rect 4632 9432 4660 9460
rect 5092 9432 5120 9463
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 5718 9500 5724 9512
rect 5592 9472 5724 9500
rect 5592 9460 5598 9472
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 5905 9503 5963 9509
rect 5905 9469 5917 9503
rect 5951 9500 5963 9503
rect 6178 9500 6184 9512
rect 5951 9472 6184 9500
rect 5951 9469 5963 9472
rect 5905 9463 5963 9469
rect 4632 9404 5120 9432
rect 1274 9395 1332 9401
rect 5258 9392 5264 9444
rect 5316 9392 5322 9444
rect 5353 9435 5411 9441
rect 5353 9401 5365 9435
rect 5399 9401 5411 9435
rect 5353 9395 5411 9401
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9364 4675 9367
rect 4890 9364 4896 9376
rect 4663 9336 4896 9364
rect 4663 9333 4675 9336
rect 4617 9327 4675 9333
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5368 9364 5396 9395
rect 5442 9364 5448 9376
rect 5368 9336 5448 9364
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5629 9367 5687 9373
rect 5629 9333 5641 9367
rect 5675 9364 5687 9367
rect 5718 9364 5724 9376
rect 5675 9336 5724 9364
rect 5675 9333 5687 9336
rect 5629 9327 5687 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 5828 9364 5856 9463
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 6730 9500 6736 9512
rect 6687 9472 6736 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 9033 9503 9091 9509
rect 9033 9500 9045 9503
rect 7708 9472 9045 9500
rect 7708 9460 7714 9472
rect 9033 9469 9045 9472
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9289 9503 9347 9509
rect 9289 9500 9301 9503
rect 9180 9472 9301 9500
rect 9180 9460 9186 9472
rect 9289 9469 9301 9472
rect 9335 9469 9347 9503
rect 9289 9463 9347 9469
rect 10410 9460 10416 9512
rect 10468 9500 10474 9512
rect 10686 9500 10692 9512
rect 10468 9472 10692 9500
rect 10468 9460 10474 9472
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 11054 9460 11060 9512
rect 11112 9460 11118 9512
rect 11256 9509 11284 9540
rect 12345 9537 12357 9571
rect 12391 9537 12403 9571
rect 12345 9531 12403 9537
rect 11241 9503 11299 9509
rect 11241 9469 11253 9503
rect 11287 9469 11299 9503
rect 11241 9463 11299 9469
rect 11330 9460 11336 9512
rect 11388 9460 11394 9512
rect 11422 9460 11428 9512
rect 11480 9460 11486 9512
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 12250 9500 12256 9512
rect 11664 9472 12256 9500
rect 11664 9460 11670 9472
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 6196 9432 6224 9460
rect 6886 9435 6944 9441
rect 6886 9432 6898 9435
rect 6196 9404 6898 9432
rect 6886 9401 6898 9404
rect 6932 9401 6944 9435
rect 6886 9395 6944 9401
rect 8036 9404 10548 9432
rect 6178 9364 6184 9376
rect 5828 9336 6184 9364
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 8036 9373 8064 9404
rect 8021 9367 8079 9373
rect 8021 9333 8033 9367
rect 8067 9333 8079 9367
rect 8021 9327 8079 9333
rect 10410 9324 10416 9376
rect 10468 9324 10474 9376
rect 10520 9364 10548 9404
rect 10778 9392 10784 9444
rect 10836 9432 10842 9444
rect 11440 9432 11468 9460
rect 10836 9404 11468 9432
rect 11532 9404 11744 9432
rect 10836 9392 10842 9404
rect 11532 9364 11560 9404
rect 10520 9336 11560 9364
rect 11716 9364 11744 9404
rect 11790 9392 11796 9444
rect 11848 9432 11854 9444
rect 11974 9432 11980 9444
rect 11848 9404 11980 9432
rect 11848 9392 11854 9404
rect 11974 9392 11980 9404
rect 12032 9392 12038 9444
rect 12360 9432 12388 9531
rect 12526 9528 12532 9580
rect 12584 9528 12590 9580
rect 15841 9571 15899 9577
rect 12820 9540 14780 9568
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9500 12679 9503
rect 12710 9500 12716 9512
rect 12667 9472 12716 9500
rect 12667 9469 12679 9472
rect 12621 9463 12679 9469
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 12820 9432 12848 9540
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 13740 9432 13768 9463
rect 13998 9460 14004 9512
rect 14056 9460 14062 9512
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9500 14151 9503
rect 14274 9500 14280 9512
rect 14139 9472 14280 9500
rect 14139 9469 14151 9472
rect 14093 9463 14151 9469
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 12360 9404 12848 9432
rect 12912 9404 13768 9432
rect 12912 9364 12940 9404
rect 13814 9392 13820 9444
rect 13872 9432 13878 9444
rect 13909 9435 13967 9441
rect 13909 9432 13921 9435
rect 13872 9404 13921 9432
rect 13872 9392 13878 9404
rect 13909 9401 13921 9404
rect 13955 9432 13967 9435
rect 14292 9432 14320 9460
rect 14752 9432 14780 9540
rect 15841 9537 15853 9571
rect 15887 9568 15899 9571
rect 16666 9568 16672 9580
rect 15887 9540 16672 9568
rect 15887 9537 15899 9540
rect 15841 9531 15899 9537
rect 16666 9528 16672 9540
rect 16724 9568 16730 9580
rect 17129 9571 17187 9577
rect 17129 9568 17141 9571
rect 16724 9540 17141 9568
rect 16724 9528 16730 9540
rect 17129 9537 17141 9540
rect 17175 9537 17187 9571
rect 18782 9568 18788 9580
rect 17129 9531 17187 9537
rect 18708 9540 18788 9568
rect 15166 9472 16804 9500
rect 15166 9432 15194 9472
rect 16776 9444 16804 9472
rect 17034 9460 17040 9512
rect 17092 9460 17098 9512
rect 18708 9509 18736 9540
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 17396 9503 17454 9509
rect 17396 9500 17408 9503
rect 17328 9472 17408 9500
rect 13955 9404 14044 9432
rect 14292 9404 14697 9432
rect 14752 9404 15194 9432
rect 13955 9401 13967 9404
rect 13909 9395 13967 9401
rect 14016 9376 14044 9404
rect 11716 9336 12940 9364
rect 13173 9367 13231 9373
rect 13173 9333 13185 9367
rect 13219 9364 13231 9367
rect 13630 9364 13636 9376
rect 13219 9336 13636 9364
rect 13219 9333 13231 9336
rect 13173 9327 13231 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 13998 9324 14004 9376
rect 14056 9324 14062 9376
rect 14274 9324 14280 9376
rect 14332 9324 14338 9376
rect 14458 9324 14464 9376
rect 14516 9324 14522 9376
rect 14669 9364 14697 9404
rect 15286 9392 15292 9444
rect 15344 9432 15350 9444
rect 15574 9435 15632 9441
rect 15574 9432 15586 9435
rect 15344 9404 15586 9432
rect 15344 9392 15350 9404
rect 15574 9401 15586 9404
rect 15620 9401 15632 9435
rect 15574 9395 15632 9401
rect 16758 9392 16764 9444
rect 16816 9392 16822 9444
rect 16945 9435 17003 9441
rect 16945 9401 16957 9435
rect 16991 9432 17003 9435
rect 17328 9432 17356 9472
rect 17396 9469 17408 9472
rect 17442 9500 17454 9503
rect 18693 9503 18751 9509
rect 18693 9500 18705 9503
rect 17442 9472 18705 9500
rect 17442 9469 17454 9472
rect 17396 9463 17454 9469
rect 18693 9469 18705 9472
rect 18739 9469 18751 9503
rect 18693 9463 18751 9469
rect 16991 9404 17356 9432
rect 16991 9401 17003 9404
rect 16945 9395 17003 9401
rect 15930 9364 15936 9376
rect 14669 9336 15936 9364
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 18230 9324 18236 9376
rect 18288 9364 18294 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 18288 9336 18521 9364
rect 18288 9324 18294 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 552 9274 19571 9296
rect 552 9222 5112 9274
rect 5164 9222 5176 9274
rect 5228 9222 5240 9274
rect 5292 9222 5304 9274
rect 5356 9222 5368 9274
rect 5420 9222 9827 9274
rect 9879 9222 9891 9274
rect 9943 9222 9955 9274
rect 10007 9222 10019 9274
rect 10071 9222 10083 9274
rect 10135 9222 14542 9274
rect 14594 9222 14606 9274
rect 14658 9222 14670 9274
rect 14722 9222 14734 9274
rect 14786 9222 14798 9274
rect 14850 9222 19257 9274
rect 19309 9222 19321 9274
rect 19373 9222 19385 9274
rect 19437 9222 19449 9274
rect 19501 9222 19513 9274
rect 19565 9222 19571 9274
rect 552 9200 19571 9222
rect 1397 9163 1455 9169
rect 1397 9129 1409 9163
rect 1443 9160 1455 9163
rect 1578 9160 1584 9172
rect 1443 9132 1584 9160
rect 1443 9129 1455 9132
rect 1397 9123 1455 9129
rect 1578 9120 1584 9132
rect 1636 9160 1642 9172
rect 1946 9160 1952 9172
rect 1636 9132 1952 9160
rect 1636 9120 1642 9132
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 3142 9120 3148 9172
rect 3200 9160 3206 9172
rect 3200 9132 4752 9160
rect 3200 9120 3206 9132
rect 4154 9092 4160 9104
rect 1596 9064 4160 9092
rect 1026 8984 1032 9036
rect 1084 8984 1090 9036
rect 1118 8984 1124 9036
rect 1176 9024 1182 9036
rect 1305 9027 1363 9033
rect 1305 9024 1317 9027
rect 1176 8996 1317 9024
rect 1176 8984 1182 8996
rect 1305 8993 1317 8996
rect 1351 8993 1363 9027
rect 1305 8987 1363 8993
rect 1044 8956 1072 8984
rect 1486 8956 1492 8968
rect 1044 8928 1492 8956
rect 1486 8916 1492 8928
rect 1544 8956 1550 8968
rect 1596 8965 1624 9064
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 3068 9033 3096 9064
rect 4154 9052 4160 9064
rect 4212 9052 4218 9104
rect 4724 9101 4752 9132
rect 4798 9120 4804 9172
rect 4856 9120 4862 9172
rect 5077 9163 5135 9169
rect 5077 9129 5089 9163
rect 5123 9160 5135 9163
rect 5534 9160 5540 9172
rect 5123 9132 5540 9160
rect 5123 9129 5135 9132
rect 5077 9123 5135 9129
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 5902 9120 5908 9172
rect 5960 9120 5966 9172
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 9030 9120 9036 9172
rect 9088 9160 9094 9172
rect 9088 9132 9536 9160
rect 9088 9120 9094 9132
rect 4709 9095 4767 9101
rect 4709 9061 4721 9095
rect 4755 9061 4767 9095
rect 4816 9092 4844 9120
rect 4816 9064 5580 9092
rect 4709 9055 4767 9061
rect 1837 9027 1895 9033
rect 1837 9024 1849 9027
rect 1728 8996 1849 9024
rect 1728 8984 1734 8996
rect 1837 8993 1849 8996
rect 1883 8993 1895 9027
rect 1837 8987 1895 8993
rect 3053 9027 3111 9033
rect 3053 8993 3065 9027
rect 3099 8993 3111 9027
rect 3309 9027 3367 9033
rect 3309 9024 3321 9027
rect 3053 8987 3111 8993
rect 3160 8996 3321 9024
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 1544 8928 1593 8956
rect 1544 8916 1550 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 3160 8956 3188 8996
rect 3309 8993 3321 8996
rect 3355 8993 3367 9027
rect 3309 8987 3367 8993
rect 4522 8984 4528 9036
rect 4580 8984 4586 9036
rect 4798 8984 4804 9036
rect 4856 8984 4862 9036
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 2648 8928 3188 8956
rect 2648 8916 2654 8928
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 4908 8956 4936 8987
rect 4764 8928 4936 8956
rect 4764 8916 4770 8928
rect 5184 8900 5212 9064
rect 5350 8984 5356 9036
rect 5408 8984 5414 9036
rect 5552 9033 5580 9064
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 8993 5595 9027
rect 5537 8987 5595 8993
rect 5626 8984 5632 9036
rect 5684 8984 5690 9036
rect 5920 9024 5948 9120
rect 7208 9092 7236 9120
rect 6564 9064 7236 9092
rect 7828 9095 7886 9101
rect 5997 9027 6055 9033
rect 5997 9024 6009 9027
rect 5920 8996 6009 9024
rect 5997 8993 6009 8996
rect 6043 9024 6055 9027
rect 6089 9027 6147 9033
rect 6089 9024 6101 9027
rect 6043 8996 6101 9024
rect 6043 8993 6055 8996
rect 5997 8987 6055 8993
rect 6089 8993 6101 8996
rect 6135 8993 6147 9027
rect 6089 8987 6147 8993
rect 6270 8984 6276 9036
rect 6328 9024 6334 9036
rect 6564 9033 6592 9064
rect 7828 9061 7840 9095
rect 7874 9092 7886 9095
rect 7926 9092 7932 9104
rect 7874 9064 7932 9092
rect 7874 9061 7886 9064
rect 7828 9055 7886 9061
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 9309 9095 9367 9101
rect 9309 9061 9321 9095
rect 9355 9061 9367 9095
rect 9309 9055 9367 9061
rect 6549 9027 6607 9033
rect 6549 9024 6561 9027
rect 6328 8996 6561 9024
rect 6328 8984 6334 8996
rect 6549 8993 6561 8996
rect 6595 8993 6607 9027
rect 6549 8987 6607 8993
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 7156 8996 7573 9024
rect 7156 8984 7162 8996
rect 7561 8993 7573 8996
rect 7607 9024 7619 9027
rect 7650 9024 7656 9036
rect 7607 8996 7656 9024
rect 7607 8993 7619 8996
rect 7561 8987 7619 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 8754 8984 8760 9036
rect 8812 9024 8818 9036
rect 9033 9027 9091 9033
rect 9033 9024 9045 9027
rect 8812 8996 9045 9024
rect 8812 8984 8818 8996
rect 9033 8993 9045 8996
rect 9079 8993 9091 9027
rect 9033 8987 9091 8993
rect 9214 8984 9220 9036
rect 9272 8984 9278 9036
rect 9324 8956 9352 9055
rect 9401 9027 9459 9033
rect 9401 8993 9413 9027
rect 9447 9022 9459 9027
rect 9508 9022 9536 9132
rect 9582 9120 9588 9172
rect 9640 9120 9646 9172
rect 11146 9120 11152 9172
rect 11204 9120 11210 9172
rect 11330 9120 11336 9172
rect 11388 9160 11394 9172
rect 11698 9160 11704 9172
rect 11388 9132 11704 9160
rect 11388 9120 11394 9132
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 12069 9163 12127 9169
rect 12069 9129 12081 9163
rect 12115 9160 12127 9163
rect 12526 9160 12532 9172
rect 12115 9132 12532 9160
rect 12115 9129 12127 9132
rect 12069 9123 12127 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 12618 9120 12624 9172
rect 12676 9160 12682 9172
rect 13265 9163 13323 9169
rect 12676 9132 12848 9160
rect 12676 9120 12682 9132
rect 11164 9092 11192 9120
rect 11241 9095 11299 9101
rect 11241 9092 11253 9095
rect 9447 8994 9536 9022
rect 9646 9064 11008 9092
rect 11164 9064 11253 9092
rect 9447 8993 9459 8994
rect 9401 8987 9459 8993
rect 9646 8956 9674 9064
rect 10229 9027 10287 9033
rect 10229 8993 10241 9027
rect 10275 9024 10287 9027
rect 10318 9024 10324 9036
rect 10275 8996 10324 9024
rect 10275 8993 10287 8996
rect 10229 8987 10287 8993
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10413 9027 10471 9033
rect 10413 8993 10425 9027
rect 10459 8993 10471 9027
rect 10413 8987 10471 8993
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 9024 10655 9027
rect 10686 9024 10692 9036
rect 10643 8996 10692 9024
rect 10643 8993 10655 8996
rect 10597 8987 10655 8993
rect 10428 8956 10456 8987
rect 8956 8928 9260 8956
rect 5166 8848 5172 8900
rect 5224 8848 5230 8900
rect 5261 8891 5319 8897
rect 5261 8857 5273 8891
rect 5307 8888 5319 8891
rect 5442 8888 5448 8900
rect 5307 8860 5448 8888
rect 5307 8857 5319 8860
rect 5261 8851 5319 8857
rect 5442 8848 5448 8860
rect 5500 8888 5506 8900
rect 8956 8897 8984 8928
rect 6181 8891 6239 8897
rect 6181 8888 6193 8891
rect 5500 8860 6193 8888
rect 5500 8848 5506 8860
rect 6181 8857 6193 8860
rect 6227 8857 6239 8891
rect 6181 8851 6239 8857
rect 8941 8891 8999 8897
rect 8941 8857 8953 8891
rect 8987 8857 8999 8891
rect 9232 8888 9260 8928
rect 9304 8928 9352 8956
rect 9416 8928 9674 8956
rect 10060 8928 10456 8956
rect 9304 8888 9332 8928
rect 9416 8900 9444 8928
rect 9232 8860 9332 8888
rect 8941 8851 8999 8857
rect 9398 8848 9404 8900
rect 9456 8848 9462 8900
rect 2958 8780 2964 8832
rect 3016 8780 3022 8832
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 5534 8820 5540 8832
rect 4479 8792 5540 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 5905 8823 5963 8829
rect 5905 8789 5917 8823
rect 5951 8820 5963 8823
rect 5994 8820 6000 8832
rect 5951 8792 6000 8820
rect 5951 8789 5963 8792
rect 5905 8783 5963 8789
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 6270 8780 6276 8832
rect 6328 8820 6334 8832
rect 6457 8823 6515 8829
rect 6457 8820 6469 8823
rect 6328 8792 6469 8820
rect 6328 8780 6334 8792
rect 6457 8789 6469 8792
rect 6503 8789 6515 8823
rect 6457 8783 6515 8789
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 9214 8820 9220 8832
rect 8904 8792 9220 8820
rect 8904 8780 8910 8792
rect 9214 8780 9220 8792
rect 9272 8820 9278 8832
rect 10060 8820 10088 8928
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 10520 8888 10548 8987
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 10980 9033 11008 9064
rect 11241 9061 11253 9064
rect 11287 9061 11299 9095
rect 11422 9092 11428 9104
rect 11241 9055 11299 9061
rect 11348 9064 11428 9092
rect 10965 9027 11023 9033
rect 10965 8993 10977 9027
rect 11011 8993 11023 9027
rect 10965 8987 11023 8993
rect 11146 8984 11152 9036
rect 11204 8984 11210 9036
rect 11348 9033 11376 9064
rect 11422 9052 11428 9064
rect 11480 9092 11486 9104
rect 12434 9092 12440 9104
rect 11480 9064 12020 9092
rect 11480 9052 11486 9064
rect 11992 9036 12020 9064
rect 12268 9064 12440 9092
rect 11333 9027 11391 9033
rect 11333 8993 11345 9027
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 11514 8984 11520 9036
rect 11572 8984 11578 9036
rect 11606 8984 11612 9036
rect 11664 8984 11670 9036
rect 11882 8984 11888 9036
rect 11940 8984 11946 9036
rect 11974 8984 11980 9036
rect 12032 8984 12038 9036
rect 12268 9033 12296 9064
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 8993 12311 9027
rect 12253 8987 12311 8993
rect 12342 8984 12348 9036
rect 12400 8984 12406 9036
rect 12710 8984 12716 9036
rect 12768 8984 12774 9036
rect 12820 9024 12848 9132
rect 13265 9129 13277 9163
rect 13311 9160 13323 9163
rect 14090 9160 14096 9172
rect 13311 9132 14096 9160
rect 13311 9129 13323 9132
rect 13265 9123 13323 9129
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 14274 9120 14280 9172
rect 14332 9120 14338 9172
rect 14458 9120 14464 9172
rect 14516 9120 14522 9172
rect 14645 9163 14703 9169
rect 14645 9129 14657 9163
rect 14691 9160 14703 9163
rect 14691 9132 15516 9160
rect 14691 9129 14703 9132
rect 14645 9123 14703 9129
rect 13538 9052 13544 9104
rect 13596 9092 13602 9104
rect 13725 9095 13783 9101
rect 13725 9092 13737 9095
rect 13596 9064 13737 9092
rect 13596 9052 13602 9064
rect 13725 9061 13737 9064
rect 13771 9061 13783 9095
rect 13725 9055 13783 9061
rect 12897 9027 12955 9033
rect 12897 9024 12909 9027
rect 12820 8996 12909 9024
rect 12897 8993 12909 8996
rect 12943 8993 12955 9027
rect 12897 8987 12955 8993
rect 13262 8984 13268 9036
rect 13320 9024 13326 9036
rect 13449 9027 13507 9033
rect 13449 9024 13461 9027
rect 13320 8996 13461 9024
rect 13320 8984 13326 8996
rect 13449 8993 13461 8996
rect 13495 8993 13507 9027
rect 13449 8987 13507 8993
rect 13633 9027 13691 9033
rect 13633 8993 13645 9027
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 11532 8956 11560 8984
rect 11112 8928 11560 8956
rect 11793 8959 11851 8965
rect 11112 8916 11118 8928
rect 11793 8925 11805 8959
rect 11839 8925 11851 8959
rect 12360 8956 12388 8984
rect 13648 8956 13676 8987
rect 13814 8984 13820 9036
rect 13872 8984 13878 9036
rect 14090 8984 14096 9036
rect 14148 9024 14154 9036
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 14148 8996 14197 9024
rect 14148 8984 14154 8996
rect 14185 8993 14197 8996
rect 14231 8993 14243 9027
rect 14292 9024 14320 9120
rect 14476 9092 14504 9120
rect 15194 9092 15200 9104
rect 14476 9064 14780 9092
rect 14752 9033 14780 9064
rect 14844 9064 15200 9092
rect 14369 9027 14427 9033
rect 14369 9024 14381 9027
rect 14292 8996 14381 9024
rect 14185 8987 14243 8993
rect 14369 8993 14381 8996
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 14461 9027 14519 9033
rect 14461 8993 14473 9027
rect 14507 8993 14519 9027
rect 14461 8987 14519 8993
rect 14737 9027 14795 9033
rect 14737 8993 14749 9027
rect 14783 8993 14795 9027
rect 14737 8987 14795 8993
rect 13722 8956 13728 8968
rect 12360 8928 13299 8956
rect 13648 8928 13728 8956
rect 11793 8919 11851 8925
rect 10468 8860 10548 8888
rect 10781 8891 10839 8897
rect 10468 8848 10474 8860
rect 10781 8857 10793 8891
rect 10827 8888 10839 8891
rect 11808 8888 11836 8919
rect 13170 8888 13176 8900
rect 10827 8860 11744 8888
rect 11808 8860 13176 8888
rect 10827 8857 10839 8860
rect 10781 8851 10839 8857
rect 9272 8792 10088 8820
rect 11517 8823 11575 8829
rect 9272 8780 9278 8792
rect 11517 8789 11529 8823
rect 11563 8820 11575 8823
rect 11609 8823 11667 8829
rect 11609 8820 11621 8823
rect 11563 8792 11621 8820
rect 11563 8789 11575 8792
rect 11517 8783 11575 8789
rect 11609 8789 11621 8792
rect 11655 8789 11667 8823
rect 11716 8820 11744 8860
rect 13170 8848 13176 8860
rect 13228 8848 13234 8900
rect 13271 8888 13299 8928
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 14274 8956 14280 8968
rect 14056 8928 14280 8956
rect 14056 8916 14062 8928
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 14476 8956 14504 8987
rect 14844 8956 14872 9064
rect 15194 9052 15200 9064
rect 15252 9052 15258 9104
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 8993 14979 9027
rect 14921 8987 14979 8993
rect 14476 8928 14872 8956
rect 14936 8956 14964 8987
rect 15286 8984 15292 9036
rect 15344 8984 15350 9036
rect 15488 9033 15516 9132
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 18141 9163 18199 9169
rect 18141 9160 18153 9163
rect 16264 9132 18153 9160
rect 16264 9120 16270 9132
rect 18141 9129 18153 9132
rect 18187 9129 18199 9163
rect 18141 9123 18199 9129
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 18877 9163 18935 9169
rect 18877 9160 18889 9163
rect 18564 9132 18889 9160
rect 18564 9120 18570 9132
rect 18877 9129 18889 9132
rect 18923 9129 18935 9163
rect 18877 9123 18935 9129
rect 16936 9095 16994 9101
rect 16936 9061 16948 9095
rect 16982 9092 16994 9095
rect 17034 9092 17040 9104
rect 16982 9064 17040 9092
rect 16982 9061 16994 9064
rect 16936 9055 16994 9061
rect 17034 9052 17040 9064
rect 17092 9092 17098 9104
rect 17310 9092 17316 9104
rect 17092 9064 17316 9092
rect 17092 9052 17098 9064
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 15473 9027 15531 9033
rect 15473 8993 15485 9027
rect 15519 8993 15531 9027
rect 15473 8987 15531 8993
rect 16666 8984 16672 9036
rect 16724 8984 16730 9036
rect 17862 8984 17868 9036
rect 17920 9024 17926 9036
rect 18325 9027 18383 9033
rect 18325 9024 18337 9027
rect 17920 8996 18337 9024
rect 17920 8984 17926 8996
rect 18325 8993 18337 8996
rect 18371 8993 18383 9027
rect 18325 8987 18383 8993
rect 18414 8984 18420 9036
rect 18472 8984 18478 9036
rect 18506 8984 18512 9036
rect 18564 8984 18570 9036
rect 18693 9027 18751 9033
rect 18693 8993 18705 9027
rect 18739 8993 18751 9027
rect 18693 8987 18751 8993
rect 18785 9027 18843 9033
rect 18785 8993 18797 9027
rect 18831 8993 18843 9027
rect 18785 8987 18843 8993
rect 15838 8956 15844 8968
rect 14936 8928 15844 8956
rect 14936 8888 14964 8928
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 15930 8916 15936 8968
rect 15988 8916 15994 8968
rect 18708 8956 18736 8987
rect 18064 8928 18736 8956
rect 18064 8897 18092 8928
rect 13271 8860 14964 8888
rect 18049 8891 18107 8897
rect 18049 8857 18061 8891
rect 18095 8857 18107 8891
rect 18800 8888 18828 8987
rect 18049 8851 18107 8857
rect 18708 8860 18828 8888
rect 18708 8832 18736 8860
rect 12618 8820 12624 8832
rect 11716 8792 12624 8820
rect 11609 8783 11667 8789
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 14001 8823 14059 8829
rect 14001 8789 14013 8823
rect 14047 8820 14059 8823
rect 14185 8823 14243 8829
rect 14185 8820 14197 8823
rect 14047 8792 14197 8820
rect 14047 8789 14059 8792
rect 14001 8783 14059 8789
rect 14185 8789 14197 8792
rect 14231 8789 14243 8823
rect 14185 8783 14243 8789
rect 18690 8780 18696 8832
rect 18748 8780 18754 8832
rect 552 8730 19412 8752
rect 552 8678 2755 8730
rect 2807 8678 2819 8730
rect 2871 8678 2883 8730
rect 2935 8678 2947 8730
rect 2999 8678 3011 8730
rect 3063 8678 7470 8730
rect 7522 8678 7534 8730
rect 7586 8678 7598 8730
rect 7650 8678 7662 8730
rect 7714 8678 7726 8730
rect 7778 8678 12185 8730
rect 12237 8678 12249 8730
rect 12301 8678 12313 8730
rect 12365 8678 12377 8730
rect 12429 8678 12441 8730
rect 12493 8678 16900 8730
rect 16952 8678 16964 8730
rect 17016 8678 17028 8730
rect 17080 8678 17092 8730
rect 17144 8678 17156 8730
rect 17208 8678 19412 8730
rect 552 8656 19412 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 2317 8619 2375 8625
rect 2317 8616 2329 8619
rect 1452 8588 2329 8616
rect 1452 8576 1458 8588
rect 2317 8585 2329 8588
rect 2363 8585 2375 8619
rect 2317 8579 2375 8585
rect 4706 8576 4712 8628
rect 4764 8616 4770 8628
rect 5626 8616 5632 8628
rect 4764 8588 5632 8616
rect 4764 8576 4770 8588
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 8570 8576 8576 8628
rect 8628 8616 8634 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8628 8588 9045 8616
rect 8628 8576 8634 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 9398 8616 9404 8628
rect 9033 8579 9091 8585
rect 9140 8588 9404 8616
rect 6012 8548 6040 8576
rect 5460 8520 6040 8548
rect 7377 8551 7435 8557
rect 2590 8480 2596 8492
rect 2424 8452 2596 8480
rect 1026 8372 1032 8424
rect 1084 8412 1090 8424
rect 1397 8415 1455 8421
rect 1397 8412 1409 8415
rect 1084 8384 1409 8412
rect 1084 8372 1090 8384
rect 1397 8381 1409 8384
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 1670 8372 1676 8424
rect 1728 8372 1734 8424
rect 2424 8421 2452 8452
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8412 2007 8415
rect 2409 8415 2467 8421
rect 1995 8384 2084 8412
rect 1995 8381 2007 8384
rect 1949 8375 2007 8381
rect 1118 8304 1124 8356
rect 1176 8344 1182 8356
rect 1305 8347 1363 8353
rect 1305 8344 1317 8347
rect 1176 8316 1317 8344
rect 1176 8304 1182 8316
rect 1305 8313 1317 8316
rect 1351 8344 1363 8347
rect 1581 8347 1639 8353
rect 1581 8344 1593 8347
rect 1351 8316 1593 8344
rect 1351 8313 1363 8316
rect 1305 8307 1363 8313
rect 1581 8313 1593 8316
rect 1627 8313 1639 8347
rect 1581 8307 1639 8313
rect 2056 8288 2084 8384
rect 2409 8381 2421 8415
rect 2455 8381 2467 8415
rect 2409 8375 2467 8381
rect 4614 8372 4620 8424
rect 4672 8412 4678 8424
rect 4893 8415 4951 8421
rect 4672 8384 4844 8412
rect 4672 8372 4678 8384
rect 1210 8236 1216 8288
rect 1268 8276 1274 8288
rect 1857 8279 1915 8285
rect 1857 8276 1869 8279
rect 1268 8248 1869 8276
rect 1268 8236 1274 8248
rect 1857 8245 1869 8248
rect 1903 8245 1915 8279
rect 1857 8239 1915 8245
rect 2038 8236 2044 8288
rect 2096 8236 2102 8288
rect 4525 8279 4583 8285
rect 4525 8245 4537 8279
rect 4571 8276 4583 8279
rect 4706 8276 4712 8288
rect 4571 8248 4712 8276
rect 4571 8245 4583 8248
rect 4525 8239 4583 8245
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 4816 8285 4844 8384
rect 4893 8381 4905 8415
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 4908 8344 4936 8375
rect 5166 8372 5172 8424
rect 5224 8372 5230 8424
rect 5460 8421 5488 8520
rect 7377 8517 7389 8551
rect 7423 8548 7435 8551
rect 9140 8548 9168 8588
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 9582 8616 9588 8628
rect 9539 8588 9588 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 10965 8619 11023 8625
rect 10965 8585 10977 8619
rect 11011 8616 11023 8619
rect 11054 8616 11060 8628
rect 11011 8588 11060 8616
rect 11011 8585 11023 8588
rect 10965 8579 11023 8585
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11664 8588 11805 8616
rect 11664 8576 11670 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 11793 8579 11851 8585
rect 11974 8576 11980 8628
rect 12032 8616 12038 8628
rect 12759 8619 12817 8625
rect 12759 8616 12771 8619
rect 12032 8588 12771 8616
rect 12032 8576 12038 8588
rect 12759 8585 12771 8588
rect 12805 8585 12817 8619
rect 17494 8616 17500 8628
rect 12759 8579 12817 8585
rect 13576 8588 17500 8616
rect 7423 8520 9168 8548
rect 7423 8517 7435 8520
rect 7377 8511 7435 8517
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 9766 8548 9772 8560
rect 9364 8520 9772 8548
rect 9364 8508 9370 8520
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 11330 8548 11336 8560
rect 10796 8520 11336 8548
rect 10796 8480 10824 8520
rect 11330 8508 11336 8520
rect 11388 8508 11394 8560
rect 13576 8548 13604 8588
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 17681 8619 17739 8625
rect 17681 8585 17693 8619
rect 17727 8616 17739 8619
rect 17770 8616 17776 8628
rect 17727 8588 17776 8616
rect 17727 8585 17739 8588
rect 17681 8579 17739 8585
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 11540 8520 13604 8548
rect 8588 8452 10824 8480
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 5534 8372 5540 8424
rect 5592 8412 5598 8424
rect 5721 8415 5779 8421
rect 5721 8412 5733 8415
rect 5592 8384 5733 8412
rect 5592 8372 5598 8384
rect 5721 8381 5733 8384
rect 5767 8381 5779 8415
rect 5721 8375 5779 8381
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6270 8421 6276 8424
rect 5997 8415 6055 8421
rect 5997 8412 6009 8415
rect 5960 8384 6009 8412
rect 5960 8372 5966 8384
rect 5997 8381 6009 8384
rect 6043 8381 6055 8415
rect 6264 8412 6276 8421
rect 6231 8384 6276 8412
rect 5997 8375 6055 8381
rect 6264 8375 6276 8384
rect 6270 8372 6276 8375
rect 6328 8372 6334 8424
rect 7834 8372 7840 8424
rect 7892 8372 7898 8424
rect 8386 8372 8392 8424
rect 8444 8372 8450 8424
rect 7852 8344 7880 8372
rect 8588 8353 8616 8452
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11112 8452 11468 8480
rect 11112 8440 11118 8452
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8412 8815 8415
rect 8846 8412 8852 8424
rect 8803 8384 8852 8412
rect 8803 8381 8815 8384
rect 8757 8375 8815 8381
rect 8573 8347 8631 8353
rect 8573 8344 8585 8347
rect 4908 8316 5396 8344
rect 7852 8316 8585 8344
rect 5368 8285 5396 8316
rect 8573 8313 8585 8316
rect 8619 8313 8631 8347
rect 8573 8307 8631 8313
rect 8662 8304 8668 8356
rect 8720 8304 8726 8356
rect 4801 8279 4859 8285
rect 4801 8245 4813 8279
rect 4847 8276 4859 8279
rect 5077 8279 5135 8285
rect 5077 8276 5089 8279
rect 4847 8248 5089 8276
rect 4847 8245 4859 8248
rect 4801 8239 4859 8245
rect 5077 8245 5089 8248
rect 5123 8245 5135 8279
rect 5077 8239 5135 8245
rect 5353 8279 5411 8285
rect 5353 8245 5365 8279
rect 5399 8276 5411 8279
rect 5442 8276 5448 8288
rect 5399 8248 5448 8276
rect 5399 8245 5411 8248
rect 5353 8239 5411 8245
rect 5442 8236 5448 8248
rect 5500 8276 5506 8288
rect 5629 8279 5687 8285
rect 5629 8276 5641 8279
rect 5500 8248 5641 8276
rect 5500 8236 5506 8248
rect 5629 8245 5641 8248
rect 5675 8245 5687 8279
rect 5629 8239 5687 8245
rect 8478 8236 8484 8288
rect 8536 8276 8542 8288
rect 8772 8276 8800 8375
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 8956 8384 9045 8412
rect 8956 8285 8984 8384
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 9214 8372 9220 8424
rect 9272 8372 9278 8424
rect 9306 8372 9312 8424
rect 9364 8372 9370 8424
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8412 10011 8415
rect 9999 8384 11008 8412
rect 9999 8381 10011 8384
rect 9953 8375 10011 8381
rect 10045 8347 10103 8353
rect 10045 8313 10057 8347
rect 10091 8344 10103 8347
rect 10321 8347 10379 8353
rect 10091 8316 10272 8344
rect 10091 8313 10103 8316
rect 10045 8307 10103 8313
rect 8536 8248 8800 8276
rect 8941 8279 8999 8285
rect 8536 8236 8542 8248
rect 8941 8245 8953 8279
rect 8987 8245 8999 8279
rect 8941 8239 8999 8245
rect 10134 8236 10140 8288
rect 10192 8236 10198 8288
rect 10244 8276 10272 8316
rect 10321 8313 10333 8347
rect 10367 8344 10379 8347
rect 10686 8344 10692 8356
rect 10367 8316 10692 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 10980 8288 11008 8384
rect 11238 8372 11244 8424
rect 11296 8372 11302 8424
rect 11440 8421 11468 8452
rect 11540 8421 11568 8520
rect 16022 8508 16028 8560
rect 16080 8508 16086 8560
rect 17310 8508 17316 8560
rect 17368 8548 17374 8560
rect 18417 8551 18475 8557
rect 18417 8548 18429 8551
rect 17368 8520 18429 8548
rect 17368 8508 17374 8520
rect 18417 8517 18429 8520
rect 18463 8517 18475 8551
rect 18417 8511 18475 8517
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 11900 8452 12081 8480
rect 11900 8424 11928 8452
rect 12069 8449 12081 8452
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12158 8440 12164 8492
rect 12216 8440 12222 8492
rect 13078 8480 13084 8492
rect 12268 8452 13084 8480
rect 12268 8424 12296 8452
rect 13078 8440 13084 8452
rect 13136 8480 13142 8492
rect 13136 8452 13400 8480
rect 13136 8440 13142 8452
rect 11425 8415 11483 8421
rect 11425 8381 11437 8415
rect 11471 8381 11483 8415
rect 11425 8375 11483 8381
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8381 11575 8415
rect 11517 8375 11575 8381
rect 11606 8372 11612 8424
rect 11664 8421 11670 8424
rect 11664 8415 11691 8421
rect 11679 8381 11691 8415
rect 11664 8375 11691 8381
rect 11664 8372 11670 8375
rect 11790 8372 11796 8424
rect 11848 8372 11854 8424
rect 11882 8372 11888 8424
rect 11940 8372 11946 8424
rect 11977 8415 12035 8421
rect 11977 8381 11989 8415
rect 12023 8381 12035 8415
rect 11977 8375 12035 8381
rect 11057 8347 11115 8353
rect 11057 8313 11069 8347
rect 11103 8344 11115 8347
rect 11808 8344 11836 8372
rect 11992 8344 12020 8375
rect 12250 8372 12256 8424
rect 12308 8372 12314 8424
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 13262 8412 13268 8424
rect 12584 8384 13268 8412
rect 12584 8372 12590 8384
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 11103 8316 11468 8344
rect 11808 8316 12020 8344
rect 12437 8347 12495 8353
rect 11103 8313 11115 8316
rect 11057 8307 11115 8313
rect 11440 8288 11468 8316
rect 12437 8313 12449 8347
rect 12483 8344 12495 8347
rect 13372 8344 13400 8452
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 16040 8480 16068 8508
rect 15528 8452 16436 8480
rect 15528 8440 15534 8452
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8412 13599 8415
rect 13630 8412 13636 8424
rect 13587 8384 13636 8412
rect 13587 8381 13599 8384
rect 13541 8375 13599 8381
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 13808 8415 13866 8421
rect 13808 8381 13820 8415
rect 13854 8412 13866 8415
rect 14182 8412 14188 8424
rect 13854 8384 14188 8412
rect 13854 8381 13866 8384
rect 13808 8375 13866 8381
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 15194 8412 15200 8424
rect 14976 8384 15200 8412
rect 14976 8372 14982 8384
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 16022 8372 16028 8424
rect 16080 8372 16086 8424
rect 16298 8372 16304 8424
rect 16356 8372 16362 8424
rect 16408 8421 16436 8452
rect 16666 8440 16672 8492
rect 16724 8480 16730 8492
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 16724 8452 17417 8480
rect 16724 8440 16730 8452
rect 17405 8449 17417 8452
rect 17451 8480 17463 8483
rect 17678 8480 17684 8492
rect 17451 8452 17684 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18138 8480 18144 8492
rect 18012 8452 18144 8480
rect 18012 8440 18018 8452
rect 18138 8440 18144 8452
rect 18196 8480 18202 8492
rect 18196 8452 18368 8480
rect 18196 8440 18202 8452
rect 16393 8415 16451 8421
rect 16393 8381 16405 8415
rect 16439 8381 16451 8415
rect 16393 8375 16451 8381
rect 17862 8372 17868 8424
rect 17920 8372 17926 8424
rect 18230 8372 18236 8424
rect 18288 8372 18294 8424
rect 18340 8421 18368 8452
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8381 18383 8415
rect 18432 8412 18460 8511
rect 18693 8415 18751 8421
rect 18693 8412 18705 8415
rect 18432 8384 18705 8412
rect 18325 8375 18383 8381
rect 18693 8381 18705 8384
rect 18739 8381 18751 8415
rect 18693 8375 18751 8381
rect 13998 8344 14004 8356
rect 12483 8316 13216 8344
rect 13372 8316 14004 8344
rect 12483 8313 12495 8316
rect 12437 8307 12495 8313
rect 10410 8276 10416 8288
rect 10244 8248 10416 8276
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 10962 8236 10968 8288
rect 11020 8236 11026 8288
rect 11422 8236 11428 8288
rect 11480 8236 11486 8288
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 12158 8276 12164 8288
rect 12032 8248 12164 8276
rect 12032 8236 12038 8248
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 13188 8276 13216 8316
rect 13998 8304 14004 8316
rect 14056 8304 14062 8356
rect 15562 8304 15568 8356
rect 15620 8344 15626 8356
rect 16209 8347 16267 8353
rect 16209 8344 16221 8347
rect 15620 8316 16221 8344
rect 15620 8304 15626 8316
rect 16209 8313 16221 8316
rect 16255 8313 16267 8347
rect 16209 8307 16267 8313
rect 16666 8304 16672 8356
rect 16724 8304 16730 8356
rect 17954 8304 17960 8356
rect 18012 8304 18018 8356
rect 18046 8304 18052 8356
rect 18104 8344 18110 8356
rect 18506 8344 18512 8356
rect 18104 8316 18512 8344
rect 18104 8304 18110 8316
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 13814 8276 13820 8288
rect 13188 8248 13820 8276
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 13906 8236 13912 8288
rect 13964 8276 13970 8288
rect 14458 8276 14464 8288
rect 13964 8248 14464 8276
rect 13964 8236 13970 8248
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 14918 8236 14924 8288
rect 14976 8236 14982 8288
rect 16390 8236 16396 8288
rect 16448 8276 16454 8288
rect 16577 8279 16635 8285
rect 16577 8276 16589 8279
rect 16448 8248 16589 8276
rect 16448 8236 16454 8248
rect 16577 8245 16589 8248
rect 16623 8245 16635 8279
rect 16577 8239 16635 8245
rect 18690 8236 18696 8288
rect 18748 8276 18754 8288
rect 18785 8279 18843 8285
rect 18785 8276 18797 8279
rect 18748 8248 18797 8276
rect 18748 8236 18754 8248
rect 18785 8245 18797 8248
rect 18831 8245 18843 8279
rect 18785 8239 18843 8245
rect 552 8186 19571 8208
rect 552 8134 5112 8186
rect 5164 8134 5176 8186
rect 5228 8134 5240 8186
rect 5292 8134 5304 8186
rect 5356 8134 5368 8186
rect 5420 8134 9827 8186
rect 9879 8134 9891 8186
rect 9943 8134 9955 8186
rect 10007 8134 10019 8186
rect 10071 8134 10083 8186
rect 10135 8134 14542 8186
rect 14594 8134 14606 8186
rect 14658 8134 14670 8186
rect 14722 8134 14734 8186
rect 14786 8134 14798 8186
rect 14850 8134 19257 8186
rect 19309 8134 19321 8186
rect 19373 8134 19385 8186
rect 19437 8134 19449 8186
rect 19501 8134 19513 8186
rect 19565 8134 19571 8186
rect 552 8112 19571 8134
rect 1210 8032 1216 8084
rect 1268 8032 1274 8084
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 1765 8075 1823 8081
rect 1765 8072 1777 8075
rect 1728 8044 1777 8072
rect 1728 8032 1734 8044
rect 1765 8041 1777 8044
rect 1811 8072 1823 8075
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 1811 8044 2329 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 3326 8072 3332 8084
rect 2317 8035 2375 8041
rect 2424 8044 3332 8072
rect 1029 7939 1087 7945
rect 1029 7905 1041 7939
rect 1075 7936 1087 7939
rect 1228 7936 1256 8032
rect 1688 8004 1716 8032
rect 1320 7976 1716 8004
rect 1320 7945 1348 7976
rect 1075 7908 1256 7936
rect 1305 7939 1363 7945
rect 1075 7905 1087 7908
rect 1029 7899 1087 7905
rect 1305 7905 1317 7939
rect 1351 7905 1363 7939
rect 1305 7899 1363 7905
rect 1394 7896 1400 7948
rect 1452 7896 1458 7948
rect 1489 7939 1547 7945
rect 1489 7905 1501 7939
rect 1535 7936 1547 7939
rect 1578 7936 1584 7948
rect 1535 7908 1584 7936
rect 1535 7905 1547 7908
rect 1489 7899 1547 7905
rect 1578 7896 1584 7908
rect 1636 7936 1642 7948
rect 2424 7945 2452 8044
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 4614 8032 4620 8084
rect 4672 8032 4678 8084
rect 5534 8072 5540 8084
rect 4908 8044 5540 8072
rect 4522 7964 4528 8016
rect 4580 7964 4586 8016
rect 1673 7939 1731 7945
rect 1673 7936 1685 7939
rect 1636 7908 1685 7936
rect 1636 7896 1642 7908
rect 1673 7905 1685 7908
rect 1719 7905 1731 7939
rect 2133 7939 2191 7945
rect 2133 7936 2145 7939
rect 1673 7899 1731 7905
rect 2056 7908 2145 7936
rect 934 7760 940 7812
rect 992 7800 998 7812
rect 1302 7800 1308 7812
rect 992 7772 1308 7800
rect 992 7760 998 7772
rect 1302 7760 1308 7772
rect 1360 7760 1366 7812
rect 1412 7732 1440 7896
rect 2056 7880 2084 7908
rect 2133 7905 2145 7908
rect 2179 7905 2191 7939
rect 2133 7899 2191 7905
rect 2409 7939 2467 7945
rect 2409 7905 2421 7939
rect 2455 7905 2467 7939
rect 2409 7899 2467 7905
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7905 2835 7939
rect 2777 7899 2835 7905
rect 2038 7828 2044 7880
rect 2096 7868 2102 7880
rect 2685 7871 2743 7877
rect 2685 7868 2697 7871
rect 2096 7840 2697 7868
rect 2096 7828 2102 7840
rect 2685 7837 2697 7840
rect 2731 7837 2743 7871
rect 2792 7868 2820 7899
rect 3142 7896 3148 7948
rect 3200 7896 3206 7948
rect 3973 7939 4031 7945
rect 3973 7905 3985 7939
rect 4019 7905 4031 7939
rect 3973 7899 4031 7905
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7936 4399 7939
rect 4540 7936 4568 7964
rect 4632 7945 4660 8032
rect 4908 7945 4936 8044
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 8849 8075 8907 8081
rect 5776 8044 8800 8072
rect 5776 8032 5782 8044
rect 7282 8013 7288 8016
rect 7276 8004 7288 8013
rect 7243 7976 7288 8004
rect 7276 7967 7288 7976
rect 7282 7964 7288 7967
rect 7340 7964 7346 8016
rect 8772 8004 8800 8044
rect 8849 8041 8861 8075
rect 8895 8072 8907 8075
rect 9030 8072 9036 8084
rect 8895 8044 9036 8072
rect 8895 8041 8907 8044
rect 8849 8035 8907 8041
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 9582 8072 9588 8084
rect 9456 8044 9588 8072
rect 9456 8032 9462 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10686 8072 10692 8084
rect 10100 8044 10692 8072
rect 10100 8032 10106 8044
rect 10686 8032 10692 8044
rect 10744 8072 10750 8084
rect 10744 8044 12112 8072
rect 10744 8032 10750 8044
rect 11054 8004 11060 8016
rect 8772 7976 11060 8004
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 11149 8007 11207 8013
rect 11149 7973 11161 8007
rect 11195 8004 11207 8007
rect 11330 8004 11336 8016
rect 11195 7976 11336 8004
rect 11195 7973 11207 7976
rect 11149 7967 11207 7973
rect 11330 7964 11336 7976
rect 11388 7964 11394 8016
rect 11532 7976 11836 8004
rect 4387 7908 4568 7936
rect 4617 7939 4675 7945
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 4617 7905 4629 7939
rect 4663 7905 4675 7939
rect 4617 7899 4675 7905
rect 4893 7939 4951 7945
rect 4893 7905 4905 7939
rect 4939 7905 4951 7939
rect 4893 7899 4951 7905
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7905 5227 7939
rect 5169 7899 5227 7905
rect 3234 7868 3240 7880
rect 2792 7840 3240 7868
rect 2685 7831 2743 7837
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 3988 7868 4016 7899
rect 4522 7868 4528 7880
rect 3988 7840 4528 7868
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 5184 7868 5212 7899
rect 5442 7896 5448 7948
rect 5500 7896 5506 7948
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7936 7067 7939
rect 7098 7936 7104 7948
rect 7055 7908 7104 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 8938 7896 8944 7948
rect 8996 7896 9002 7948
rect 9585 7939 9643 7945
rect 9585 7905 9597 7939
rect 9631 7936 9643 7939
rect 9631 7908 9996 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 4764 7840 5479 7868
rect 4764 7828 4770 7840
rect 2130 7760 2136 7812
rect 2188 7800 2194 7812
rect 3053 7803 3111 7809
rect 3053 7800 3065 7803
rect 2188 7772 3065 7800
rect 2188 7760 2194 7772
rect 3053 7769 3065 7772
rect 3099 7769 3111 7803
rect 3053 7763 3111 7769
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 4120 7772 4844 7800
rect 4120 7760 4126 7772
rect 2041 7735 2099 7741
rect 2041 7732 2053 7735
rect 1412 7704 2053 7732
rect 2041 7701 2053 7704
rect 2087 7701 2099 7735
rect 2041 7695 2099 7701
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 3927 7704 4261 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 4249 7701 4261 7704
rect 4295 7732 4307 7735
rect 4338 7732 4344 7744
rect 4295 7704 4344 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 4522 7692 4528 7744
rect 4580 7692 4586 7744
rect 4816 7741 4844 7772
rect 4890 7760 4896 7812
rect 4948 7800 4954 7812
rect 5353 7803 5411 7809
rect 5353 7800 5365 7803
rect 4948 7772 5365 7800
rect 4948 7760 4954 7772
rect 5353 7769 5365 7772
rect 5399 7769 5411 7803
rect 5451 7800 5479 7840
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 9600 7868 9628 7899
rect 9968 7880 9996 7908
rect 10042 7896 10048 7948
rect 10100 7896 10106 7948
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7905 10195 7939
rect 10137 7899 10195 7905
rect 10229 7939 10287 7945
rect 10229 7905 10241 7939
rect 10275 7936 10287 7939
rect 10410 7936 10416 7948
rect 10275 7908 10416 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 8904 7840 9628 7868
rect 9677 7871 9735 7877
rect 8904 7828 8910 7840
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 6270 7800 6276 7812
rect 5451 7772 6276 7800
rect 5353 7763 5411 7769
rect 6270 7760 6276 7772
rect 6328 7760 6334 7812
rect 9122 7760 9128 7812
rect 9180 7800 9186 7812
rect 9490 7800 9496 7812
rect 9180 7772 9496 7800
rect 9180 7760 9186 7772
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 9582 7760 9588 7812
rect 9640 7800 9646 7812
rect 9692 7800 9720 7831
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 10152 7868 10180 7899
rect 10410 7896 10416 7908
rect 10468 7896 10474 7948
rect 11532 7945 11560 7976
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7936 10563 7939
rect 11517 7939 11575 7945
rect 10551 7908 11468 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 10962 7868 10968 7880
rect 10152 7840 10968 7868
rect 10962 7828 10968 7840
rect 11020 7868 11026 7880
rect 11057 7871 11115 7877
rect 11057 7868 11069 7871
rect 11020 7840 11069 7868
rect 11020 7828 11026 7840
rect 11057 7837 11069 7840
rect 11103 7837 11115 7871
rect 11440 7868 11468 7908
rect 11517 7905 11529 7939
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 11609 7939 11667 7945
rect 11609 7905 11621 7939
rect 11655 7936 11667 7939
rect 11698 7936 11704 7948
rect 11655 7908 11704 7936
rect 11655 7905 11667 7908
rect 11609 7899 11667 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 11808 7936 11836 7976
rect 11882 7936 11888 7948
rect 11808 7908 11888 7936
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 12084 7945 12112 8044
rect 12342 8032 12348 8084
rect 12400 8032 12406 8084
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12676 8044 13032 8072
rect 12676 8032 12682 8044
rect 12158 7964 12164 8016
rect 12216 8004 12222 8016
rect 12216 7976 12388 8004
rect 12216 7964 12222 7976
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7936 12127 7939
rect 12360 7936 12388 7976
rect 12434 7964 12440 8016
rect 12492 8004 12498 8016
rect 12897 8007 12955 8013
rect 12897 8004 12909 8007
rect 12492 7976 12909 8004
rect 12492 7964 12498 7976
rect 12897 7973 12909 7976
rect 12943 7973 12955 8007
rect 13004 8004 13032 8044
rect 13078 8032 13084 8084
rect 13136 8072 13142 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13136 8044 13645 8072
rect 13136 8032 13142 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 14918 8032 14924 8084
rect 14976 8032 14982 8084
rect 15102 8032 15108 8084
rect 15160 8032 15166 8084
rect 15381 8075 15439 8081
rect 15381 8072 15393 8075
rect 15212 8044 15393 8072
rect 14936 8004 14964 8032
rect 15013 8007 15071 8013
rect 15013 8004 15025 8007
rect 13004 7976 13308 8004
rect 12897 7967 12955 7973
rect 12713 7939 12771 7945
rect 12713 7936 12725 7939
rect 12115 7908 12296 7936
rect 12360 7934 12434 7936
rect 12544 7934 12725 7936
rect 12360 7908 12725 7934
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 11790 7868 11796 7880
rect 11440 7840 11796 7868
rect 11057 7831 11115 7837
rect 11330 7800 11336 7812
rect 9640 7772 11336 7800
rect 9640 7760 9646 7772
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 11532 7744 11560 7840
rect 11790 7828 11796 7840
rect 11848 7868 11854 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11848 7840 12173 7868
rect 11848 7828 11854 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12268 7868 12296 7908
rect 12406 7906 12572 7908
rect 12713 7905 12725 7908
rect 12759 7905 12771 7939
rect 12713 7899 12771 7905
rect 12802 7896 12808 7948
rect 12860 7896 12866 7948
rect 13078 7896 13084 7948
rect 13136 7896 13142 7948
rect 13280 7945 13308 7976
rect 13372 7976 14412 8004
rect 14936 7976 15025 8004
rect 13372 7945 13400 7976
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7905 13875 7939
rect 13817 7899 13875 7905
rect 13446 7868 13452 7880
rect 12268 7840 13452 7868
rect 12161 7831 12219 7837
rect 13446 7828 13452 7840
rect 13504 7868 13510 7880
rect 13832 7868 13860 7899
rect 13998 7896 14004 7948
rect 14056 7936 14062 7948
rect 14093 7939 14151 7945
rect 14093 7936 14105 7939
rect 14056 7908 14105 7936
rect 14056 7896 14062 7908
rect 14093 7905 14105 7908
rect 14139 7936 14151 7939
rect 14182 7936 14188 7948
rect 14139 7908 14188 7936
rect 14139 7905 14151 7908
rect 14093 7899 14151 7905
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 14277 7939 14335 7945
rect 14277 7905 14289 7939
rect 14323 7905 14335 7939
rect 14277 7899 14335 7905
rect 13504 7840 13860 7868
rect 13504 7828 13510 7840
rect 13906 7828 13912 7880
rect 13964 7828 13970 7880
rect 12250 7760 12256 7812
rect 12308 7800 12314 7812
rect 12308 7772 12434 7800
rect 12308 7760 12314 7772
rect 4801 7735 4859 7741
rect 4801 7701 4813 7735
rect 4847 7732 4859 7735
rect 5077 7735 5135 7741
rect 5077 7732 5089 7735
rect 4847 7704 5089 7732
rect 4847 7701 4859 7704
rect 4801 7695 4859 7701
rect 5077 7701 5089 7704
rect 5123 7701 5135 7735
rect 5077 7695 5135 7701
rect 8386 7692 8392 7744
rect 8444 7692 8450 7744
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 11146 7732 11152 7744
rect 10836 7704 11152 7732
rect 10836 7692 10842 7704
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11514 7692 11520 7744
rect 11572 7692 11578 7744
rect 11698 7692 11704 7744
rect 11756 7732 11762 7744
rect 12158 7732 12164 7744
rect 11756 7704 12164 7732
rect 11756 7692 11762 7704
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 12406 7732 12434 7772
rect 12710 7760 12716 7812
rect 12768 7800 12774 7812
rect 12768 7772 13216 7800
rect 12768 7760 12774 7772
rect 13081 7735 13139 7741
rect 13081 7732 13093 7735
rect 12406 7704 13093 7732
rect 13081 7701 13093 7704
rect 13127 7701 13139 7735
rect 13188 7732 13216 7772
rect 13262 7760 13268 7812
rect 13320 7800 13326 7812
rect 14292 7800 14320 7899
rect 13320 7772 14320 7800
rect 13320 7760 13326 7772
rect 13541 7735 13599 7741
rect 13541 7732 13553 7735
rect 13188 7704 13553 7732
rect 13081 7695 13139 7701
rect 13541 7701 13553 7704
rect 13587 7701 13599 7735
rect 13541 7695 13599 7701
rect 13998 7692 14004 7744
rect 14056 7692 14062 7744
rect 14384 7732 14412 7976
rect 15013 7973 15025 7976
rect 15059 7973 15071 8007
rect 15120 8004 15148 8032
rect 15212 8004 15240 8044
rect 15381 8041 15393 8044
rect 15427 8041 15439 8075
rect 15381 8035 15439 8041
rect 16574 8032 16580 8084
rect 16632 8032 16638 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 16684 8044 17693 8072
rect 16684 8004 16712 8044
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 17681 8035 17739 8041
rect 15120 7976 15240 8004
rect 15304 7976 15884 8004
rect 15013 7967 15071 7973
rect 14550 7896 14556 7948
rect 14608 7936 14614 7948
rect 14737 7939 14795 7945
rect 14737 7936 14749 7939
rect 14608 7908 14749 7936
rect 14608 7896 14614 7908
rect 14737 7905 14749 7908
rect 14783 7905 14795 7939
rect 14737 7899 14795 7905
rect 14918 7896 14924 7948
rect 14976 7896 14982 7948
rect 15105 7939 15163 7945
rect 15105 7905 15117 7939
rect 15151 7905 15163 7939
rect 15105 7899 15163 7905
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7868 14519 7871
rect 15010 7868 15016 7880
rect 14507 7840 15016 7868
rect 14507 7837 14519 7840
rect 14461 7831 14519 7837
rect 15010 7828 15016 7840
rect 15068 7868 15074 7880
rect 15120 7868 15148 7899
rect 15068 7840 15148 7868
rect 15068 7828 15074 7840
rect 15304 7809 15332 7976
rect 15562 7896 15568 7948
rect 15620 7896 15626 7948
rect 15654 7896 15660 7948
rect 15712 7896 15718 7948
rect 15749 7939 15807 7945
rect 15749 7905 15761 7939
rect 15795 7905 15807 7939
rect 15749 7899 15807 7905
rect 15289 7803 15347 7809
rect 15289 7769 15301 7803
rect 15335 7769 15347 7803
rect 15764 7800 15792 7899
rect 15856 7868 15884 7976
rect 15948 7976 16712 8004
rect 17129 8007 17187 8013
rect 15948 7945 15976 7976
rect 17129 7973 17141 8007
rect 17175 8004 17187 8007
rect 17310 8004 17316 8016
rect 17175 7976 17316 8004
rect 17175 7973 17187 7976
rect 17129 7967 17187 7973
rect 17310 7964 17316 7976
rect 17368 7964 17374 8016
rect 18966 8004 18972 8016
rect 17696 7976 18972 8004
rect 17696 7948 17724 7976
rect 18966 7964 18972 7976
rect 19024 8004 19030 8016
rect 19024 7976 19104 8004
rect 19024 7964 19030 7976
rect 15933 7939 15991 7945
rect 15933 7905 15945 7939
rect 15979 7905 15991 7939
rect 15933 7899 15991 7905
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7905 16175 7939
rect 16117 7899 16175 7905
rect 16132 7868 16160 7899
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 16393 7939 16451 7945
rect 16393 7936 16405 7939
rect 16264 7908 16405 7936
rect 16264 7896 16270 7908
rect 16393 7905 16405 7908
rect 16439 7936 16451 7939
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 16439 7908 16865 7936
rect 16439 7905 16451 7908
rect 16393 7899 16451 7905
rect 16853 7905 16865 7908
rect 16899 7905 16911 7939
rect 16853 7899 16911 7905
rect 17218 7896 17224 7948
rect 17276 7896 17282 7948
rect 17678 7896 17684 7948
rect 17736 7896 17742 7948
rect 18506 7896 18512 7948
rect 18564 7936 18570 7948
rect 19076 7945 19104 7976
rect 18794 7939 18852 7945
rect 18794 7936 18806 7939
rect 18564 7908 18806 7936
rect 18564 7896 18570 7908
rect 18794 7905 18806 7908
rect 18840 7905 18852 7939
rect 18794 7899 18852 7905
rect 19061 7939 19119 7945
rect 19061 7905 19073 7939
rect 19107 7905 19119 7939
rect 19061 7899 19119 7905
rect 15856 7840 16160 7868
rect 16298 7828 16304 7880
rect 16356 7828 16362 7880
rect 15838 7800 15844 7812
rect 15764 7772 15844 7800
rect 15289 7763 15347 7769
rect 15838 7760 15844 7772
rect 15896 7800 15902 7812
rect 18046 7800 18052 7812
rect 15896 7772 18052 7800
rect 15896 7760 15902 7772
rect 18046 7760 18052 7772
rect 18104 7760 18110 7812
rect 15378 7732 15384 7744
rect 14384 7704 15384 7732
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 16390 7692 16396 7744
rect 16448 7692 16454 7744
rect 552 7642 19412 7664
rect 552 7590 2755 7642
rect 2807 7590 2819 7642
rect 2871 7590 2883 7642
rect 2935 7590 2947 7642
rect 2999 7590 3011 7642
rect 3063 7590 7470 7642
rect 7522 7590 7534 7642
rect 7586 7590 7598 7642
rect 7650 7590 7662 7642
rect 7714 7590 7726 7642
rect 7778 7590 12185 7642
rect 12237 7590 12249 7642
rect 12301 7590 12313 7642
rect 12365 7590 12377 7642
rect 12429 7590 12441 7642
rect 12493 7590 16900 7642
rect 16952 7590 16964 7642
rect 17016 7590 17028 7642
rect 17080 7590 17092 7642
rect 17144 7590 17156 7642
rect 17208 7590 19412 7642
rect 552 7568 19412 7590
rect 1026 7488 1032 7540
rect 1084 7488 1090 7540
rect 1305 7531 1363 7537
rect 1305 7497 1317 7531
rect 1351 7528 1363 7531
rect 1578 7528 1584 7540
rect 1351 7500 1584 7528
rect 1351 7497 1363 7500
rect 1305 7491 1363 7497
rect 1121 7327 1179 7333
rect 1121 7293 1133 7327
rect 1167 7324 1179 7327
rect 1320 7324 1348 7491
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2130 7488 2136 7540
rect 2188 7488 2194 7540
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 2590 7528 2596 7540
rect 2455 7500 2596 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2148 7392 2176 7488
rect 1412 7364 2176 7392
rect 1412 7333 1440 7364
rect 1167 7296 1348 7324
rect 1397 7327 1455 7333
rect 1167 7293 1179 7296
rect 1121 7287 1179 7293
rect 1397 7293 1409 7327
rect 1443 7293 1455 7327
rect 1397 7287 1455 7293
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7293 1731 7327
rect 1673 7287 1731 7293
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 2148 7324 2176 7364
rect 1995 7296 2176 7324
rect 2225 7327 2283 7333
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 2424 7324 2452 7491
rect 2590 7488 2596 7500
rect 2648 7528 2654 7540
rect 2685 7531 2743 7537
rect 2685 7528 2697 7531
rect 2648 7500 2697 7528
rect 2648 7488 2654 7500
rect 2685 7497 2697 7500
rect 2731 7497 2743 7531
rect 2685 7491 2743 7497
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 3326 7528 3332 7540
rect 2924 7500 3332 7528
rect 2924 7488 2930 7500
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 5902 7528 5908 7540
rect 5000 7500 5908 7528
rect 4522 7460 4528 7472
rect 3068 7432 4528 7460
rect 2271 7296 2452 7324
rect 2501 7327 2559 7333
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 2501 7293 2513 7327
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 1688 7256 1716 7287
rect 1857 7259 1915 7265
rect 1857 7256 1869 7259
rect 1688 7228 1869 7256
rect 1857 7225 1869 7228
rect 1903 7256 1915 7259
rect 2516 7256 2544 7287
rect 2590 7284 2596 7336
rect 2648 7324 2654 7336
rect 3068 7333 3096 7432
rect 4522 7420 4528 7432
rect 4580 7460 4586 7472
rect 4801 7463 4859 7469
rect 4801 7460 4813 7463
rect 4580 7432 4813 7460
rect 4580 7420 4586 7432
rect 4801 7429 4813 7432
rect 4847 7429 4859 7463
rect 4801 7423 4859 7429
rect 4062 7392 4068 7404
rect 3620 7364 4068 7392
rect 3620 7333 3648 7364
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 5000 7401 5028 7500
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 8202 7528 8208 7540
rect 7055 7500 8208 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 9953 7531 10011 7537
rect 9953 7528 9965 7531
rect 8496 7500 9965 7528
rect 8496 7404 8524 7500
rect 9953 7497 9965 7500
rect 9999 7497 10011 7531
rect 9953 7491 10011 7497
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 11238 7528 11244 7540
rect 10560 7500 11244 7528
rect 10560 7488 10566 7500
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 11330 7488 11336 7540
rect 11388 7528 11394 7540
rect 12434 7528 12440 7540
rect 11388 7500 12440 7528
rect 11388 7488 11394 7500
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 13722 7528 13728 7540
rect 12768 7500 13728 7528
rect 12768 7488 12774 7500
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14093 7531 14151 7537
rect 14093 7528 14105 7531
rect 14056 7500 14105 7528
rect 14056 7488 14062 7500
rect 14093 7497 14105 7500
rect 14139 7497 14151 7531
rect 14093 7491 14151 7497
rect 14182 7488 14188 7540
rect 14240 7528 14246 7540
rect 14461 7531 14519 7537
rect 14461 7528 14473 7531
rect 14240 7500 14473 7528
rect 14240 7488 14246 7500
rect 14461 7497 14473 7500
rect 14507 7497 14519 7531
rect 14461 7491 14519 7497
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 15194 7528 15200 7540
rect 14783 7500 15200 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 10410 7460 10416 7472
rect 8864 7432 10416 7460
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4212 7364 4445 7392
rect 4212 7352 4218 7364
rect 4433 7361 4445 7364
rect 4479 7392 4491 7395
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4479 7364 4997 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 4985 7361 4997 7364
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 6288 7364 6868 7392
rect 2777 7327 2835 7333
rect 2777 7324 2789 7327
rect 2648 7296 2789 7324
rect 2648 7284 2654 7296
rect 2777 7293 2789 7296
rect 2823 7293 2835 7327
rect 2777 7287 2835 7293
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 4890 7284 4896 7336
rect 4948 7284 4954 7336
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 5994 7324 6000 7336
rect 5684 7296 6000 7324
rect 5684 7284 5690 7296
rect 5994 7284 6000 7296
rect 6052 7324 6058 7336
rect 6288 7324 6316 7364
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 6052 7296 6316 7324
rect 6380 7296 6469 7324
rect 6052 7284 6058 7296
rect 3234 7256 3240 7268
rect 1903 7228 2452 7256
rect 2516 7228 3240 7256
rect 1903 7225 1915 7228
rect 1857 7219 1915 7225
rect 1581 7191 1639 7197
rect 1581 7157 1593 7191
rect 1627 7188 1639 7191
rect 2038 7188 2044 7200
rect 1627 7160 2044 7188
rect 1627 7157 1639 7160
rect 1581 7151 1639 7157
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 2424 7188 2452 7228
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 3697 7259 3755 7265
rect 3697 7225 3709 7259
rect 3743 7256 3755 7259
rect 4982 7256 4988 7268
rect 3743 7228 4988 7256
rect 3743 7225 3755 7228
rect 3697 7219 3755 7225
rect 4982 7216 4988 7228
rect 5040 7216 5046 7268
rect 5252 7259 5310 7265
rect 5252 7225 5264 7259
rect 5298 7256 5310 7259
rect 5442 7256 5448 7268
rect 5298 7228 5448 7256
rect 5298 7225 5310 7228
rect 5252 7219 5310 7225
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 2866 7188 2872 7200
rect 2424 7160 2872 7188
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 2961 7191 3019 7197
rect 2961 7157 2973 7191
rect 3007 7188 3019 7191
rect 3142 7188 3148 7200
rect 3007 7160 3148 7188
rect 3007 7157 3019 7160
rect 2961 7151 3019 7157
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7188 3571 7191
rect 4890 7188 4896 7200
rect 3559 7160 4896 7188
rect 3559 7157 3571 7160
rect 3513 7151 3571 7157
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 6380 7197 6408 7296
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 6840 7333 6868 7364
rect 7098 7352 7104 7404
rect 7156 7392 7162 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7156 7364 7941 7392
rect 7156 7352 7162 7364
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8478 7352 8484 7404
rect 8536 7352 8542 7404
rect 8864 7401 8892 7432
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7361 8907 7395
rect 8849 7355 8907 7361
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6604 7296 6653 7324
rect 6604 7284 6610 7296
rect 6641 7293 6653 7296
rect 6687 7293 6699 7327
rect 6641 7287 6699 7293
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 9309 7327 9367 7333
rect 7239 7296 8064 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 6733 7259 6791 7265
rect 6733 7225 6745 7259
rect 6779 7225 6791 7259
rect 6733 7219 6791 7225
rect 6365 7191 6423 7197
rect 6365 7157 6377 7191
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 6748 7188 6776 7219
rect 8036 7200 8064 7296
rect 9309 7293 9321 7327
rect 9355 7324 9367 7327
rect 9508 7324 9536 7432
rect 10410 7420 10416 7432
rect 10468 7460 10474 7472
rect 10468 7432 12020 7460
rect 10468 7420 10474 7432
rect 9355 7296 9536 7324
rect 9692 7364 10088 7392
rect 9355 7293 9367 7296
rect 9309 7287 9367 7293
rect 8757 7259 8815 7265
rect 8757 7225 8769 7259
rect 8803 7225 8815 7259
rect 8757 7219 8815 7225
rect 6512 7160 6776 7188
rect 6512 7148 6518 7160
rect 8018 7148 8024 7200
rect 8076 7148 8082 7200
rect 8570 7148 8576 7200
rect 8628 7148 8634 7200
rect 8772 7188 8800 7219
rect 8846 7216 8852 7268
rect 8904 7256 8910 7268
rect 8941 7259 8999 7265
rect 8941 7256 8953 7259
rect 8904 7228 8953 7256
rect 8904 7216 8910 7228
rect 8941 7225 8953 7228
rect 8987 7225 8999 7259
rect 8941 7219 8999 7225
rect 9030 7216 9036 7268
rect 9088 7216 9094 7268
rect 9217 7259 9275 7265
rect 9217 7225 9229 7259
rect 9263 7256 9275 7259
rect 9692 7256 9720 7364
rect 10060 7336 10088 7364
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7324 9827 7327
rect 9815 7296 9996 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 9968 7268 9996 7296
rect 10042 7284 10048 7336
rect 10100 7324 10106 7336
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 10100 7296 10149 7324
rect 10100 7284 10106 7296
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 10226 7284 10232 7336
rect 10284 7324 10290 7336
rect 10704 7333 10732 7432
rect 11992 7404 12020 7432
rect 12894 7420 12900 7472
rect 12952 7460 12958 7472
rect 13541 7463 13599 7469
rect 13541 7460 13553 7463
rect 12952 7432 13553 7460
rect 12952 7420 12958 7432
rect 13541 7429 13553 7432
rect 13587 7429 13599 7463
rect 13541 7423 13599 7429
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11790 7392 11796 7404
rect 11195 7364 11796 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 11974 7352 11980 7404
rect 12032 7352 12038 7404
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 12526 7392 12532 7404
rect 12207 7364 12532 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 10284 7296 10425 7324
rect 10284 7284 10290 7296
rect 10413 7293 10425 7296
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 10962 7324 10968 7336
rect 10919 7296 10968 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 9263 7228 9720 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 9048 7188 9076 7216
rect 8772 7160 9076 7188
rect 9582 7148 9588 7200
rect 9640 7148 9646 7200
rect 9692 7197 9720 7228
rect 9950 7216 9956 7268
rect 10008 7256 10014 7268
rect 10428 7256 10456 7287
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11238 7284 11244 7336
rect 11296 7284 11302 7336
rect 11514 7284 11520 7336
rect 11572 7324 11578 7336
rect 11609 7327 11667 7333
rect 11609 7324 11621 7327
rect 11572 7296 11621 7324
rect 11572 7284 11578 7296
rect 11609 7293 11621 7296
rect 11655 7293 11667 7327
rect 11609 7287 11667 7293
rect 11146 7256 11152 7268
rect 10008 7228 11152 7256
rect 10008 7216 10014 7228
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 9677 7191 9735 7197
rect 9677 7157 9689 7191
rect 9723 7157 9735 7191
rect 9677 7151 9735 7157
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10229 7191 10287 7197
rect 10229 7188 10241 7191
rect 9916 7160 10241 7188
rect 9916 7148 9922 7160
rect 10229 7157 10241 7160
rect 10275 7188 10287 7191
rect 10410 7188 10416 7200
rect 10275 7160 10416 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 11624 7188 11652 7287
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 11756 7296 11836 7324
rect 11756 7284 11762 7296
rect 11808 7256 11836 7296
rect 11882 7284 11888 7336
rect 11940 7324 11946 7336
rect 12176 7324 12204 7355
rect 12526 7352 12532 7364
rect 12584 7392 12590 7404
rect 12584 7364 12848 7392
rect 12584 7352 12590 7364
rect 12820 7333 12848 7364
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 13173 7395 13231 7401
rect 13173 7392 13185 7395
rect 13044 7364 13185 7392
rect 13044 7352 13050 7364
rect 13173 7361 13185 7364
rect 13219 7361 13231 7395
rect 13173 7355 13231 7361
rect 13262 7352 13268 7404
rect 13320 7392 13326 7404
rect 14016 7392 14044 7488
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 14918 7460 14924 7472
rect 14608 7432 14924 7460
rect 14608 7420 14614 7432
rect 14918 7420 14924 7432
rect 14976 7420 14982 7472
rect 13320 7364 14044 7392
rect 13320 7352 13326 7364
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 15028 7392 15056 7500
rect 15194 7488 15200 7500
rect 15252 7488 15258 7540
rect 16298 7488 16304 7540
rect 16356 7488 16362 7540
rect 18233 7531 18291 7537
rect 18233 7497 18245 7531
rect 18279 7528 18291 7531
rect 18506 7528 18512 7540
rect 18279 7500 18512 7528
rect 18279 7497 18291 7500
rect 18233 7491 18291 7497
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 18874 7488 18880 7540
rect 18932 7488 18938 7540
rect 14240 7364 15056 7392
rect 14240 7352 14246 7364
rect 15838 7352 15844 7404
rect 15896 7352 15902 7404
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7392 18015 7395
rect 18690 7392 18696 7404
rect 18003 7364 18696 7392
rect 18003 7361 18015 7364
rect 17957 7355 18015 7361
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 11940 7296 12204 7324
rect 12253 7327 12311 7333
rect 11940 7284 11946 7296
rect 12253 7293 12265 7327
rect 12299 7293 12311 7327
rect 12253 7287 12311 7293
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 12851 7296 13921 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 13909 7293 13921 7296
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14829 7327 14887 7333
rect 14829 7293 14841 7327
rect 14875 7293 14887 7327
rect 15856 7311 15884 7352
rect 16117 7327 16175 7333
rect 14829 7287 14887 7293
rect 15841 7305 15899 7311
rect 12268 7256 12296 7287
rect 11808 7228 12296 7256
rect 12713 7259 12771 7265
rect 12713 7225 12725 7259
rect 12759 7225 12771 7259
rect 12713 7219 12771 7225
rect 13265 7259 13323 7265
rect 13265 7225 13277 7259
rect 13311 7225 13323 7259
rect 13265 7219 13323 7225
rect 13725 7259 13783 7265
rect 13725 7225 13737 7259
rect 13771 7256 13783 7259
rect 13814 7256 13820 7268
rect 13771 7228 13820 7256
rect 13771 7225 13783 7228
rect 13725 7219 13783 7225
rect 12526 7188 12532 7200
rect 11624 7160 12532 7188
rect 12526 7148 12532 7160
rect 12584 7188 12590 7200
rect 12728 7188 12756 7219
rect 12584 7160 12756 7188
rect 12584 7148 12590 7160
rect 12802 7148 12808 7200
rect 12860 7188 12866 7200
rect 13280 7188 13308 7219
rect 13814 7216 13820 7228
rect 13872 7216 13878 7268
rect 14292 7188 14320 7287
rect 14458 7216 14464 7268
rect 14516 7256 14522 7268
rect 14844 7256 14872 7287
rect 15841 7271 15853 7305
rect 15887 7271 15899 7305
rect 16117 7293 16129 7327
rect 16163 7324 16175 7327
rect 16298 7324 16304 7336
rect 16163 7296 16304 7324
rect 16163 7293 16175 7296
rect 16117 7287 16175 7293
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 17218 7284 17224 7336
rect 17276 7324 17282 7336
rect 17506 7327 17564 7333
rect 17506 7324 17518 7327
rect 17276 7296 17518 7324
rect 17276 7284 17282 7296
rect 17506 7293 17518 7296
rect 17552 7293 17564 7327
rect 17506 7287 17564 7293
rect 17678 7284 17684 7336
rect 17736 7324 17742 7336
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 17736 7296 17785 7324
rect 17736 7284 17742 7296
rect 17773 7293 17785 7296
rect 17819 7293 17831 7327
rect 17773 7287 17831 7293
rect 17862 7284 17868 7336
rect 17920 7284 17926 7336
rect 18325 7327 18383 7333
rect 18325 7293 18337 7327
rect 18371 7324 18383 7327
rect 18708 7324 18736 7352
rect 18777 7327 18835 7333
rect 18777 7324 18789 7327
rect 18371 7296 18644 7324
rect 18708 7296 18789 7324
rect 18371 7293 18383 7296
rect 18325 7287 18383 7293
rect 15841 7265 15899 7271
rect 14516 7228 14872 7256
rect 14516 7216 14522 7228
rect 18616 7200 18644 7296
rect 18777 7293 18789 7296
rect 18823 7293 18835 7327
rect 18777 7287 18835 7293
rect 12860 7160 14320 7188
rect 15933 7191 15991 7197
rect 12860 7148 12866 7160
rect 15933 7157 15945 7191
rect 15979 7188 15991 7191
rect 16393 7191 16451 7197
rect 16393 7188 16405 7191
rect 15979 7160 16405 7188
rect 15979 7157 15991 7160
rect 15933 7151 15991 7157
rect 16393 7157 16405 7160
rect 16439 7157 16451 7191
rect 16393 7151 16451 7157
rect 18598 7148 18604 7200
rect 18656 7148 18662 7200
rect 552 7098 19571 7120
rect 552 7046 5112 7098
rect 5164 7046 5176 7098
rect 5228 7046 5240 7098
rect 5292 7046 5304 7098
rect 5356 7046 5368 7098
rect 5420 7046 9827 7098
rect 9879 7046 9891 7098
rect 9943 7046 9955 7098
rect 10007 7046 10019 7098
rect 10071 7046 10083 7098
rect 10135 7046 14542 7098
rect 14594 7046 14606 7098
rect 14658 7046 14670 7098
rect 14722 7046 14734 7098
rect 14786 7046 14798 7098
rect 14850 7046 19257 7098
rect 19309 7046 19321 7098
rect 19373 7046 19385 7098
rect 19437 7046 19449 7098
rect 19501 7046 19513 7098
rect 19565 7046 19571 7098
rect 552 7024 19571 7046
rect 3234 6944 3240 6996
rect 3292 6984 3298 6996
rect 3329 6987 3387 6993
rect 3329 6984 3341 6987
rect 3292 6956 3341 6984
rect 3292 6944 3298 6956
rect 3329 6953 3341 6956
rect 3375 6953 3387 6987
rect 3329 6947 3387 6953
rect 4062 6944 4068 6996
rect 4120 6944 4126 6996
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 5224 6956 8064 6984
rect 5224 6944 5230 6956
rect 1320 6888 1624 6916
rect 1118 6808 1124 6860
rect 1176 6808 1182 6860
rect 1210 6808 1216 6860
rect 1268 6848 1274 6860
rect 1320 6848 1348 6888
rect 1268 6820 1348 6848
rect 1397 6851 1455 6857
rect 1268 6808 1274 6820
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1486 6848 1492 6860
rect 1443 6820 1492 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 1596 6848 1624 6888
rect 1653 6851 1711 6857
rect 1653 6848 1665 6851
rect 1596 6820 1665 6848
rect 1653 6817 1665 6820
rect 1699 6817 1711 6851
rect 1653 6811 1711 6817
rect 2590 6808 2596 6860
rect 2648 6848 2654 6860
rect 4080 6857 4108 6944
rect 8036 6928 8064 6956
rect 8386 6944 8392 6996
rect 8444 6944 8450 6996
rect 9861 6987 9919 6993
rect 9861 6984 9873 6987
rect 8956 6956 9873 6984
rect 4890 6876 4896 6928
rect 4948 6876 4954 6928
rect 6104 6888 6316 6916
rect 2953 6851 3011 6857
rect 2953 6848 2965 6851
rect 2648 6820 2965 6848
rect 2648 6808 2654 6820
rect 2953 6817 2965 6820
rect 2999 6817 3011 6851
rect 2953 6811 3011 6817
rect 3421 6851 3479 6857
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 3697 6851 3755 6857
rect 3467 6820 3648 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 934 6672 940 6724
rect 992 6712 998 6724
rect 1394 6712 1400 6724
rect 992 6684 1400 6712
rect 992 6672 998 6684
rect 1394 6672 1400 6684
rect 1452 6672 1458 6724
rect 2777 6715 2835 6721
rect 2777 6681 2789 6715
rect 2823 6712 2835 6715
rect 3510 6712 3516 6724
rect 2823 6684 3516 6712
rect 2823 6681 2835 6684
rect 2777 6675 2835 6681
rect 3510 6672 3516 6684
rect 3568 6672 3574 6724
rect 1029 6647 1087 6653
rect 1029 6644 1041 6647
rect 492 6616 1041 6644
rect 492 6440 520 6616
rect 1029 6613 1041 6616
rect 1075 6613 1087 6647
rect 1029 6607 1087 6613
rect 1118 6604 1124 6656
rect 1176 6644 1182 6656
rect 1578 6644 1584 6656
rect 1176 6616 1584 6644
rect 1176 6604 1182 6616
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 3142 6644 3148 6656
rect 3099 6616 3148 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 3620 6653 3648 6820
rect 3697 6817 3709 6851
rect 3743 6817 3755 6851
rect 3697 6811 3755 6817
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 3712 6780 3740 6811
rect 4154 6808 4160 6860
rect 4212 6808 4218 6860
rect 4424 6851 4482 6857
rect 4424 6817 4436 6851
rect 4470 6848 4482 6851
rect 4908 6848 4936 6876
rect 6104 6848 6132 6888
rect 6178 6857 6184 6860
rect 4470 6820 4936 6848
rect 5460 6820 6132 6848
rect 4470 6817 4482 6820
rect 4424 6811 4482 6817
rect 3712 6752 4108 6780
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 3970 6644 3976 6656
rect 3651 6616 3976 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4080 6644 4108 6752
rect 5460 6656 5488 6820
rect 6172 6811 6184 6857
rect 6178 6808 6184 6811
rect 6236 6808 6242 6860
rect 6288 6848 6316 6888
rect 8018 6876 8024 6928
rect 8076 6876 8082 6928
rect 8404 6916 8432 6944
rect 8665 6919 8723 6925
rect 8665 6916 8677 6919
rect 8404 6888 8677 6916
rect 8665 6885 8677 6888
rect 8711 6885 8723 6919
rect 8665 6879 8723 6885
rect 8956 6860 8984 6956
rect 9861 6953 9873 6956
rect 9907 6953 9919 6987
rect 12618 6984 12624 6996
rect 9861 6947 9919 6953
rect 11532 6956 11836 6984
rect 9674 6876 9680 6928
rect 9732 6916 9738 6928
rect 11532 6916 11560 6956
rect 11698 6916 11704 6928
rect 9732 6888 10456 6916
rect 9732 6876 9738 6888
rect 6288 6820 7328 6848
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 4430 6644 4436 6656
rect 4080 6616 4436 6644
rect 4430 6604 4436 6616
rect 4488 6604 4494 6656
rect 5442 6604 5448 6656
rect 5500 6604 5506 6656
rect 5534 6604 5540 6656
rect 5592 6604 5598 6656
rect 5920 6644 5948 6743
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7300 6780 7328 6820
rect 7374 6808 7380 6860
rect 7432 6848 7438 6860
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7432 6820 7665 6848
rect 7432 6808 7438 6820
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 8386 6808 8392 6860
rect 8444 6808 8450 6860
rect 8478 6808 8484 6860
rect 8536 6848 8542 6860
rect 8573 6851 8631 6857
rect 8573 6848 8585 6851
rect 8536 6820 8585 6848
rect 8536 6808 8542 6820
rect 8573 6817 8585 6820
rect 8619 6817 8631 6851
rect 8573 6811 8631 6817
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6848 8815 6851
rect 8938 6848 8944 6860
rect 8803 6820 8944 6848
rect 8803 6817 8815 6820
rect 8757 6811 8815 6817
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 9033 6851 9091 6857
rect 9033 6817 9045 6851
rect 9079 6817 9091 6851
rect 9033 6811 9091 6817
rect 9048 6780 9076 6811
rect 9122 6808 9128 6860
rect 9180 6848 9186 6860
rect 9217 6851 9275 6857
rect 9217 6848 9229 6851
rect 9180 6820 9229 6848
rect 9180 6808 9186 6820
rect 9217 6817 9229 6820
rect 9263 6817 9275 6851
rect 9217 6811 9275 6817
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 6972 6752 7236 6780
rect 7300 6752 9076 6780
rect 9324 6780 9352 6811
rect 9398 6808 9404 6860
rect 9456 6808 9462 6860
rect 9953 6851 10011 6857
rect 9953 6817 9965 6851
rect 9999 6848 10011 6851
rect 9999 6820 10180 6848
rect 9999 6817 10011 6820
rect 9953 6811 10011 6817
rect 9582 6780 9588 6792
rect 9324 6752 9588 6780
rect 6972 6740 6978 6752
rect 7098 6672 7104 6724
rect 7156 6672 7162 6724
rect 7208 6712 7236 6752
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 7561 6715 7619 6721
rect 7561 6712 7573 6715
rect 7208 6684 7573 6712
rect 7561 6681 7573 6684
rect 7607 6681 7619 6715
rect 7561 6675 7619 6681
rect 9214 6672 9220 6724
rect 9272 6712 9278 6724
rect 10152 6712 10180 6820
rect 10226 6808 10232 6860
rect 10284 6808 10290 6860
rect 10428 6857 10456 6888
rect 11440 6888 11560 6916
rect 11624 6888 11704 6916
rect 10413 6851 10471 6857
rect 10413 6817 10425 6851
rect 10459 6848 10471 6851
rect 10962 6848 10968 6860
rect 10459 6820 10968 6848
rect 10459 6817 10471 6820
rect 10413 6811 10471 6817
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11440 6857 11468 6888
rect 11624 6857 11652 6888
rect 11698 6876 11704 6888
rect 11756 6876 11762 6928
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6817 11483 6851
rect 11425 6811 11483 6817
rect 11609 6851 11667 6857
rect 11609 6817 11621 6851
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 11238 6780 11244 6792
rect 10827 6752 11244 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 11532 6712 11560 6740
rect 9272 6684 9628 6712
rect 10152 6684 11560 6712
rect 9272 6672 9278 6684
rect 7116 6644 7144 6672
rect 5920 6616 7144 6644
rect 7282 6604 7288 6656
rect 7340 6604 7346 6656
rect 8941 6647 8999 6653
rect 8941 6613 8953 6647
rect 8987 6644 8999 6647
rect 9398 6644 9404 6656
rect 8987 6616 9404 6644
rect 8987 6613 8999 6616
rect 8941 6607 8999 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9600 6653 9628 6684
rect 11164 6656 11192 6684
rect 9585 6647 9643 6653
rect 9585 6613 9597 6647
rect 9631 6613 9643 6647
rect 9585 6607 9643 6613
rect 11146 6604 11152 6656
rect 11204 6604 11210 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11624 6644 11652 6811
rect 11701 6783 11759 6789
rect 11701 6749 11713 6783
rect 11747 6749 11759 6783
rect 11808 6780 11836 6956
rect 12452 6956 12624 6984
rect 11885 6919 11943 6925
rect 11885 6885 11897 6919
rect 11931 6885 11943 6919
rect 11885 6879 11943 6885
rect 11900 6848 11928 6879
rect 12452 6848 12480 6956
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 13357 6987 13415 6993
rect 13357 6953 13369 6987
rect 13403 6984 13415 6987
rect 13906 6984 13912 6996
rect 13403 6956 13912 6984
rect 13403 6953 13415 6956
rect 13357 6947 13415 6953
rect 11900 6820 12480 6848
rect 12526 6808 12532 6860
rect 12584 6808 12590 6860
rect 12618 6808 12624 6860
rect 12676 6848 12682 6860
rect 12802 6848 12808 6860
rect 12676 6820 12808 6848
rect 12676 6808 12682 6820
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 13173 6851 13231 6857
rect 13173 6848 13185 6851
rect 12952 6820 13185 6848
rect 12952 6808 12958 6820
rect 13173 6817 13185 6820
rect 13219 6817 13231 6851
rect 13173 6811 13231 6817
rect 13262 6808 13268 6860
rect 13320 6808 13326 6860
rect 11882 6780 11888 6792
rect 11808 6752 11888 6780
rect 11701 6743 11759 6749
rect 11296 6616 11652 6644
rect 11716 6644 11744 6743
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 12032 6752 12081 6780
rect 12032 6740 12038 6752
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6780 12219 6783
rect 12710 6780 12716 6792
rect 12207 6752 12716 6780
rect 12207 6749 12219 6752
rect 12161 6743 12219 6749
rect 12084 6712 12112 6743
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6780 13139 6783
rect 13280 6780 13308 6808
rect 13127 6752 13308 6780
rect 13127 6749 13139 6752
rect 13081 6743 13139 6749
rect 13372 6712 13400 6947
rect 13906 6944 13912 6956
rect 13964 6944 13970 6996
rect 17494 6944 17500 6996
rect 17552 6944 17558 6996
rect 16206 6916 16212 6928
rect 12084 6684 13400 6712
rect 13556 6888 16212 6916
rect 13170 6644 13176 6656
rect 11716 6616 13176 6644
rect 11296 6604 11302 6616
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 13262 6604 13268 6656
rect 13320 6644 13326 6656
rect 13556 6644 13584 6888
rect 16206 6876 16212 6888
rect 16264 6876 16270 6928
rect 16485 6919 16543 6925
rect 16485 6885 16497 6919
rect 16531 6916 16543 6919
rect 18046 6916 18052 6928
rect 16531 6888 18052 6916
rect 16531 6885 16543 6888
rect 16485 6879 16543 6885
rect 18046 6876 18052 6888
rect 18104 6876 18110 6928
rect 13900 6851 13958 6857
rect 13900 6817 13912 6851
rect 13946 6848 13958 6851
rect 14458 6848 14464 6860
rect 13946 6820 14464 6848
rect 13946 6817 13958 6820
rect 13900 6811 13958 6817
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 16666 6848 16672 6860
rect 15252 6820 16672 6848
rect 15252 6808 15258 6820
rect 16666 6808 16672 6820
rect 16724 6848 16730 6860
rect 17221 6851 17279 6857
rect 17221 6848 17233 6851
rect 16724 6820 17233 6848
rect 16724 6808 16730 6820
rect 17221 6817 17233 6820
rect 17267 6817 17279 6851
rect 17221 6811 17279 6817
rect 18598 6808 18604 6860
rect 18656 6857 18662 6860
rect 18656 6848 18668 6857
rect 18877 6851 18935 6857
rect 18656 6820 18701 6848
rect 18656 6811 18668 6820
rect 18877 6817 18889 6851
rect 18923 6848 18935 6851
rect 18966 6848 18972 6860
rect 18923 6820 18972 6848
rect 18923 6817 18935 6820
rect 18877 6811 18935 6817
rect 18656 6808 18662 6811
rect 18966 6808 18972 6820
rect 19024 6808 19030 6860
rect 13630 6740 13636 6792
rect 13688 6740 13694 6792
rect 13320 6616 13584 6644
rect 13320 6604 13326 6616
rect 15010 6604 15016 6656
rect 15068 6604 15074 6656
rect 552 6554 19412 6576
rect 552 6502 2755 6554
rect 2807 6502 2819 6554
rect 2871 6502 2883 6554
rect 2935 6502 2947 6554
rect 2999 6502 3011 6554
rect 3063 6502 7470 6554
rect 7522 6502 7534 6554
rect 7586 6502 7598 6554
rect 7650 6502 7662 6554
rect 7714 6502 7726 6554
rect 7778 6502 12185 6554
rect 12237 6502 12249 6554
rect 12301 6502 12313 6554
rect 12365 6502 12377 6554
rect 12429 6502 12441 6554
rect 12493 6502 16900 6554
rect 16952 6502 16964 6554
rect 17016 6502 17028 6554
rect 17080 6502 17092 6554
rect 17144 6502 17156 6554
rect 17208 6502 19412 6554
rect 552 6480 19412 6502
rect 1213 6443 1271 6449
rect 1213 6440 1225 6443
rect 492 6412 1225 6440
rect 1213 6409 1225 6412
rect 1259 6409 1271 6443
rect 1213 6403 1271 6409
rect 937 6375 995 6381
rect 937 6341 949 6375
rect 983 6372 995 6375
rect 1026 6372 1032 6384
rect 983 6344 1032 6372
rect 983 6341 995 6344
rect 937 6335 995 6341
rect 1026 6332 1032 6344
rect 1084 6332 1090 6384
rect 1228 6372 1256 6403
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 2961 6443 3019 6449
rect 1452 6412 2176 6440
rect 1452 6400 1458 6412
rect 1228 6344 1440 6372
rect 1412 6304 1440 6344
rect 1412 6276 1900 6304
rect 1872 6248 1900 6276
rect 934 6196 940 6248
rect 992 6236 998 6248
rect 1029 6239 1087 6245
rect 1029 6236 1041 6239
rect 992 6208 1041 6236
rect 992 6196 998 6208
rect 1029 6205 1041 6208
rect 1075 6205 1087 6239
rect 1029 6199 1087 6205
rect 1302 6196 1308 6248
rect 1360 6196 1366 6248
rect 1578 6196 1584 6248
rect 1636 6196 1642 6248
rect 1854 6196 1860 6248
rect 1912 6196 1918 6248
rect 2148 6245 2176 6412
rect 2961 6409 2973 6443
rect 3007 6440 3019 6443
rect 3234 6440 3240 6452
rect 3007 6412 3240 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 3510 6400 3516 6452
rect 3568 6400 3574 6452
rect 5534 6400 5540 6452
rect 5592 6400 5598 6452
rect 7098 6440 7104 6452
rect 6840 6412 7104 6440
rect 3528 6372 3556 6400
rect 5442 6372 5448 6384
rect 3528 6344 5448 6372
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 3510 6304 3516 6316
rect 3068 6276 3516 6304
rect 3068 6245 3096 6276
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6205 2191 6239
rect 2133 6199 2191 6205
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6205 3111 6239
rect 3053 6199 3111 6205
rect 3142 6196 3148 6248
rect 3200 6236 3206 6248
rect 3970 6245 3976 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3200 6208 3433 6236
rect 3200 6196 3206 6208
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3965 6236 3976 6245
rect 3931 6208 3976 6236
rect 3421 6199 3479 6205
rect 3965 6199 3976 6208
rect 3970 6196 3976 6199
rect 4028 6196 4034 6248
rect 4890 6196 4896 6248
rect 4948 6196 4954 6248
rect 4985 6239 5043 6245
rect 4985 6205 4997 6239
rect 5031 6236 5043 6239
rect 5166 6236 5172 6248
rect 5031 6208 5172 6236
rect 5031 6205 5043 6208
rect 4985 6199 5043 6205
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6205 5319 6239
rect 5552 6236 5580 6400
rect 6840 6313 6868 6412
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 9122 6400 9128 6452
rect 9180 6440 9186 6452
rect 9582 6440 9588 6452
rect 9180 6412 9588 6440
rect 9180 6400 9186 6412
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 12158 6440 12164 6452
rect 10468 6412 12164 6440
rect 10468 6400 10474 6412
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 15746 6440 15752 6452
rect 12584 6412 15752 6440
rect 12584 6400 12590 6412
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 15841 6443 15899 6449
rect 15841 6409 15853 6443
rect 15887 6440 15899 6443
rect 16117 6443 16175 6449
rect 16117 6440 16129 6443
rect 15887 6412 16129 6440
rect 15887 6409 15899 6412
rect 15841 6403 15899 6409
rect 16117 6409 16129 6412
rect 16163 6409 16175 6443
rect 16117 6403 16175 6409
rect 16482 6400 16488 6452
rect 16540 6400 16546 6452
rect 18138 6400 18144 6452
rect 18196 6440 18202 6452
rect 18417 6443 18475 6449
rect 18417 6440 18429 6443
rect 18196 6412 18429 6440
rect 18196 6400 18202 6412
rect 18417 6409 18429 6412
rect 18463 6409 18475 6443
rect 18417 6403 18475 6409
rect 9306 6332 9312 6384
rect 9364 6372 9370 6384
rect 9401 6375 9459 6381
rect 9401 6372 9413 6375
rect 9364 6344 9413 6372
rect 9364 6332 9370 6344
rect 9401 6341 9413 6344
rect 9447 6341 9459 6375
rect 10962 6372 10968 6384
rect 9401 6335 9459 6341
rect 9488 6344 10968 6372
rect 6825 6307 6883 6313
rect 5828 6276 6592 6304
rect 5629 6239 5687 6245
rect 5629 6236 5641 6239
rect 5552 6208 5641 6236
rect 5261 6199 5319 6205
rect 5629 6205 5641 6208
rect 5675 6205 5687 6239
rect 5629 6199 5687 6205
rect 1949 6171 2007 6177
rect 1949 6168 1961 6171
rect 1228 6140 1961 6168
rect 1228 6112 1256 6140
rect 1949 6137 1961 6140
rect 1995 6168 2007 6171
rect 2225 6171 2283 6177
rect 2225 6168 2237 6171
rect 1995 6140 2237 6168
rect 1995 6137 2007 6140
rect 1949 6131 2007 6137
rect 2225 6137 2237 6140
rect 2271 6137 2283 6171
rect 2225 6131 2283 6137
rect 4246 6128 4252 6180
rect 4304 6128 4310 6180
rect 4908 6168 4936 6196
rect 5276 6168 5304 6199
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 5828 6245 5856 6276
rect 6564 6248 6592 6276
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 9488 6304 9516 6344
rect 10962 6332 10968 6344
rect 11020 6332 11026 6384
rect 13814 6332 13820 6384
rect 13872 6372 13878 6384
rect 13872 6344 14780 6372
rect 13872 6332 13878 6344
rect 6825 6267 6883 6273
rect 8312 6276 9516 6304
rect 5813 6239 5871 6245
rect 5813 6236 5825 6239
rect 5776 6208 5825 6236
rect 5776 6196 5782 6208
rect 5813 6205 5825 6208
rect 5859 6205 5871 6239
rect 5813 6199 5871 6205
rect 5994 6196 6000 6248
rect 6052 6196 6058 6248
rect 6546 6196 6552 6248
rect 6604 6196 6610 6248
rect 7092 6239 7150 6245
rect 7092 6205 7104 6239
rect 7138 6236 7150 6239
rect 7374 6236 7380 6248
rect 7138 6208 7380 6236
rect 7138 6205 7150 6208
rect 7092 6199 7150 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 8312 6236 8340 6276
rect 9582 6264 9588 6316
rect 9640 6304 9646 6316
rect 10778 6304 10784 6316
rect 9640 6276 10784 6304
rect 9640 6264 9646 6276
rect 10778 6264 10784 6276
rect 10836 6304 10842 6316
rect 11425 6307 11483 6313
rect 10836 6276 11275 6304
rect 10836 6264 10842 6276
rect 7760 6208 8340 6236
rect 4908 6140 5304 6168
rect 5902 6128 5908 6180
rect 5960 6128 5966 6180
rect 6564 6168 6592 6196
rect 7760 6168 7788 6208
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8444 6208 8861 6236
rect 8444 6196 8450 6208
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8849 6199 8907 6205
rect 8956 6208 9137 6236
rect 6564 6140 7788 6168
rect 7834 6128 7840 6180
rect 7892 6168 7898 6180
rect 8956 6168 8984 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 9217 6239 9275 6245
rect 9217 6205 9229 6239
rect 9263 6236 9275 6239
rect 9674 6236 9680 6248
rect 9263 6208 9680 6236
rect 9263 6205 9275 6208
rect 9217 6199 9275 6205
rect 9674 6196 9680 6208
rect 9732 6236 9738 6248
rect 11149 6239 11207 6245
rect 11149 6236 11161 6239
rect 9732 6208 11161 6236
rect 9732 6196 9738 6208
rect 11149 6205 11161 6208
rect 11195 6205 11207 6239
rect 11247 6236 11275 6276
rect 11425 6273 11437 6307
rect 11471 6304 11483 6307
rect 11514 6304 11520 6316
rect 11471 6276 11520 6304
rect 11471 6273 11483 6276
rect 11425 6267 11483 6273
rect 11514 6264 11520 6276
rect 11572 6304 11578 6316
rect 11974 6304 11980 6316
rect 11572 6276 11980 6304
rect 11572 6264 11578 6276
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 13446 6304 13452 6316
rect 12492 6276 13452 6304
rect 12492 6264 12498 6276
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 13740 6276 14657 6304
rect 11247 6208 11560 6236
rect 11149 6199 11207 6205
rect 7892 6140 8984 6168
rect 9033 6171 9091 6177
rect 7892 6128 7898 6140
rect 9033 6137 9045 6171
rect 9079 6137 9091 6171
rect 9033 6131 9091 6137
rect 1210 6060 1216 6112
rect 1268 6060 1274 6112
rect 1302 6060 1308 6112
rect 1360 6100 1366 6112
rect 1673 6103 1731 6109
rect 1673 6100 1685 6103
rect 1360 6072 1685 6100
rect 1360 6060 1366 6072
rect 1673 6069 1685 6072
rect 1719 6069 1731 6103
rect 1673 6063 1731 6069
rect 2590 6060 2596 6112
rect 2648 6100 2654 6112
rect 3881 6103 3939 6109
rect 3881 6100 3893 6103
rect 2648 6072 3893 6100
rect 2648 6060 2654 6072
rect 3881 6069 3893 6072
rect 3927 6100 3939 6103
rect 5169 6103 5227 6109
rect 5169 6100 5181 6103
rect 3927 6072 5181 6100
rect 3927 6069 3939 6072
rect 3881 6063 3939 6069
rect 5169 6069 5181 6072
rect 5215 6100 5227 6103
rect 5442 6100 5448 6112
rect 5215 6072 5448 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 6181 6103 6239 6109
rect 6181 6069 6193 6103
rect 6227 6100 6239 6103
rect 7006 6100 7012 6112
rect 6227 6072 7012 6100
rect 6227 6069 6239 6072
rect 6181 6063 6239 6069
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 8202 6060 8208 6112
rect 8260 6060 8266 6112
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 9048 6100 9076 6131
rect 9398 6128 9404 6180
rect 9456 6168 9462 6180
rect 11532 6177 11560 6208
rect 11882 6196 11888 6248
rect 11940 6196 11946 6248
rect 12986 6196 12992 6248
rect 13044 6236 13050 6248
rect 13630 6236 13636 6248
rect 13044 6208 13636 6236
rect 13044 6196 13050 6208
rect 13630 6196 13636 6208
rect 13688 6236 13694 6248
rect 13740 6236 13768 6276
rect 14645 6273 14657 6276
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 13688 6208 13768 6236
rect 13688 6196 13694 6208
rect 13906 6196 13912 6248
rect 13964 6236 13970 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13964 6208 14105 6236
rect 13964 6196 13970 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 14185 6239 14243 6245
rect 14185 6205 14197 6239
rect 14231 6205 14243 6239
rect 14185 6199 14243 6205
rect 14277 6239 14335 6245
rect 14277 6205 14289 6239
rect 14323 6205 14335 6239
rect 14277 6199 14335 6205
rect 11517 6171 11575 6177
rect 9456 6140 11468 6168
rect 9456 6128 9462 6140
rect 9582 6100 9588 6112
rect 8628 6072 9588 6100
rect 8628 6060 8634 6072
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 11440 6100 11468 6140
rect 11517 6137 11529 6171
rect 11563 6168 11575 6171
rect 11606 6168 11612 6180
rect 11563 6140 11612 6168
rect 11563 6137 11575 6140
rect 11517 6131 11575 6137
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 11790 6128 11796 6180
rect 11848 6168 11854 6180
rect 11977 6171 12035 6177
rect 11977 6168 11989 6171
rect 11848 6140 11989 6168
rect 11848 6128 11854 6140
rect 11977 6137 11989 6140
rect 12023 6168 12035 6171
rect 12618 6168 12624 6180
rect 12023 6140 12624 6168
rect 12023 6137 12035 6140
rect 11977 6131 12035 6137
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 12802 6128 12808 6180
rect 12860 6168 12866 6180
rect 14200 6168 14228 6199
rect 12860 6140 14228 6168
rect 14292 6168 14320 6199
rect 14458 6196 14464 6248
rect 14516 6196 14522 6248
rect 14752 6168 14780 6344
rect 15470 6332 15476 6384
rect 15528 6372 15534 6384
rect 16025 6375 16083 6381
rect 15528 6344 15976 6372
rect 15528 6332 15534 6344
rect 15562 6264 15568 6316
rect 15620 6264 15626 6316
rect 15580 6236 15608 6264
rect 15166 6208 15700 6236
rect 15166 6168 15194 6208
rect 14292 6140 15194 6168
rect 15473 6171 15531 6177
rect 12860 6128 12866 6140
rect 15473 6137 15485 6171
rect 15519 6137 15531 6171
rect 15473 6131 15531 6137
rect 13262 6100 13268 6112
rect 11440 6072 13268 6100
rect 13262 6060 13268 6072
rect 13320 6060 13326 6112
rect 13909 6103 13967 6109
rect 13909 6069 13921 6103
rect 13955 6100 13967 6103
rect 14458 6100 14464 6112
rect 13955 6072 14464 6100
rect 13955 6069 13967 6072
rect 13909 6063 13967 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 15488 6100 15516 6131
rect 15562 6128 15568 6180
rect 15620 6128 15626 6180
rect 15672 6168 15700 6208
rect 15746 6196 15752 6248
rect 15804 6196 15810 6248
rect 15838 6196 15844 6248
rect 15896 6196 15902 6248
rect 15948 6236 15976 6344
rect 16025 6341 16037 6375
rect 16071 6372 16083 6375
rect 16500 6372 16528 6400
rect 16071 6344 16528 6372
rect 16071 6341 16083 6344
rect 16025 6335 16083 6341
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 18598 6304 18604 6316
rect 16172 6276 16436 6304
rect 16172 6264 16178 6276
rect 16408 6245 16436 6276
rect 18248 6276 18604 6304
rect 16301 6239 16359 6245
rect 16301 6236 16313 6239
rect 15948 6208 16313 6236
rect 16301 6205 16313 6208
rect 16347 6205 16359 6239
rect 16301 6199 16359 6205
rect 16393 6239 16451 6245
rect 16393 6205 16405 6239
rect 16439 6205 16451 6239
rect 16393 6199 16451 6205
rect 16666 6196 16672 6248
rect 16724 6196 16730 6248
rect 17218 6196 17224 6248
rect 17276 6196 17282 6248
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6236 17371 6239
rect 17770 6236 17776 6248
rect 17359 6208 17776 6236
rect 17359 6205 17371 6208
rect 17313 6199 17371 6205
rect 17770 6196 17776 6208
rect 17828 6196 17834 6248
rect 18248 6245 18276 6276
rect 18598 6264 18604 6276
rect 18656 6304 18662 6316
rect 18785 6307 18843 6313
rect 18785 6304 18797 6307
rect 18656 6276 18797 6304
rect 18656 6264 18662 6276
rect 18785 6273 18797 6276
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6236 17923 6239
rect 18233 6239 18291 6245
rect 18233 6236 18245 6239
rect 17911 6208 18245 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 18233 6205 18245 6208
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 18322 6196 18328 6248
rect 18380 6196 18386 6248
rect 18414 6196 18420 6248
rect 18472 6236 18478 6248
rect 18693 6239 18751 6245
rect 18693 6236 18705 6239
rect 18472 6208 18705 6236
rect 18472 6196 18478 6208
rect 18693 6205 18705 6208
rect 18739 6205 18751 6239
rect 18693 6199 18751 6205
rect 16485 6171 16543 6177
rect 16485 6168 16497 6171
rect 15672 6140 16497 6168
rect 16485 6137 16497 6140
rect 16531 6137 16543 6171
rect 16485 6131 16543 6137
rect 15252 6072 15516 6100
rect 15252 6060 15258 6072
rect 552 6010 19571 6032
rect 552 5958 5112 6010
rect 5164 5958 5176 6010
rect 5228 5958 5240 6010
rect 5292 5958 5304 6010
rect 5356 5958 5368 6010
rect 5420 5958 9827 6010
rect 9879 5958 9891 6010
rect 9943 5958 9955 6010
rect 10007 5958 10019 6010
rect 10071 5958 10083 6010
rect 10135 5958 14542 6010
rect 14594 5958 14606 6010
rect 14658 5958 14670 6010
rect 14722 5958 14734 6010
rect 14786 5958 14798 6010
rect 14850 5958 19257 6010
rect 19309 5958 19321 6010
rect 19373 5958 19385 6010
rect 19437 5958 19449 6010
rect 19501 5958 19513 6010
rect 19565 5958 19571 6010
rect 552 5936 19571 5958
rect 1302 5856 1308 5908
rect 1360 5896 1366 5908
rect 1397 5899 1455 5905
rect 1397 5896 1409 5899
rect 1360 5868 1409 5896
rect 1360 5856 1366 5868
rect 1397 5865 1409 5868
rect 1443 5865 1455 5899
rect 1397 5859 1455 5865
rect 1854 5856 1860 5908
rect 1912 5856 1918 5908
rect 1946 5856 1952 5908
rect 2004 5856 2010 5908
rect 2961 5899 3019 5905
rect 2961 5865 2973 5899
rect 3007 5896 3019 5899
rect 3326 5896 3332 5908
rect 3007 5868 3332 5896
rect 3007 5865 3019 5868
rect 2961 5859 3019 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 6362 5856 6368 5908
rect 6420 5856 6426 5908
rect 6822 5856 6828 5908
rect 6880 5856 6886 5908
rect 8202 5856 8208 5908
rect 8260 5856 8266 5908
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 8846 5896 8852 5908
rect 8435 5868 8852 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 8996 5868 9321 5896
rect 8996 5856 9002 5868
rect 1872 5828 1900 5856
rect 1780 5800 1900 5828
rect 1780 5769 1808 5800
rect 1305 5763 1363 5769
rect 1305 5729 1317 5763
rect 1351 5729 1363 5763
rect 1305 5723 1363 5729
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5729 1823 5763
rect 1765 5723 1823 5729
rect 1210 5652 1216 5704
rect 1268 5692 1274 5704
rect 1320 5692 1348 5723
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 1964 5760 1992 5856
rect 3160 5800 4200 5828
rect 3160 5769 3188 5800
rect 4172 5772 4200 5800
rect 4890 5788 4896 5840
rect 4948 5828 4954 5840
rect 6089 5831 6147 5837
rect 6089 5828 6101 5831
rect 4948 5800 6101 5828
rect 4948 5788 4954 5800
rect 6089 5797 6101 5800
rect 6135 5797 6147 5831
rect 6840 5828 6868 5856
rect 7254 5831 7312 5837
rect 7254 5828 7266 5831
rect 6840 5800 7266 5828
rect 6089 5791 6147 5797
rect 7254 5797 7266 5800
rect 7300 5797 7312 5831
rect 8220 5828 8248 5856
rect 8757 5831 8815 5837
rect 8757 5828 8769 5831
rect 8220 5800 8769 5828
rect 7254 5791 7312 5797
rect 8757 5797 8769 5800
rect 8803 5797 8815 5831
rect 8757 5791 8815 5797
rect 3418 5769 3424 5772
rect 1912 5732 1992 5760
rect 3145 5763 3203 5769
rect 3053 5753 3111 5759
rect 1912 5720 1918 5732
rect 3053 5719 3065 5753
rect 3099 5719 3111 5753
rect 3145 5729 3157 5763
rect 3191 5729 3203 5763
rect 3412 5760 3424 5769
rect 3379 5732 3424 5760
rect 3145 5723 3203 5729
rect 3412 5723 3424 5732
rect 3418 5720 3424 5723
rect 3476 5720 3482 5772
rect 4154 5720 4160 5772
rect 4212 5720 4218 5772
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5729 4675 5763
rect 4617 5723 4675 5729
rect 3053 5713 3111 5719
rect 1268 5664 1348 5692
rect 1268 5652 1274 5664
rect 1670 5516 1676 5568
rect 1728 5516 1734 5568
rect 1946 5516 1952 5568
rect 2004 5516 2010 5568
rect 3068 5556 3096 5713
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 4632 5692 4660 5723
rect 5718 5720 5724 5772
rect 5776 5720 5782 5772
rect 5810 5720 5816 5772
rect 5868 5720 5874 5772
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5729 6055 5763
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 5997 5723 6055 5729
rect 6104 5732 6193 5760
rect 4488 5664 4660 5692
rect 5736 5692 5764 5720
rect 6012 5692 6040 5723
rect 6104 5704 6132 5732
rect 6181 5729 6193 5732
rect 6227 5760 6239 5763
rect 6730 5760 6736 5772
rect 6227 5732 6736 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 6822 5720 6828 5772
rect 6880 5760 6886 5772
rect 7009 5763 7067 5769
rect 7009 5760 7021 5763
rect 6880 5732 7021 5760
rect 6880 5720 6886 5732
rect 7009 5729 7021 5732
rect 7055 5760 7067 5763
rect 7098 5760 7104 5772
rect 7055 5732 7104 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 8478 5720 8484 5772
rect 8536 5720 8542 5772
rect 8570 5720 8576 5772
rect 8628 5760 8634 5772
rect 8665 5763 8723 5769
rect 8665 5760 8677 5763
rect 8628 5732 8677 5760
rect 8628 5720 8634 5732
rect 8665 5729 8677 5732
rect 8711 5729 8723 5763
rect 8665 5723 8723 5729
rect 8849 5763 8907 5769
rect 8849 5729 8861 5763
rect 8895 5758 8907 5763
rect 8956 5758 8984 5856
rect 9293 5828 9321 5868
rect 9398 5856 9404 5908
rect 9456 5896 9462 5908
rect 10778 5896 10784 5908
rect 9456 5868 10784 5896
rect 9456 5856 9462 5868
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 11698 5896 11704 5908
rect 11247 5868 11704 5896
rect 9293 5800 9536 5828
rect 8895 5730 8984 5758
rect 8895 5729 8907 5730
rect 8849 5723 8907 5729
rect 5736 5664 6040 5692
rect 4488 5652 4494 5664
rect 6086 5652 6092 5704
rect 6144 5652 6150 5704
rect 8680 5692 8708 5723
rect 9122 5720 9128 5772
rect 9180 5720 9186 5772
rect 9309 5763 9367 5769
rect 9309 5729 9321 5763
rect 9355 5729 9367 5763
rect 9309 5723 9367 5729
rect 9324 5692 9352 5723
rect 9398 5720 9404 5772
rect 9456 5720 9462 5772
rect 9508 5769 9536 5800
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5760 11207 5763
rect 11247 5760 11275 5868
rect 11698 5856 11704 5868
rect 11756 5896 11762 5908
rect 12434 5896 12440 5908
rect 11756 5868 12440 5896
rect 11756 5856 11762 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 12526 5856 12532 5908
rect 12584 5896 12590 5908
rect 13906 5896 13912 5908
rect 12584 5868 13912 5896
rect 12584 5856 12590 5868
rect 13906 5856 13912 5868
rect 13964 5896 13970 5908
rect 14274 5896 14280 5908
rect 13964 5868 14280 5896
rect 13964 5856 13970 5868
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 15010 5896 15016 5908
rect 14669 5868 15016 5896
rect 12158 5788 12164 5840
rect 12216 5828 12222 5840
rect 12253 5831 12311 5837
rect 12253 5828 12265 5831
rect 12216 5800 12265 5828
rect 12216 5788 12222 5800
rect 12253 5797 12265 5800
rect 12299 5797 12311 5831
rect 12253 5791 12311 5797
rect 13256 5831 13314 5837
rect 13256 5797 13268 5831
rect 13302 5828 13314 5831
rect 14182 5828 14188 5840
rect 13302 5800 14188 5828
rect 13302 5797 13314 5800
rect 13256 5791 13314 5797
rect 14182 5788 14188 5800
rect 14240 5788 14246 5840
rect 11195 5732 11275 5760
rect 11195 5729 11207 5732
rect 11149 5723 11207 5729
rect 11330 5720 11336 5772
rect 11388 5720 11394 5772
rect 11514 5720 11520 5772
rect 11572 5720 11578 5772
rect 11701 5763 11759 5769
rect 11701 5729 11713 5763
rect 11747 5729 11759 5763
rect 11701 5723 11759 5729
rect 8680 5664 9352 5692
rect 4709 5627 4767 5633
rect 4709 5624 4721 5627
rect 4080 5596 4721 5624
rect 4080 5568 4108 5596
rect 4709 5593 4721 5596
rect 4755 5593 4767 5627
rect 4709 5587 4767 5593
rect 9324 5568 9352 5664
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11348 5692 11376 5720
rect 11716 5692 11744 5723
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12437 5763 12495 5769
rect 12437 5760 12449 5763
rect 12032 5732 12449 5760
rect 12032 5720 12038 5732
rect 12437 5729 12449 5732
rect 12483 5729 12495 5763
rect 12437 5723 12495 5729
rect 14274 5720 14280 5772
rect 14332 5760 14338 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 14332 5732 14565 5760
rect 14332 5720 14338 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14669 5760 14697 5868
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 15562 5896 15568 5908
rect 15151 5868 15568 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 15654 5856 15660 5908
rect 15712 5856 15718 5908
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 15804 5868 16681 5896
rect 15804 5856 15810 5868
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 16669 5859 16727 5865
rect 17037 5899 17095 5905
rect 17037 5865 17049 5899
rect 17083 5896 17095 5899
rect 17494 5896 17500 5908
rect 17083 5868 17500 5896
rect 17083 5865 17095 5868
rect 17037 5859 17095 5865
rect 17494 5856 17500 5868
rect 17552 5856 17558 5908
rect 17770 5856 17776 5908
rect 17828 5896 17834 5908
rect 17865 5899 17923 5905
rect 17865 5896 17877 5899
rect 17828 5868 17877 5896
rect 17828 5856 17834 5868
rect 17865 5865 17877 5868
rect 17911 5865 17923 5899
rect 17865 5859 17923 5865
rect 18141 5899 18199 5905
rect 18141 5865 18153 5899
rect 18187 5896 18199 5899
rect 18322 5896 18328 5908
rect 18187 5868 18328 5896
rect 18187 5865 18199 5868
rect 18141 5859 18199 5865
rect 14734 5788 14740 5840
rect 14792 5828 14798 5840
rect 15286 5828 15292 5840
rect 14792 5800 15292 5828
rect 14792 5788 14798 5800
rect 15286 5788 15292 5800
rect 15344 5828 15350 5840
rect 15672 5828 15700 5856
rect 15344 5800 15608 5828
rect 15672 5800 17172 5828
rect 15344 5788 15350 5800
rect 14829 5763 14887 5769
rect 14829 5760 14841 5763
rect 14669 5732 14841 5760
rect 14553 5723 14611 5729
rect 14829 5729 14841 5732
rect 14875 5729 14887 5763
rect 14829 5723 14887 5729
rect 14921 5763 14979 5769
rect 14921 5729 14933 5763
rect 14967 5760 14979 5763
rect 15102 5760 15108 5772
rect 14967 5732 15108 5760
rect 14967 5729 14979 5732
rect 14921 5723 14979 5729
rect 15102 5720 15108 5732
rect 15160 5760 15166 5772
rect 15580 5769 15608 5800
rect 15381 5763 15439 5769
rect 15381 5760 15393 5763
rect 15160 5732 15393 5760
rect 15160 5720 15166 5732
rect 15381 5729 15393 5732
rect 15427 5729 15439 5763
rect 15381 5723 15439 5729
rect 15473 5763 15531 5769
rect 15473 5729 15485 5763
rect 15519 5729 15531 5763
rect 15473 5723 15531 5729
rect 15565 5763 15623 5769
rect 15565 5729 15577 5763
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 11112 5664 11376 5692
rect 11648 5664 11744 5692
rect 11112 5652 11118 5664
rect 9674 5584 9680 5636
rect 9732 5584 9738 5636
rect 10594 5584 10600 5636
rect 10652 5624 10658 5636
rect 10962 5624 10968 5636
rect 10652 5596 10968 5624
rect 10652 5584 10658 5596
rect 10962 5584 10968 5596
rect 11020 5584 11026 5636
rect 3510 5556 3516 5568
rect 3068 5528 3516 5556
rect 3510 5516 3516 5528
rect 3568 5556 3574 5568
rect 4062 5556 4068 5568
rect 3568 5528 4068 5556
rect 3568 5516 3574 5528
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4525 5559 4583 5565
rect 4525 5525 4537 5559
rect 4571 5556 4583 5559
rect 7926 5556 7932 5568
rect 4571 5528 7932 5556
rect 4571 5525 4583 5528
rect 4525 5519 4583 5525
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 9030 5516 9036 5568
rect 9088 5516 9094 5568
rect 9306 5516 9312 5568
rect 9364 5516 9370 5568
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 10502 5556 10508 5568
rect 9456 5528 10508 5556
rect 9456 5516 9462 5528
rect 10502 5516 10508 5528
rect 10560 5516 10566 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 11648 5556 11676 5664
rect 12986 5652 12992 5704
rect 13044 5652 13050 5704
rect 15488 5692 15516 5723
rect 15654 5720 15660 5772
rect 15712 5760 15718 5772
rect 15749 5763 15807 5769
rect 15749 5760 15761 5763
rect 15712 5732 15761 5760
rect 15712 5720 15718 5732
rect 15749 5729 15761 5732
rect 15795 5729 15807 5763
rect 15749 5723 15807 5729
rect 16298 5720 16304 5772
rect 16356 5720 16362 5772
rect 16482 5720 16488 5772
rect 16540 5720 16546 5772
rect 16592 5769 16620 5800
rect 17144 5769 17172 5800
rect 17218 5788 17224 5840
rect 17276 5828 17282 5840
rect 17313 5831 17371 5837
rect 17313 5828 17325 5831
rect 17276 5800 17325 5828
rect 17276 5788 17282 5800
rect 17313 5797 17325 5800
rect 17359 5828 17371 5831
rect 17589 5831 17647 5837
rect 17589 5828 17601 5831
rect 17359 5800 17601 5828
rect 17359 5797 17371 5800
rect 17313 5791 17371 5797
rect 17589 5797 17601 5800
rect 17635 5797 17647 5831
rect 18156 5828 18184 5859
rect 18322 5856 18328 5868
rect 18380 5896 18386 5908
rect 18417 5899 18475 5905
rect 18417 5896 18429 5899
rect 18380 5868 18429 5896
rect 18380 5856 18386 5868
rect 18417 5865 18429 5868
rect 18463 5865 18475 5899
rect 18417 5859 18475 5865
rect 17589 5791 17647 5797
rect 17696 5800 18184 5828
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5729 16635 5763
rect 16577 5723 16635 5729
rect 16853 5763 16911 5769
rect 16853 5729 16865 5763
rect 16899 5729 16911 5763
rect 16853 5723 16911 5729
rect 17129 5763 17187 5769
rect 17129 5729 17141 5763
rect 17175 5729 17187 5763
rect 17129 5723 17187 5729
rect 14384 5664 15516 5692
rect 16316 5692 16344 5720
rect 16868 5692 16896 5723
rect 17402 5720 17408 5772
rect 17460 5720 17466 5772
rect 17696 5769 17724 5800
rect 17681 5763 17739 5769
rect 17681 5729 17693 5763
rect 17727 5729 17739 5763
rect 17681 5723 17739 5729
rect 17957 5763 18015 5769
rect 17957 5729 17969 5763
rect 18003 5760 18015 5763
rect 18138 5760 18144 5772
rect 18003 5732 18144 5760
rect 18003 5729 18015 5732
rect 17957 5723 18015 5729
rect 18138 5720 18144 5732
rect 18196 5720 18202 5772
rect 18233 5763 18291 5769
rect 18233 5729 18245 5763
rect 18279 5760 18291 5763
rect 18322 5760 18328 5772
rect 18279 5732 18328 5760
rect 18279 5729 18291 5732
rect 18233 5723 18291 5729
rect 18322 5720 18328 5732
rect 18380 5720 18386 5772
rect 18506 5720 18512 5772
rect 18564 5720 18570 5772
rect 16316 5664 16896 5692
rect 11790 5584 11796 5636
rect 11848 5624 11854 5636
rect 14384 5633 14412 5664
rect 11977 5627 12035 5633
rect 11977 5624 11989 5627
rect 11848 5596 11989 5624
rect 11848 5584 11854 5596
rect 11977 5593 11989 5596
rect 12023 5593 12035 5627
rect 11977 5587 12035 5593
rect 14369 5627 14427 5633
rect 14369 5593 14381 5627
rect 14415 5593 14427 5627
rect 14369 5587 14427 5593
rect 10744 5528 11676 5556
rect 15197 5559 15255 5565
rect 10744 5516 10750 5528
rect 15197 5525 15209 5559
rect 15243 5556 15255 5559
rect 15378 5556 15384 5568
rect 15243 5528 15384 5556
rect 15243 5525 15255 5528
rect 15197 5519 15255 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 16114 5516 16120 5568
rect 16172 5516 16178 5568
rect 552 5466 19412 5488
rect 552 5414 2755 5466
rect 2807 5414 2819 5466
rect 2871 5414 2883 5466
rect 2935 5414 2947 5466
rect 2999 5414 3011 5466
rect 3063 5414 7470 5466
rect 7522 5414 7534 5466
rect 7586 5414 7598 5466
rect 7650 5414 7662 5466
rect 7714 5414 7726 5466
rect 7778 5414 12185 5466
rect 12237 5414 12249 5466
rect 12301 5414 12313 5466
rect 12365 5414 12377 5466
rect 12429 5414 12441 5466
rect 12493 5414 16900 5466
rect 16952 5414 16964 5466
rect 17016 5414 17028 5466
rect 17080 5414 17092 5466
rect 17144 5414 17156 5466
rect 17208 5414 19412 5466
rect 552 5392 19412 5414
rect 1397 5355 1455 5361
rect 1397 5321 1409 5355
rect 1443 5352 1455 5355
rect 1486 5352 1492 5364
rect 1443 5324 1492 5352
rect 1443 5321 1455 5324
rect 1397 5315 1455 5321
rect 1486 5312 1492 5324
rect 1544 5352 1550 5364
rect 1854 5352 1860 5364
rect 1544 5324 1860 5352
rect 1544 5312 1550 5324
rect 1854 5312 1860 5324
rect 1912 5312 1918 5364
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5321 3111 5355
rect 3053 5315 3111 5321
rect 6549 5355 6607 5361
rect 6549 5321 6561 5355
rect 6595 5352 6607 5355
rect 7834 5352 7840 5364
rect 6595 5324 7840 5352
rect 6595 5321 6607 5324
rect 6549 5315 6607 5321
rect 3068 5228 3096 5315
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 7926 5312 7932 5364
rect 7984 5352 7990 5364
rect 9398 5352 9404 5364
rect 7984 5324 9404 5352
rect 7984 5312 7990 5324
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 9490 5312 9496 5364
rect 9548 5312 9554 5364
rect 10778 5352 10784 5364
rect 9646 5324 10784 5352
rect 6730 5244 6736 5296
rect 6788 5284 6794 5296
rect 9646 5284 9674 5324
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 10965 5355 11023 5361
rect 10965 5352 10977 5355
rect 10928 5324 10977 5352
rect 10928 5312 10934 5324
rect 10965 5321 10977 5324
rect 11011 5321 11023 5355
rect 10965 5315 11023 5321
rect 11072 5324 13288 5352
rect 6788 5256 9674 5284
rect 6788 5244 6794 5256
rect 9858 5244 9864 5296
rect 9916 5284 9922 5296
rect 10594 5284 10600 5296
rect 9916 5256 10600 5284
rect 9916 5244 9922 5256
rect 10594 5244 10600 5256
rect 10652 5284 10658 5296
rect 11072 5284 11100 5324
rect 10652 5256 11100 5284
rect 10652 5244 10658 5256
rect 11330 5244 11336 5296
rect 11388 5284 11394 5296
rect 11974 5284 11980 5296
rect 11388 5256 11980 5284
rect 11388 5244 11394 5256
rect 11974 5244 11980 5256
rect 12032 5244 12038 5296
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 13260 5284 13288 5324
rect 13354 5312 13360 5364
rect 13412 5352 13418 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 13412 5324 13553 5352
rect 13412 5312 13418 5324
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 13541 5315 13599 5321
rect 14090 5312 14096 5364
rect 14148 5312 14154 5364
rect 14366 5312 14372 5364
rect 14424 5312 14430 5364
rect 14458 5312 14464 5364
rect 14516 5352 14522 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 14516 5324 15301 5352
rect 14516 5312 14522 5324
rect 15289 5321 15301 5324
rect 15335 5321 15347 5355
rect 15289 5315 15347 5321
rect 13814 5284 13820 5296
rect 12124 5256 13216 5284
rect 13260 5256 13820 5284
rect 12124 5244 12130 5256
rect 1121 5219 1179 5225
rect 1121 5185 1133 5219
rect 1167 5216 1179 5219
rect 1394 5216 1400 5228
rect 1167 5188 1400 5216
rect 1167 5185 1179 5188
rect 1121 5179 1179 5185
rect 1394 5176 1400 5188
rect 1452 5176 1458 5228
rect 3050 5176 3056 5228
rect 3108 5176 3114 5228
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 12084 5216 12112 5244
rect 8076 5188 12112 5216
rect 8076 5176 8082 5188
rect 1210 5108 1216 5160
rect 1268 5108 1274 5160
rect 1302 5108 1308 5160
rect 1360 5108 1366 5160
rect 1673 5151 1731 5157
rect 1673 5148 1685 5151
rect 1596 5120 1685 5148
rect 1596 5024 1624 5120
rect 1673 5117 1685 5120
rect 1719 5148 1731 5151
rect 3697 5151 3755 5157
rect 3697 5148 3709 5151
rect 1719 5120 3709 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 3697 5117 3709 5120
rect 3743 5148 3755 5151
rect 4246 5148 4252 5160
rect 3743 5120 4252 5148
rect 3743 5117 3755 5120
rect 3697 5111 3755 5117
rect 4246 5108 4252 5120
rect 4304 5148 4310 5160
rect 4982 5148 4988 5160
rect 4304 5120 4988 5148
rect 4304 5108 4310 5120
rect 4982 5108 4988 5120
rect 5040 5148 5046 5160
rect 5442 5157 5448 5160
rect 5169 5151 5227 5157
rect 5169 5148 5181 5151
rect 5040 5120 5181 5148
rect 5040 5108 5046 5120
rect 5169 5117 5181 5120
rect 5215 5117 5227 5151
rect 5169 5111 5227 5117
rect 5436 5111 5448 5157
rect 5442 5108 5448 5111
rect 5500 5108 5506 5160
rect 9324 5157 9352 5188
rect 9309 5151 9367 5157
rect 6472 5120 9168 5148
rect 1946 5089 1952 5092
rect 1940 5080 1952 5089
rect 1907 5052 1952 5080
rect 1940 5043 1952 5052
rect 1946 5040 1952 5043
rect 2004 5040 2010 5092
rect 3964 5083 4022 5089
rect 3964 5049 3976 5083
rect 4010 5080 4022 5083
rect 4062 5080 4068 5092
rect 4010 5052 4068 5080
rect 4010 5049 4022 5052
rect 3964 5043 4022 5049
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 1578 4972 1584 5024
rect 1636 4972 1642 5024
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 6472 5012 6500 5120
rect 8573 5083 8631 5089
rect 8573 5049 8585 5083
rect 8619 5080 8631 5083
rect 9030 5080 9036 5092
rect 8619 5052 9036 5080
rect 8619 5049 8631 5052
rect 8573 5043 8631 5049
rect 9030 5040 9036 5052
rect 9088 5040 9094 5092
rect 9140 5080 9168 5120
rect 9309 5117 9321 5151
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10045 5151 10103 5157
rect 9732 5120 9996 5148
rect 9732 5108 9738 5120
rect 9769 5083 9827 5089
rect 9769 5080 9781 5083
rect 9140 5052 9781 5080
rect 9769 5049 9781 5052
rect 9815 5049 9827 5083
rect 9769 5043 9827 5049
rect 9858 5040 9864 5092
rect 9916 5040 9922 5092
rect 5123 4984 6500 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 9876 5012 9904 5040
rect 9640 4984 9904 5012
rect 9968 5012 9996 5120
rect 10045 5117 10057 5151
rect 10091 5148 10103 5151
rect 10226 5148 10232 5160
rect 10091 5120 10232 5148
rect 10091 5117 10103 5120
rect 10045 5111 10103 5117
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 10410 5108 10416 5160
rect 10468 5108 10474 5160
rect 10502 5108 10508 5160
rect 10560 5148 10566 5160
rect 10689 5151 10747 5157
rect 10689 5148 10701 5151
rect 10560 5120 10701 5148
rect 10560 5108 10566 5120
rect 10689 5117 10701 5120
rect 10735 5117 10747 5151
rect 10689 5111 10747 5117
rect 10781 5151 10839 5157
rect 10781 5117 10793 5151
rect 10827 5117 10839 5151
rect 10781 5111 10839 5117
rect 10594 5040 10600 5092
rect 10652 5040 10658 5092
rect 10686 5012 10692 5024
rect 9968 4984 10692 5012
rect 9640 4972 9646 4984
rect 10686 4972 10692 4984
rect 10744 5012 10750 5024
rect 10796 5012 10824 5111
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 11425 5151 11483 5157
rect 11425 5148 11437 5151
rect 11112 5120 11437 5148
rect 11112 5108 11118 5120
rect 11425 5117 11437 5120
rect 11471 5117 11483 5151
rect 11425 5111 11483 5117
rect 11517 5151 11575 5157
rect 11517 5117 11529 5151
rect 11563 5148 11575 5151
rect 11698 5148 11704 5160
rect 11563 5120 11704 5148
rect 11563 5117 11575 5120
rect 11517 5111 11575 5117
rect 11698 5108 11704 5120
rect 11756 5108 11762 5160
rect 11977 5151 12035 5157
rect 11977 5148 11989 5151
rect 11808 5120 11989 5148
rect 11808 5092 11836 5120
rect 11977 5117 11989 5120
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 12066 5108 12072 5160
rect 12124 5148 12130 5160
rect 13188 5148 13216 5256
rect 13814 5244 13820 5256
rect 13872 5244 13878 5296
rect 14384 5284 14412 5312
rect 15105 5287 15163 5293
rect 15105 5284 15117 5287
rect 14384 5256 15117 5284
rect 15105 5253 15117 5256
rect 15151 5253 15163 5287
rect 15105 5247 15163 5253
rect 15194 5216 15200 5228
rect 13372 5188 15200 5216
rect 13372 5157 13400 5188
rect 15194 5176 15200 5188
rect 15252 5176 15258 5228
rect 15473 5219 15531 5225
rect 15473 5185 15485 5219
rect 15519 5216 15531 5219
rect 16114 5216 16120 5228
rect 15519 5188 16120 5216
rect 15519 5185 15531 5188
rect 15473 5179 15531 5185
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 13357 5151 13415 5157
rect 13357 5148 13369 5151
rect 12124 5120 13124 5148
rect 13188 5120 13369 5148
rect 12124 5108 12130 5120
rect 11238 5040 11244 5092
rect 11296 5080 11302 5092
rect 11333 5083 11391 5089
rect 11333 5080 11345 5083
rect 11296 5052 11345 5080
rect 11296 5040 11302 5052
rect 11333 5049 11345 5052
rect 11379 5049 11391 5083
rect 11333 5043 11391 5049
rect 10744 4984 10824 5012
rect 11348 5012 11376 5043
rect 11790 5040 11796 5092
rect 11848 5040 11854 5092
rect 11885 5083 11943 5089
rect 11885 5049 11897 5083
rect 11931 5080 11943 5083
rect 12434 5080 12440 5092
rect 11931 5052 12440 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 12434 5040 12440 5052
rect 12492 5040 12498 5092
rect 12526 5040 12532 5092
rect 12584 5040 12590 5092
rect 12894 5040 12900 5092
rect 12952 5040 12958 5092
rect 13096 5080 13124 5120
rect 13357 5117 13369 5120
rect 13403 5117 13415 5151
rect 13357 5111 13415 5117
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5117 13783 5151
rect 13725 5111 13783 5117
rect 13740 5080 13768 5111
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 13872 5120 14013 5148
rect 13872 5108 13878 5120
rect 14001 5117 14013 5120
rect 14047 5117 14059 5151
rect 14001 5111 14059 5117
rect 14277 5151 14335 5157
rect 14277 5117 14289 5151
rect 14323 5117 14335 5151
rect 14277 5111 14335 5117
rect 14292 5080 14320 5111
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14424 5120 14565 5148
rect 14424 5108 14430 5120
rect 14553 5117 14565 5120
rect 14599 5148 14611 5151
rect 14734 5148 14740 5160
rect 14599 5120 14740 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 14734 5108 14740 5120
rect 14792 5108 14798 5160
rect 15286 5108 15292 5160
rect 15344 5108 15350 5160
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 15436 5120 15577 5148
rect 15436 5108 15442 5120
rect 15565 5117 15577 5120
rect 15611 5117 15623 5151
rect 15565 5111 15623 5117
rect 18046 5108 18052 5160
rect 18104 5148 18110 5160
rect 18141 5151 18199 5157
rect 18141 5148 18153 5151
rect 18104 5120 18153 5148
rect 18104 5108 18110 5120
rect 18141 5117 18153 5120
rect 18187 5117 18199 5151
rect 18141 5111 18199 5117
rect 18233 5151 18291 5157
rect 18233 5117 18245 5151
rect 18279 5117 18291 5151
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18233 5111 18291 5117
rect 18340 5120 18705 5148
rect 16298 5080 16304 5092
rect 13096 5052 16304 5080
rect 16298 5040 16304 5052
rect 16356 5040 16362 5092
rect 17402 5040 17408 5092
rect 17460 5080 17466 5092
rect 17874 5083 17932 5089
rect 17874 5080 17886 5083
rect 17460 5052 17886 5080
rect 17460 5040 17466 5052
rect 17874 5049 17886 5052
rect 17920 5080 17932 5083
rect 18248 5080 18276 5111
rect 17920 5052 18276 5080
rect 17920 5049 17932 5052
rect 17874 5043 17932 5049
rect 12912 5012 12940 5040
rect 11348 4984 12940 5012
rect 10744 4972 10750 4984
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 13909 5015 13967 5021
rect 13909 5012 13921 5015
rect 13872 4984 13921 5012
rect 13872 4972 13878 4984
rect 13909 4981 13921 4984
rect 13955 4981 13967 5015
rect 13909 4975 13967 4981
rect 14458 4972 14464 5024
rect 14516 4972 14522 5024
rect 16758 4972 16764 5024
rect 16816 4972 16822 5024
rect 18138 4972 18144 5024
rect 18196 5012 18202 5024
rect 18340 5021 18368 5120
rect 18693 5117 18705 5120
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 18325 5015 18383 5021
rect 18325 5012 18337 5015
rect 18196 4984 18337 5012
rect 18196 4972 18202 4984
rect 18325 4981 18337 4984
rect 18371 4981 18383 5015
rect 18325 4975 18383 4981
rect 18782 4972 18788 5024
rect 18840 4972 18846 5024
rect 552 4922 19571 4944
rect 552 4870 5112 4922
rect 5164 4870 5176 4922
rect 5228 4870 5240 4922
rect 5292 4870 5304 4922
rect 5356 4870 5368 4922
rect 5420 4870 9827 4922
rect 9879 4870 9891 4922
rect 9943 4870 9955 4922
rect 10007 4870 10019 4922
rect 10071 4870 10083 4922
rect 10135 4870 14542 4922
rect 14594 4870 14606 4922
rect 14658 4870 14670 4922
rect 14722 4870 14734 4922
rect 14786 4870 14798 4922
rect 14850 4870 19257 4922
rect 19309 4870 19321 4922
rect 19373 4870 19385 4922
rect 19437 4870 19449 4922
rect 19501 4870 19513 4922
rect 19565 4870 19571 4922
rect 552 4848 19571 4870
rect 1302 4768 1308 4820
rect 1360 4768 1366 4820
rect 1397 4811 1455 4817
rect 1397 4777 1409 4811
rect 1443 4808 1455 4811
rect 1670 4808 1676 4820
rect 1443 4780 1676 4808
rect 1443 4777 1455 4780
rect 1397 4771 1455 4777
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 2961 4811 3019 4817
rect 2961 4777 2973 4811
rect 3007 4777 3019 4811
rect 2961 4771 3019 4777
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5810 4808 5816 4820
rect 5307 4780 5816 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 1213 4675 1271 4681
rect 1213 4641 1225 4675
rect 1259 4672 1271 4675
rect 1320 4672 1348 4768
rect 1826 4743 1884 4749
rect 1826 4740 1838 4743
rect 1412 4712 1838 4740
rect 1412 4684 1440 4712
rect 1826 4709 1838 4712
rect 1872 4709 1884 4743
rect 2976 4740 3004 4771
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 7469 4811 7527 4817
rect 7469 4777 7481 4811
rect 7515 4808 7527 4811
rect 8478 4808 8484 4820
rect 7515 4780 8484 4808
rect 7515 4777 7527 4780
rect 7469 4771 7527 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 9401 4811 9459 4817
rect 9401 4777 9413 4811
rect 9447 4808 9459 4811
rect 10410 4808 10416 4820
rect 9447 4780 10416 4808
rect 9447 4777 9459 4780
rect 9401 4771 9459 4777
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 10962 4768 10968 4820
rect 11020 4808 11026 4820
rect 12161 4811 12219 4817
rect 12161 4808 12173 4811
rect 11020 4780 12173 4808
rect 11020 4768 11026 4780
rect 12161 4777 12173 4780
rect 12207 4777 12219 4811
rect 12161 4771 12219 4777
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 14366 4808 14372 4820
rect 12400 4780 14372 4808
rect 12400 4768 12406 4780
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 15933 4811 15991 4817
rect 15933 4777 15945 4811
rect 15979 4808 15991 4811
rect 16022 4808 16028 4820
rect 15979 4780 16028 4808
rect 15979 4777 15991 4780
rect 15933 4771 15991 4777
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 16758 4768 16764 4820
rect 16816 4768 16822 4820
rect 17681 4811 17739 4817
rect 17681 4808 17693 4811
rect 16887 4780 17693 4808
rect 9064 4743 9122 4749
rect 2976 4712 7328 4740
rect 1826 4703 1884 4709
rect 1259 4644 1348 4672
rect 1259 4641 1271 4644
rect 1213 4635 1271 4641
rect 1394 4632 1400 4684
rect 1452 4632 1458 4684
rect 1486 4632 1492 4684
rect 1544 4632 1550 4684
rect 4148 4675 4206 4681
rect 4148 4641 4160 4675
rect 4194 4672 4206 4675
rect 4430 4672 4436 4684
rect 4194 4644 4436 4672
rect 4194 4641 4206 4644
rect 4148 4635 4206 4641
rect 4430 4632 4436 4644
rect 4488 4632 4494 4684
rect 6362 4681 6368 4684
rect 6356 4635 6368 4681
rect 6362 4632 6368 4635
rect 6420 4632 6426 4684
rect 7300 4672 7328 4712
rect 9064 4709 9076 4743
rect 9110 4740 9122 4743
rect 10686 4740 10692 4752
rect 9110 4712 10692 4740
rect 9110 4709 9122 4712
rect 9064 4703 9122 4709
rect 10686 4700 10692 4712
rect 10744 4700 10750 4752
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 11793 4743 11851 4749
rect 11793 4740 11805 4743
rect 11388 4712 11805 4740
rect 11388 4700 11394 4712
rect 11793 4709 11805 4712
rect 11839 4709 11851 4743
rect 11793 4703 11851 4709
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 12437 4743 12495 4749
rect 12437 4740 12449 4743
rect 12124 4712 12449 4740
rect 12124 4700 12130 4712
rect 12437 4709 12449 4712
rect 12483 4709 12495 4743
rect 12437 4703 12495 4709
rect 12529 4743 12587 4749
rect 12529 4709 12541 4743
rect 12575 4740 12587 4743
rect 12618 4740 12624 4752
rect 12575 4712 12624 4740
rect 12575 4709 12587 4712
rect 12529 4703 12587 4709
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 16776 4740 16804 4768
rect 13832 4712 16804 4740
rect 7300 4644 9674 4672
rect 1578 4564 1584 4616
rect 1636 4564 1642 4616
rect 3881 4607 3939 4613
rect 3881 4604 3893 4607
rect 2746 4576 3893 4604
rect 1118 4428 1124 4480
rect 1176 4428 1182 4480
rect 1596 4468 1624 4564
rect 2590 4468 2596 4480
rect 1596 4440 2596 4468
rect 2590 4428 2596 4440
rect 2648 4468 2654 4480
rect 2746 4468 2774 4576
rect 3881 4573 3893 4576
rect 3927 4573 3939 4607
rect 3881 4567 3939 4573
rect 6086 4564 6092 4616
rect 6144 4564 6150 4616
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 2648 4440 2774 4468
rect 7929 4471 7987 4477
rect 2648 4428 2654 4440
rect 7929 4437 7941 4471
rect 7975 4468 7987 4471
rect 8386 4468 8392 4480
rect 7975 4440 8392 4468
rect 7975 4437 7987 4440
rect 7929 4431 7987 4437
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 9030 4428 9036 4480
rect 9088 4468 9094 4480
rect 9324 4468 9352 4567
rect 9088 4440 9352 4468
rect 9646 4468 9674 4644
rect 10502 4632 10508 4684
rect 10560 4681 10566 4684
rect 10560 4635 10572 4681
rect 10560 4632 10566 4635
rect 10962 4632 10968 4684
rect 11020 4632 11026 4684
rect 11054 4632 11060 4684
rect 11112 4632 11118 4684
rect 11238 4632 11244 4684
rect 11296 4632 11302 4684
rect 11422 4632 11428 4684
rect 11480 4632 11486 4684
rect 11517 4675 11575 4681
rect 11517 4641 11529 4675
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 10778 4564 10784 4616
rect 10836 4564 10842 4616
rect 11532 4468 11560 4635
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11664 4644 11713 4672
rect 11664 4632 11670 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 11701 4635 11759 4641
rect 11885 4675 11943 4681
rect 11885 4641 11897 4675
rect 11931 4672 11943 4675
rect 12342 4672 12348 4684
rect 11931 4644 12348 4672
rect 11931 4641 11943 4644
rect 11885 4635 11943 4641
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 12713 4675 12771 4681
rect 12713 4641 12725 4675
rect 12759 4672 12771 4675
rect 13832 4672 13860 4712
rect 12759 4644 13860 4672
rect 14820 4675 14878 4681
rect 12759 4641 12771 4644
rect 12713 4635 12771 4641
rect 14820 4641 14832 4675
rect 14866 4672 14878 4675
rect 15378 4672 15384 4684
rect 14866 4644 15384 4672
rect 14866 4641 14878 4644
rect 14820 4635 14878 4641
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 16482 4632 16488 4684
rect 16540 4672 16546 4684
rect 16887 4672 16915 4780
rect 17681 4777 17693 4780
rect 17727 4777 17739 4811
rect 18506 4808 18512 4820
rect 17681 4771 17739 4777
rect 17926 4780 18512 4808
rect 17037 4743 17095 4749
rect 17037 4709 17049 4743
rect 17083 4740 17095 4743
rect 17402 4740 17408 4752
rect 17083 4712 17408 4740
rect 17083 4709 17095 4712
rect 17037 4703 17095 4709
rect 17402 4700 17408 4712
rect 17460 4700 17466 4752
rect 16540 4644 16915 4672
rect 16945 4675 17003 4681
rect 16540 4632 16546 4644
rect 16945 4641 16957 4675
rect 16991 4641 17003 4675
rect 16945 4635 17003 4641
rect 17497 4675 17555 4681
rect 17497 4641 17509 4675
rect 17543 4672 17555 4675
rect 17926 4672 17954 4780
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 18966 4740 18972 4752
rect 18064 4712 18972 4740
rect 18064 4684 18092 4712
rect 18966 4700 18972 4712
rect 19024 4740 19030 4752
rect 19024 4712 19104 4740
rect 19024 4700 19030 4712
rect 17543 4644 17954 4672
rect 17543 4641 17555 4644
rect 17497 4635 17555 4641
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 13044 4576 14565 4604
rect 13044 4564 13050 4576
rect 14553 4573 14565 4576
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 12069 4539 12127 4545
rect 12069 4505 12081 4539
rect 12115 4536 12127 4539
rect 13078 4536 13084 4548
rect 12115 4508 13084 4536
rect 12115 4505 12127 4508
rect 12069 4499 12127 4505
rect 13078 4496 13084 4508
rect 13136 4496 13142 4548
rect 9646 4440 11560 4468
rect 9088 4428 9094 4440
rect 11606 4428 11612 4480
rect 11664 4468 11670 4480
rect 16758 4468 16764 4480
rect 11664 4440 16764 4468
rect 11664 4428 11670 4440
rect 16758 4428 16764 4440
rect 16816 4468 16822 4480
rect 16960 4468 16988 4635
rect 18046 4632 18052 4684
rect 18104 4632 18110 4684
rect 18322 4632 18328 4684
rect 18380 4672 18386 4684
rect 18782 4672 18788 4684
rect 18840 4681 18846 4684
rect 19076 4681 19104 4712
rect 18380 4644 18788 4672
rect 18380 4632 18386 4644
rect 18782 4632 18788 4644
rect 18840 4635 18852 4681
rect 19061 4675 19119 4681
rect 19061 4641 19073 4675
rect 19107 4641 19119 4675
rect 19061 4635 19119 4641
rect 18840 4632 18846 4635
rect 16816 4440 16988 4468
rect 16816 4428 16822 4440
rect 552 4378 19412 4400
rect 552 4326 2755 4378
rect 2807 4326 2819 4378
rect 2871 4326 2883 4378
rect 2935 4326 2947 4378
rect 2999 4326 3011 4378
rect 3063 4326 7470 4378
rect 7522 4326 7534 4378
rect 7586 4326 7598 4378
rect 7650 4326 7662 4378
rect 7714 4326 7726 4378
rect 7778 4326 12185 4378
rect 12237 4326 12249 4378
rect 12301 4326 12313 4378
rect 12365 4326 12377 4378
rect 12429 4326 12441 4378
rect 12493 4326 16900 4378
rect 16952 4326 16964 4378
rect 17016 4326 17028 4378
rect 17080 4326 17092 4378
rect 17144 4326 17156 4378
rect 17208 4326 19412 4378
rect 552 4304 19412 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 1489 4267 1547 4273
rect 1489 4264 1501 4267
rect 1452 4236 1501 4264
rect 1452 4224 1458 4236
rect 1489 4233 1501 4236
rect 1535 4233 1547 4267
rect 1489 4227 1547 4233
rect 10137 4267 10195 4273
rect 10137 4233 10149 4267
rect 10183 4264 10195 4267
rect 10226 4264 10232 4276
rect 10183 4236 10232 4264
rect 10183 4233 10195 4236
rect 10137 4227 10195 4233
rect 1118 4020 1124 4072
rect 1176 4020 1182 4072
rect 1394 4020 1400 4072
rect 1452 4020 1458 4072
rect 1504 4060 1532 4227
rect 10226 4224 10232 4236
rect 10284 4224 10290 4276
rect 10502 4224 10508 4276
rect 10560 4264 10566 4276
rect 10597 4267 10655 4273
rect 10597 4264 10609 4267
rect 10560 4236 10609 4264
rect 10560 4224 10566 4236
rect 10597 4233 10609 4236
rect 10643 4264 10655 4267
rect 11514 4264 11520 4276
rect 10643 4236 11520 4264
rect 10643 4233 10655 4236
rect 10597 4227 10655 4233
rect 11514 4224 11520 4236
rect 11572 4224 11578 4276
rect 12526 4264 12532 4276
rect 11624 4236 12532 4264
rect 1946 4156 1952 4208
rect 2004 4156 2010 4208
rect 1670 4060 1676 4072
rect 1504 4032 1676 4060
rect 1670 4020 1676 4032
rect 1728 4020 1734 4072
rect 1964 4069 1992 4156
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5077 4131 5135 4137
rect 5077 4128 5089 4131
rect 5040 4100 5089 4128
rect 5040 4088 5046 4100
rect 5077 4097 5089 4100
rect 5123 4097 5135 4131
rect 5077 4091 5135 4097
rect 6822 4088 6828 4140
rect 6880 4088 6886 4140
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4029 2007 4063
rect 1949 4023 2007 4029
rect 8757 4063 8815 4069
rect 8757 4029 8769 4063
rect 8803 4060 8815 4063
rect 9024 4063 9082 4069
rect 8803 4032 8892 4060
rect 8803 4029 8815 4032
rect 8757 4023 8815 4029
rect 1136 3992 1164 4020
rect 8864 4004 8892 4032
rect 9024 4029 9036 4063
rect 9070 4060 9082 4063
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 9070 4032 10517 4060
rect 9070 4029 9082 4032
rect 9024 4023 9082 4029
rect 10505 4029 10517 4032
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 1302 3992 1308 4004
rect 1136 3964 1308 3992
rect 1302 3952 1308 3964
rect 1360 3992 1366 4004
rect 1765 3995 1823 4001
rect 1765 3992 1777 3995
rect 1360 3964 1777 3992
rect 1360 3952 1366 3964
rect 1765 3961 1777 3964
rect 1811 3961 1823 3995
rect 1765 3955 1823 3961
rect 5344 3995 5402 4001
rect 5344 3961 5356 3995
rect 5390 3992 5402 3995
rect 5442 3992 5448 4004
rect 5390 3964 5448 3992
rect 5390 3961 5402 3964
rect 5344 3955 5402 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 7092 3995 7150 4001
rect 7092 3961 7104 3995
rect 7138 3992 7150 3995
rect 7282 3992 7288 4004
rect 7138 3964 7288 3992
rect 7138 3961 7150 3964
rect 7092 3955 7150 3961
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 8128 3964 8800 3992
rect 1118 3884 1124 3936
rect 1176 3924 1182 3936
rect 2038 3924 2044 3936
rect 1176 3896 2044 3924
rect 1176 3884 1182 3896
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 8128 3924 8156 3964
rect 6503 3896 8156 3924
rect 8205 3927 8263 3933
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 8205 3893 8217 3927
rect 8251 3924 8263 3927
rect 8662 3924 8668 3936
rect 8251 3896 8668 3924
rect 8251 3893 8263 3896
rect 8205 3887 8263 3893
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 8772 3924 8800 3964
rect 8846 3952 8852 4004
rect 8904 3952 8910 4004
rect 10520 3992 10548 4023
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 11624 4069 11652 4236
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 13541 4267 13599 4273
rect 13541 4233 13553 4267
rect 13587 4264 13599 4267
rect 13998 4264 14004 4276
rect 13587 4236 14004 4264
rect 13587 4233 13599 4236
rect 13541 4227 13599 4233
rect 13998 4224 14004 4236
rect 14056 4224 14062 4276
rect 15930 4224 15936 4276
rect 15988 4264 15994 4276
rect 17218 4264 17224 4276
rect 15988 4236 17224 4264
rect 15988 4224 15994 4236
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 18322 4224 18328 4276
rect 18380 4224 18386 4276
rect 18506 4224 18512 4276
rect 18564 4264 18570 4276
rect 18785 4267 18843 4273
rect 18785 4264 18797 4267
rect 18564 4236 18797 4264
rect 18564 4224 18570 4236
rect 18785 4233 18797 4236
rect 18831 4233 18843 4267
rect 18785 4227 18843 4233
rect 16758 4156 16764 4208
rect 16816 4196 16822 4208
rect 17773 4199 17831 4205
rect 17773 4196 17785 4199
rect 16816 4168 17785 4196
rect 16816 4156 16822 4168
rect 13740 4100 13952 4128
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 10836 4032 11621 4060
rect 10836 4020 10842 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 13740 4060 13768 4100
rect 11609 4023 11667 4029
rect 11716 4032 13768 4060
rect 11716 3992 11744 4032
rect 13814 4020 13820 4072
rect 13872 4020 13878 4072
rect 13924 4060 13952 4100
rect 15378 4088 15384 4140
rect 15436 4088 15442 4140
rect 15562 4088 15568 4140
rect 15620 4128 15626 4140
rect 16301 4131 16359 4137
rect 15620 4100 15792 4128
rect 15620 4088 15626 4100
rect 14921 4063 14979 4069
rect 13924 4032 14872 4060
rect 10520 3964 11744 3992
rect 11876 3995 11934 4001
rect 11876 3961 11888 3995
rect 11922 3992 11934 3995
rect 12802 3992 12808 4004
rect 11922 3964 12808 3992
rect 11922 3961 11934 3964
rect 11876 3955 11934 3961
rect 12802 3952 12808 3964
rect 12860 3952 12866 4004
rect 13832 3992 13860 4020
rect 13004 3964 13860 3992
rect 11054 3924 11060 3936
rect 8772 3896 11060 3924
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 13004 3933 13032 3964
rect 14366 3952 14372 4004
rect 14424 3992 14430 4004
rect 14654 3995 14712 4001
rect 14654 3992 14666 3995
rect 14424 3964 14666 3992
rect 14424 3952 14430 3964
rect 14654 3961 14666 3964
rect 14700 3961 14712 3995
rect 14844 3992 14872 4032
rect 14921 4029 14933 4063
rect 14967 4060 14979 4063
rect 15194 4060 15200 4072
rect 14967 4032 15200 4060
rect 14967 4029 14979 4032
rect 14921 4023 14979 4029
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 15396 4060 15424 4088
rect 15764 4069 15792 4100
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 16347 4100 16988 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 16960 4072 16988 4100
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 15396 4032 15485 4060
rect 15473 4029 15485 4032
rect 15519 4060 15531 4063
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 15519 4032 15669 4060
rect 15519 4029 15531 4032
rect 15473 4023 15531 4029
rect 15657 4029 15669 4032
rect 15703 4029 15715 4063
rect 15657 4023 15715 4029
rect 15749 4063 15807 4069
rect 15749 4029 15761 4063
rect 15795 4029 15807 4063
rect 15749 4023 15807 4029
rect 16114 4020 16120 4072
rect 16172 4020 16178 4072
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4029 16267 4063
rect 16209 4023 16267 4029
rect 16669 4063 16727 4069
rect 16669 4029 16681 4063
rect 16715 4029 16727 4063
rect 16669 4023 16727 4029
rect 15381 3995 15439 4001
rect 15381 3992 15393 3995
rect 14844 3964 15393 3992
rect 14654 3955 14712 3961
rect 15381 3961 15393 3964
rect 15427 3992 15439 3995
rect 16025 3995 16083 4001
rect 16025 3992 16037 3995
rect 15427 3964 16037 3992
rect 15427 3961 15439 3964
rect 15381 3955 15439 3961
rect 16025 3961 16037 3964
rect 16071 3992 16083 3995
rect 16224 3992 16252 4023
rect 16071 3964 16252 3992
rect 16684 3992 16712 4023
rect 16942 4020 16948 4072
rect 17000 4020 17006 4072
rect 17236 4069 17264 4168
rect 17773 4165 17785 4168
rect 17819 4165 17831 4199
rect 17773 4159 17831 4165
rect 18049 4131 18107 4137
rect 17328 4100 17908 4128
rect 17328 4072 17356 4100
rect 17221 4063 17279 4069
rect 17221 4029 17233 4063
rect 17267 4029 17279 4063
rect 17221 4023 17279 4029
rect 17310 4020 17316 4072
rect 17368 4020 17374 4072
rect 17880 4069 17908 4100
rect 18049 4097 18061 4131
rect 18095 4128 18107 4131
rect 18524 4128 18552 4224
rect 18095 4100 18552 4128
rect 18095 4097 18107 4100
rect 18049 4091 18107 4097
rect 17405 4063 17463 4069
rect 17405 4029 17417 4063
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4060 17923 4063
rect 17957 4063 18015 4069
rect 17957 4060 17969 4063
rect 17911 4032 17969 4060
rect 17911 4029 17923 4032
rect 17865 4023 17923 4029
rect 17957 4029 17969 4032
rect 18003 4029 18015 4063
rect 17957 4023 18015 4029
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4060 18475 4063
rect 18693 4063 18751 4069
rect 18693 4060 18705 4063
rect 18463 4032 18705 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 18693 4029 18705 4032
rect 18739 4029 18751 4063
rect 18693 4023 18751 4029
rect 16853 3995 16911 4001
rect 16853 3992 16865 3995
rect 16684 3964 16865 3992
rect 16071 3961 16083 3964
rect 16025 3955 16083 3961
rect 16853 3961 16865 3964
rect 16899 3992 16911 3995
rect 17129 3995 17187 4001
rect 17129 3992 17141 3995
rect 16899 3964 17141 3992
rect 16899 3961 16911 3964
rect 16853 3955 16911 3961
rect 17129 3961 17141 3964
rect 17175 3992 17187 3995
rect 17420 3992 17448 4023
rect 17175 3964 17448 3992
rect 17497 3995 17555 4001
rect 17175 3961 17187 3964
rect 17129 3955 17187 3961
rect 17497 3961 17509 3995
rect 17543 3992 17555 3995
rect 18138 3992 18144 4004
rect 17543 3964 18144 3992
rect 17543 3961 17555 3964
rect 17497 3955 17555 3961
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 12989 3927 13047 3933
rect 12989 3893 13001 3927
rect 13035 3893 13047 3927
rect 12989 3887 13047 3893
rect 16577 3927 16635 3933
rect 16577 3893 16589 3927
rect 16623 3924 16635 3927
rect 17862 3924 17868 3936
rect 16623 3896 17868 3924
rect 16623 3893 16635 3896
rect 16577 3887 16635 3893
rect 17862 3884 17868 3896
rect 17920 3924 17926 3936
rect 18432 3924 18460 4023
rect 17920 3896 18460 3924
rect 17920 3884 17926 3896
rect 552 3834 19571 3856
rect 552 3782 5112 3834
rect 5164 3782 5176 3834
rect 5228 3782 5240 3834
rect 5292 3782 5304 3834
rect 5356 3782 5368 3834
rect 5420 3782 9827 3834
rect 9879 3782 9891 3834
rect 9943 3782 9955 3834
rect 10007 3782 10019 3834
rect 10071 3782 10083 3834
rect 10135 3782 14542 3834
rect 14594 3782 14606 3834
rect 14658 3782 14670 3834
rect 14722 3782 14734 3834
rect 14786 3782 14798 3834
rect 14850 3782 19257 3834
rect 19309 3782 19321 3834
rect 19373 3782 19385 3834
rect 19437 3782 19449 3834
rect 19501 3782 19513 3834
rect 19565 3782 19571 3834
rect 552 3760 19571 3782
rect 1118 3680 1124 3732
rect 1176 3680 1182 3732
rect 1670 3680 1676 3732
rect 1728 3680 1734 3732
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 4985 3723 5043 3729
rect 4985 3720 4997 3723
rect 4948 3692 4997 3720
rect 4948 3680 4954 3692
rect 4985 3689 4997 3692
rect 5031 3689 5043 3723
rect 4985 3683 5043 3689
rect 5445 3723 5503 3729
rect 5445 3689 5457 3723
rect 5491 3720 5503 3723
rect 5626 3720 5632 3732
rect 5491 3692 5632 3720
rect 5491 3689 5503 3692
rect 5445 3683 5503 3689
rect 5626 3680 5632 3692
rect 5684 3720 5690 3732
rect 6362 3720 6368 3732
rect 5684 3692 6368 3720
rect 5684 3680 5690 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 8113 3723 8171 3729
rect 8113 3689 8125 3723
rect 8159 3720 8171 3723
rect 9122 3720 9128 3732
rect 8159 3692 9128 3720
rect 8159 3689 8171 3692
rect 8113 3683 8171 3689
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 10318 3680 10324 3732
rect 10376 3720 10382 3732
rect 10597 3723 10655 3729
rect 10597 3720 10609 3723
rect 10376 3692 10609 3720
rect 10376 3680 10382 3692
rect 10597 3689 10609 3692
rect 10643 3689 10655 3723
rect 10597 3683 10655 3689
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 14369 3723 14427 3729
rect 10744 3692 14320 3720
rect 10744 3680 10750 3692
rect 1213 3587 1271 3593
rect 1213 3553 1225 3587
rect 1259 3553 1271 3587
rect 1213 3547 1271 3553
rect 1228 3516 1256 3547
rect 1302 3544 1308 3596
rect 1360 3544 1366 3596
rect 1688 3584 1716 3680
rect 2590 3652 2596 3664
rect 1964 3624 2596 3652
rect 1765 3587 1823 3593
rect 1765 3584 1777 3587
rect 1688 3556 1777 3584
rect 1765 3553 1777 3556
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 1578 3516 1584 3528
rect 1228 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 1964 3525 1992 3624
rect 2590 3612 2596 3624
rect 2648 3652 2654 3664
rect 6380 3652 6408 3680
rect 2648 3624 2774 3652
rect 2648 3612 2654 3624
rect 2222 3593 2228 3596
rect 2216 3584 2228 3593
rect 2183 3556 2228 3584
rect 2216 3547 2228 3556
rect 2222 3544 2228 3547
rect 2280 3544 2286 3596
rect 2746 3584 2774 3624
rect 6288 3624 6408 3652
rect 14292 3652 14320 3692
rect 14369 3689 14381 3723
rect 14415 3720 14427 3723
rect 14458 3720 14464 3732
rect 14415 3692 14464 3720
rect 14415 3689 14427 3692
rect 14369 3683 14427 3689
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 14829 3723 14887 3729
rect 14829 3720 14841 3723
rect 14669 3692 14841 3720
rect 14669 3652 14697 3692
rect 14829 3689 14841 3692
rect 14875 3720 14887 3723
rect 15102 3720 15108 3732
rect 14875 3692 15108 3720
rect 14875 3689 14887 3692
rect 14829 3683 14887 3689
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 15436 3692 15485 3720
rect 15436 3680 15442 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 16209 3723 16267 3729
rect 16209 3720 16221 3723
rect 15473 3683 15531 3689
rect 15571 3692 16221 3720
rect 14292 3624 14697 3652
rect 3605 3587 3663 3593
rect 3605 3584 3617 3587
rect 2746 3556 3617 3584
rect 3605 3553 3617 3556
rect 3651 3553 3663 3587
rect 3605 3547 3663 3553
rect 3694 3544 3700 3596
rect 3752 3584 3758 3596
rect 3861 3587 3919 3593
rect 3861 3584 3873 3587
rect 3752 3556 3873 3584
rect 3752 3544 3758 3556
rect 3861 3553 3873 3556
rect 3907 3553 3919 3587
rect 5353 3587 5411 3593
rect 5353 3584 5365 3587
rect 3861 3547 3919 3553
rect 4632 3556 5365 3584
rect 1949 3519 2007 3525
rect 1949 3516 1961 3519
rect 1728 3488 1961 3516
rect 1728 3476 1734 3488
rect 1949 3485 1961 3488
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 4632 3460 4660 3556
rect 5353 3553 5365 3556
rect 5399 3584 5411 3587
rect 5442 3584 5448 3596
rect 5399 3556 5448 3584
rect 5399 3553 5411 3556
rect 5353 3547 5411 3553
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 6086 3544 6092 3596
rect 6144 3544 6150 3596
rect 6288 3593 6316 3624
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 6362 3544 6368 3596
rect 6420 3584 6426 3596
rect 6989 3587 7047 3593
rect 6989 3584 7001 3587
rect 6420 3556 7001 3584
rect 6420 3544 6426 3556
rect 6989 3553 7001 3556
rect 7035 3553 7047 3587
rect 6989 3547 7047 3553
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 9473 3587 9531 3593
rect 9473 3584 9485 3587
rect 8812 3556 9485 3584
rect 8812 3544 8818 3556
rect 9473 3553 9485 3556
rect 9519 3553 9531 3587
rect 9473 3547 9531 3553
rect 12986 3544 12992 3596
rect 13044 3544 13050 3596
rect 13078 3544 13084 3596
rect 13136 3584 13142 3596
rect 13245 3587 13303 3593
rect 13245 3584 13257 3587
rect 13136 3556 13257 3584
rect 13136 3544 13142 3556
rect 13245 3553 13257 3556
rect 13291 3553 13303 3587
rect 13245 3547 13303 3553
rect 14366 3544 14372 3596
rect 14424 3584 14430 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14424 3556 14749 3584
rect 14424 3544 14430 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 6104 3516 6132 3544
rect 6546 3516 6552 3528
rect 6104 3488 6552 3516
rect 6546 3476 6552 3488
rect 6604 3516 6610 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6604 3488 6745 3516
rect 6604 3476 6610 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9217 3519 9275 3525
rect 9217 3516 9229 3519
rect 9088 3488 9229 3516
rect 9088 3476 9094 3488
rect 9217 3485 9229 3488
rect 9263 3485 9275 3519
rect 14752 3516 14780 3547
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 15571 3593 15599 3692
rect 16209 3689 16221 3692
rect 16255 3689 16267 3723
rect 16209 3683 16267 3689
rect 15565 3587 15623 3593
rect 15565 3584 15577 3587
rect 15160 3556 15577 3584
rect 15160 3544 15166 3556
rect 15565 3553 15577 3556
rect 15611 3553 15623 3587
rect 15565 3547 15623 3553
rect 15657 3587 15715 3593
rect 15657 3553 15669 3587
rect 15703 3553 15715 3587
rect 16117 3587 16175 3593
rect 16117 3584 16129 3587
rect 15657 3547 15715 3553
rect 15948 3556 16129 3584
rect 15286 3516 15292 3528
rect 14752 3488 15292 3516
rect 9217 3479 9275 3485
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 1397 3451 1455 3457
rect 1397 3417 1409 3451
rect 1443 3448 1455 3451
rect 1854 3448 1860 3460
rect 1443 3420 1860 3448
rect 1443 3417 1455 3420
rect 1397 3411 1455 3417
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 4614 3408 4620 3460
rect 4672 3408 4678 3460
rect 6454 3448 6460 3460
rect 5000 3420 6460 3448
rect 1673 3383 1731 3389
rect 1673 3349 1685 3383
rect 1719 3380 1731 3383
rect 1762 3380 1768 3392
rect 1719 3352 1768 3380
rect 1719 3349 1731 3352
rect 1673 3343 1731 3349
rect 1762 3340 1768 3352
rect 1820 3380 1826 3392
rect 2222 3380 2228 3392
rect 1820 3352 2228 3380
rect 1820 3340 1826 3352
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 5000 3380 5028 3420
rect 6454 3408 6460 3420
rect 6512 3408 6518 3460
rect 15378 3408 15384 3460
rect 15436 3448 15442 3460
rect 15672 3448 15700 3547
rect 15948 3528 15976 3556
rect 16117 3553 16129 3556
rect 16163 3553 16175 3587
rect 16224 3584 16252 3683
rect 16298 3680 16304 3732
rect 16356 3720 16362 3732
rect 16758 3720 16764 3732
rect 16356 3692 16764 3720
rect 16356 3680 16362 3692
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 17037 3723 17095 3729
rect 17037 3720 17049 3723
rect 17000 3692 17049 3720
rect 17000 3680 17006 3692
rect 17037 3689 17049 3692
rect 17083 3689 17095 3723
rect 17037 3683 17095 3689
rect 17494 3680 17500 3732
rect 17552 3720 17558 3732
rect 17589 3723 17647 3729
rect 17589 3720 17601 3723
rect 17552 3692 17601 3720
rect 17552 3680 17558 3692
rect 17589 3689 17601 3692
rect 17635 3689 17647 3723
rect 17589 3683 17647 3689
rect 17862 3612 17868 3664
rect 17920 3652 17926 3664
rect 18702 3655 18760 3661
rect 18702 3652 18714 3655
rect 17920 3624 18714 3652
rect 17920 3612 17926 3624
rect 18702 3621 18714 3624
rect 18748 3621 18760 3655
rect 18702 3615 18760 3621
rect 16393 3587 16451 3593
rect 16393 3584 16405 3587
rect 16224 3556 16405 3584
rect 16117 3547 16175 3553
rect 16393 3553 16405 3556
rect 16439 3553 16451 3587
rect 16393 3547 16451 3553
rect 16853 3587 16911 3593
rect 16853 3553 16865 3587
rect 16899 3584 16911 3587
rect 16945 3587 17003 3593
rect 16945 3584 16957 3587
rect 16899 3556 16957 3584
rect 16899 3553 16911 3556
rect 16853 3547 16911 3553
rect 16945 3553 16957 3556
rect 16991 3553 17003 3587
rect 16945 3547 17003 3553
rect 17221 3587 17279 3593
rect 17221 3553 17233 3587
rect 17267 3553 17279 3587
rect 17221 3547 17279 3553
rect 15930 3476 15936 3528
rect 15988 3476 15994 3528
rect 16868 3516 16896 3547
rect 16040 3488 16896 3516
rect 16040 3448 16068 3488
rect 15436 3420 15700 3448
rect 15764 3420 16068 3448
rect 15436 3408 15442 3420
rect 15764 3392 15792 3420
rect 16114 3408 16120 3460
rect 16172 3448 16178 3460
rect 16485 3451 16543 3457
rect 16485 3448 16497 3451
rect 16172 3420 16497 3448
rect 16172 3408 16178 3420
rect 16485 3417 16497 3420
rect 16531 3448 16543 3451
rect 17236 3448 17264 3547
rect 18966 3544 18972 3596
rect 19024 3544 19030 3596
rect 16531 3420 17264 3448
rect 16531 3417 16543 3420
rect 16485 3411 16543 3417
rect 3375 3352 5028 3380
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 6362 3340 6368 3392
rect 6420 3340 6426 3392
rect 15746 3340 15752 3392
rect 15804 3340 15810 3392
rect 17310 3340 17316 3392
rect 17368 3340 17374 3392
rect 552 3290 19412 3312
rect 552 3238 2755 3290
rect 2807 3238 2819 3290
rect 2871 3238 2883 3290
rect 2935 3238 2947 3290
rect 2999 3238 3011 3290
rect 3063 3238 7470 3290
rect 7522 3238 7534 3290
rect 7586 3238 7598 3290
rect 7650 3238 7662 3290
rect 7714 3238 7726 3290
rect 7778 3238 12185 3290
rect 12237 3238 12249 3290
rect 12301 3238 12313 3290
rect 12365 3238 12377 3290
rect 12429 3238 12441 3290
rect 12493 3238 16900 3290
rect 16952 3238 16964 3290
rect 17016 3238 17028 3290
rect 17080 3238 17092 3290
rect 17144 3238 17156 3290
rect 17208 3238 19412 3290
rect 552 3216 19412 3238
rect 1854 3176 1860 3188
rect 1596 3148 1860 3176
rect 1302 2932 1308 2984
rect 1360 2932 1366 2984
rect 1596 2981 1624 3148
rect 1854 3136 1860 3148
rect 1912 3136 1918 3188
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 4798 3176 4804 3188
rect 3099 3148 4804 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7340 3148 7757 3176
rect 7340 3136 7346 3148
rect 7745 3145 7757 3148
rect 7791 3176 7803 3179
rect 8386 3176 8392 3188
rect 7791 3148 8392 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 8754 3136 8760 3188
rect 8812 3136 8818 3188
rect 10873 3179 10931 3185
rect 10873 3145 10885 3179
rect 10919 3176 10931 3179
rect 11330 3176 11336 3188
rect 10919 3148 11336 3176
rect 10919 3145 10931 3148
rect 10873 3139 10931 3145
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 12802 3136 12808 3188
rect 12860 3136 12866 3188
rect 12897 3179 12955 3185
rect 12897 3145 12909 3179
rect 12943 3176 12955 3179
rect 13078 3176 13084 3188
rect 12943 3148 13084 3176
rect 12943 3145 12955 3148
rect 12897 3139 12955 3145
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 15102 3136 15108 3188
rect 15160 3136 15166 3188
rect 15286 3136 15292 3188
rect 15344 3176 15350 3188
rect 15381 3179 15439 3185
rect 15381 3176 15393 3179
rect 15344 3148 15393 3176
rect 15344 3136 15350 3148
rect 15381 3145 15393 3148
rect 15427 3145 15439 3179
rect 15381 3139 15439 3145
rect 15746 3136 15752 3188
rect 15804 3136 15810 3188
rect 16114 3136 16120 3188
rect 16172 3136 16178 3188
rect 17129 3179 17187 3185
rect 17129 3145 17141 3179
rect 17175 3176 17187 3179
rect 17218 3176 17224 3188
rect 17175 3148 17224 3176
rect 17175 3145 17187 3148
rect 17129 3139 17187 3145
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2941 1731 2975
rect 1673 2935 1731 2941
rect 1688 2848 1716 2935
rect 2222 2932 2228 2984
rect 2280 2972 2286 2984
rect 3237 2975 3295 2981
rect 3237 2972 3249 2975
rect 2280 2944 3249 2972
rect 2280 2932 2286 2944
rect 3237 2941 3249 2944
rect 3283 2941 3295 2975
rect 3237 2935 3295 2941
rect 5534 2932 5540 2984
rect 5592 2972 5598 2984
rect 5721 2975 5779 2981
rect 5721 2972 5733 2975
rect 5592 2944 5733 2972
rect 5592 2932 5598 2944
rect 5721 2941 5733 2944
rect 5767 2941 5779 2975
rect 5721 2935 5779 2941
rect 6362 2932 6368 2984
rect 6420 2972 6426 2984
rect 7009 2975 7067 2981
rect 7009 2972 7021 2975
rect 6420 2944 7021 2972
rect 6420 2932 6426 2944
rect 7009 2941 7021 2944
rect 7055 2972 7067 2975
rect 7193 2975 7251 2981
rect 7193 2972 7205 2975
rect 7055 2944 7205 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 7193 2941 7205 2944
rect 7239 2941 7251 2975
rect 7193 2935 7251 2941
rect 7650 2932 7656 2984
rect 7708 2932 7714 2984
rect 8404 2972 8432 3136
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3040 12311 3043
rect 12526 3040 12532 3052
rect 12299 3012 12532 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12820 3040 12848 3136
rect 15562 3108 15568 3120
rect 14752 3080 15568 3108
rect 14752 3040 14780 3080
rect 15562 3068 15568 3080
rect 15620 3108 15626 3120
rect 15838 3108 15844 3120
rect 15620 3080 15844 3108
rect 15620 3068 15626 3080
rect 15838 3068 15844 3080
rect 15896 3068 15902 3120
rect 15948 3080 16712 3108
rect 12820 3012 14780 3040
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 8404 2944 8677 2972
rect 8665 2941 8677 2944
rect 8711 2941 8723 2975
rect 8665 2935 8723 2941
rect 12802 2932 12808 2984
rect 12860 2932 12866 2984
rect 14752 2981 14780 3012
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3040 14887 3043
rect 14875 3012 15332 3040
rect 14875 3009 14887 3012
rect 14829 3003 14887 3009
rect 15304 2981 15332 3012
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 15289 2975 15347 2981
rect 15289 2941 15301 2975
rect 15335 2972 15347 2975
rect 15657 2975 15715 2981
rect 15657 2972 15669 2975
rect 15335 2944 15669 2972
rect 15335 2941 15347 2944
rect 15289 2935 15347 2941
rect 15657 2941 15669 2944
rect 15703 2972 15715 2975
rect 15948 2972 15976 3080
rect 16298 3040 16304 3052
rect 16224 3012 16304 3040
rect 16224 2981 16252 3012
rect 16298 3000 16304 3012
rect 16356 3040 16362 3052
rect 16356 3012 16620 3040
rect 16356 3000 16362 3012
rect 15703 2944 15976 2972
rect 16209 2975 16267 2981
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 16209 2941 16221 2975
rect 16255 2941 16267 2975
rect 16209 2935 16267 2941
rect 1946 2913 1952 2916
rect 1940 2867 1952 2913
rect 1946 2864 1952 2867
rect 2004 2864 2010 2916
rect 2406 2864 2412 2916
rect 2464 2904 2470 2916
rect 3329 2907 3387 2913
rect 3329 2904 3341 2907
rect 2464 2876 3341 2904
rect 2464 2864 2470 2876
rect 3329 2873 3341 2876
rect 3375 2873 3387 2907
rect 3329 2867 3387 2873
rect 12008 2907 12066 2913
rect 12008 2873 12020 2907
rect 12054 2904 12066 2907
rect 13262 2904 13268 2916
rect 12054 2876 13268 2904
rect 12054 2873 12066 2876
rect 12008 2867 12066 2873
rect 13262 2864 13268 2876
rect 13320 2864 13326 2916
rect 15212 2904 15240 2935
rect 16482 2932 16488 2984
rect 16540 2932 16546 2984
rect 16592 2981 16620 3012
rect 16577 2975 16635 2981
rect 16577 2941 16589 2975
rect 16623 2941 16635 2975
rect 16577 2935 16635 2941
rect 16022 2904 16028 2916
rect 15212 2876 16028 2904
rect 16022 2864 16028 2876
rect 16080 2864 16086 2916
rect 16684 2904 16712 3080
rect 18506 3000 18512 3052
rect 18564 3040 18570 3052
rect 18966 3040 18972 3052
rect 18564 3012 18972 3040
rect 18564 3000 18570 3012
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 17037 2975 17095 2981
rect 17037 2972 17049 2975
rect 16816 2944 17049 2972
rect 16816 2932 16822 2944
rect 17037 2941 17049 2944
rect 17083 2941 17095 2975
rect 17037 2935 17095 2941
rect 17770 2904 17776 2916
rect 16592 2876 16712 2904
rect 16960 2876 17776 2904
rect 16592 2848 16620 2876
rect 1210 2796 1216 2848
rect 1268 2796 1274 2848
rect 1486 2796 1492 2848
rect 1544 2796 1550 2848
rect 1670 2796 1676 2848
rect 1728 2796 1734 2848
rect 5810 2796 5816 2848
rect 5868 2796 5874 2848
rect 6914 2796 6920 2848
rect 6972 2796 6978 2848
rect 15286 2796 15292 2848
rect 15344 2836 15350 2848
rect 15930 2836 15936 2848
rect 15344 2808 15936 2836
rect 15344 2796 15350 2808
rect 15930 2796 15936 2808
rect 15988 2796 15994 2848
rect 16390 2796 16396 2848
rect 16448 2796 16454 2848
rect 16574 2796 16580 2848
rect 16632 2796 16638 2848
rect 16960 2845 16988 2876
rect 17770 2864 17776 2876
rect 17828 2904 17834 2916
rect 18242 2907 18300 2913
rect 18242 2904 18254 2907
rect 17828 2876 18254 2904
rect 17828 2864 17834 2876
rect 18242 2873 18254 2876
rect 18288 2873 18300 2907
rect 18242 2867 18300 2873
rect 16669 2839 16727 2845
rect 16669 2805 16681 2839
rect 16715 2836 16727 2839
rect 16945 2839 17003 2845
rect 16945 2836 16957 2839
rect 16715 2808 16957 2836
rect 16715 2805 16727 2808
rect 16669 2799 16727 2805
rect 16945 2805 16957 2808
rect 16991 2805 17003 2839
rect 16945 2799 17003 2805
rect 552 2746 19571 2768
rect 552 2694 5112 2746
rect 5164 2694 5176 2746
rect 5228 2694 5240 2746
rect 5292 2694 5304 2746
rect 5356 2694 5368 2746
rect 5420 2694 9827 2746
rect 9879 2694 9891 2746
rect 9943 2694 9955 2746
rect 10007 2694 10019 2746
rect 10071 2694 10083 2746
rect 10135 2694 14542 2746
rect 14594 2694 14606 2746
rect 14658 2694 14670 2746
rect 14722 2694 14734 2746
rect 14786 2694 14798 2746
rect 14850 2694 19257 2746
rect 19309 2694 19321 2746
rect 19373 2694 19385 2746
rect 19437 2694 19449 2746
rect 19501 2694 19513 2746
rect 19565 2694 19571 2746
rect 552 2672 19571 2694
rect 1486 2592 1492 2644
rect 1544 2632 1550 2644
rect 1946 2632 1952 2644
rect 1544 2604 1952 2632
rect 1544 2592 1550 2604
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 3694 2632 3700 2644
rect 2792 2604 3700 2632
rect 1673 2567 1731 2573
rect 1673 2564 1685 2567
rect 1228 2536 1685 2564
rect 1228 2508 1256 2536
rect 1673 2533 1685 2536
rect 1719 2564 1731 2567
rect 1762 2564 1768 2576
rect 1719 2536 1768 2564
rect 1719 2533 1731 2536
rect 1673 2527 1731 2533
rect 1762 2524 1768 2536
rect 1820 2524 1826 2576
rect 1854 2524 1860 2576
rect 1912 2524 1918 2576
rect 1964 2564 1992 2592
rect 1964 2536 2360 2564
rect 1210 2456 1216 2508
rect 1268 2456 1274 2508
rect 1486 2456 1492 2508
rect 1544 2456 1550 2508
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2496 1639 2499
rect 1872 2496 1900 2524
rect 1627 2468 1900 2496
rect 2041 2499 2099 2505
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 2041 2465 2053 2499
rect 2087 2496 2099 2499
rect 2222 2496 2228 2508
rect 2087 2468 2228 2496
rect 2087 2465 2099 2468
rect 2041 2459 2099 2465
rect 1121 2431 1179 2437
rect 1121 2397 1133 2431
rect 1167 2428 1179 2431
rect 1302 2428 1308 2440
rect 1167 2400 1308 2428
rect 1167 2397 1179 2400
rect 1121 2391 1179 2397
rect 1302 2388 1308 2400
rect 1360 2428 1366 2440
rect 2056 2428 2084 2459
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 2332 2505 2360 2536
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2465 2375 2499
rect 2317 2459 2375 2465
rect 2409 2499 2467 2505
rect 2409 2465 2421 2499
rect 2455 2496 2467 2499
rect 2498 2496 2504 2508
rect 2455 2468 2504 2496
rect 2455 2465 2467 2468
rect 2409 2459 2467 2465
rect 2498 2456 2504 2468
rect 2556 2496 2562 2508
rect 2792 2505 2820 2604
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 3789 2635 3847 2641
rect 3789 2601 3801 2635
rect 3835 2632 3847 2635
rect 4154 2632 4160 2644
rect 3835 2604 4160 2632
rect 3835 2601 3847 2604
rect 3789 2595 3847 2601
rect 4154 2592 4160 2604
rect 4212 2632 4218 2644
rect 4614 2632 4620 2644
rect 4212 2604 4620 2632
rect 4212 2592 4218 2604
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2632 5319 2635
rect 5626 2632 5632 2644
rect 5307 2604 5632 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6362 2592 6368 2644
rect 6420 2592 6426 2644
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 7432 2604 10364 2632
rect 7432 2592 7438 2604
rect 3145 2567 3203 2573
rect 3145 2533 3157 2567
rect 3191 2564 3203 2567
rect 3234 2564 3240 2576
rect 3191 2536 3240 2564
rect 3191 2533 3203 2536
rect 3145 2527 3203 2533
rect 3234 2524 3240 2536
rect 3292 2564 3298 2576
rect 4341 2567 4399 2573
rect 3292 2536 3740 2564
rect 3292 2524 3298 2536
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 2556 2468 2789 2496
rect 2556 2456 2562 2468
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 3053 2499 3111 2505
rect 3053 2496 3065 2499
rect 2777 2459 2835 2465
rect 2884 2468 3065 2496
rect 1360 2400 2084 2428
rect 1360 2388 1366 2400
rect 1394 2252 1400 2304
rect 1452 2252 1458 2304
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 2884 2301 2912 2468
rect 3053 2465 3065 2468
rect 3099 2465 3111 2499
rect 3053 2459 3111 2465
rect 3602 2456 3608 2508
rect 3660 2456 3666 2508
rect 3712 2505 3740 2536
rect 4341 2533 4353 2567
rect 4387 2564 4399 2567
rect 4893 2567 4951 2573
rect 4893 2564 4905 2567
rect 4387 2536 4905 2564
rect 4387 2533 4399 2536
rect 4341 2527 4399 2533
rect 4893 2533 4905 2536
rect 4939 2564 4951 2567
rect 5534 2564 5540 2576
rect 4939 2536 5540 2564
rect 4939 2533 4951 2536
rect 4893 2527 4951 2533
rect 5534 2524 5540 2536
rect 5592 2524 5598 2576
rect 3697 2499 3755 2505
rect 3697 2465 3709 2499
rect 3743 2465 3755 2499
rect 3697 2459 3755 2465
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2496 4215 2499
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 4203 2468 4261 2496
rect 4203 2465 4215 2468
rect 4157 2459 4215 2465
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2465 4583 2499
rect 4525 2459 4583 2465
rect 4172 2428 4200 2459
rect 3528 2400 4200 2428
rect 3528 2304 3556 2400
rect 4065 2363 4123 2369
rect 4065 2360 4077 2363
rect 3712 2332 4077 2360
rect 3712 2304 3740 2332
rect 4065 2329 4077 2332
rect 4111 2360 4123 2363
rect 4540 2360 4568 2459
rect 4982 2456 4988 2508
rect 5040 2456 5046 2508
rect 5644 2505 5672 2592
rect 5810 2524 5816 2576
rect 5868 2564 5874 2576
rect 6794 2567 6852 2573
rect 6794 2564 6806 2567
rect 5868 2536 6806 2564
rect 5868 2524 5874 2536
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2465 5227 2499
rect 5169 2459 5227 2465
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2465 5687 2499
rect 5828 2496 5856 2524
rect 6380 2508 6408 2536
rect 6794 2533 6806 2536
rect 6840 2533 6852 2567
rect 6794 2527 6852 2533
rect 8386 2524 8392 2576
rect 8444 2524 8450 2576
rect 8588 2536 9076 2564
rect 5997 2499 6055 2505
rect 5997 2496 6009 2499
rect 5828 2468 6009 2496
rect 5629 2459 5687 2465
rect 5997 2465 6009 2468
rect 6043 2465 6055 2499
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5997 2459 6055 2465
rect 6104 2468 6285 2496
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2428 4675 2431
rect 5184 2428 5212 2459
rect 4663 2400 5212 2428
rect 4663 2397 4675 2400
rect 4617 2391 4675 2397
rect 5000 2372 5028 2400
rect 4111 2332 4568 2360
rect 4111 2329 4123 2332
rect 4065 2323 4123 2329
rect 4982 2320 4988 2372
rect 5040 2320 5046 2372
rect 6104 2304 6132 2468
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 6362 2456 6368 2508
rect 6420 2456 6426 2508
rect 6546 2456 6552 2508
rect 6604 2456 6610 2508
rect 8297 2499 8355 2505
rect 8297 2465 8309 2499
rect 8343 2496 8355 2499
rect 8404 2496 8432 2524
rect 8588 2505 8616 2536
rect 8343 2468 8432 2496
rect 8573 2499 8631 2505
rect 8343 2465 8355 2468
rect 8297 2459 8355 2465
rect 8573 2465 8585 2499
rect 8619 2465 8631 2499
rect 8573 2459 8631 2465
rect 8202 2388 8208 2440
rect 8260 2428 8266 2440
rect 8588 2428 8616 2459
rect 8662 2456 8668 2508
rect 8720 2456 8726 2508
rect 9048 2505 9076 2536
rect 9306 2524 9312 2576
rect 9364 2564 9370 2576
rect 9585 2567 9643 2573
rect 9585 2564 9597 2567
rect 9364 2536 9597 2564
rect 9364 2524 9370 2536
rect 9585 2533 9597 2536
rect 9631 2564 9643 2567
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 9631 2536 10241 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 8757 2499 8815 2505
rect 8757 2465 8769 2499
rect 8803 2465 8815 2499
rect 8757 2459 8815 2465
rect 9033 2499 9091 2505
rect 9033 2465 9045 2499
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 8260 2400 8616 2428
rect 8260 2388 8266 2400
rect 7929 2363 7987 2369
rect 7929 2329 7941 2363
rect 7975 2360 7987 2363
rect 8680 2360 8708 2456
rect 7975 2332 8708 2360
rect 7975 2329 7987 2332
rect 7929 2323 7987 2329
rect 2869 2295 2927 2301
rect 2869 2292 2881 2295
rect 2648 2264 2881 2292
rect 2648 2252 2654 2264
rect 2869 2261 2881 2264
rect 2915 2261 2927 2295
rect 2869 2255 2927 2261
rect 3510 2252 3516 2304
rect 3568 2252 3574 2304
rect 3694 2252 3700 2304
rect 3752 2252 3758 2304
rect 5534 2252 5540 2304
rect 5592 2252 5598 2304
rect 6086 2252 6092 2304
rect 6144 2252 6150 2304
rect 8202 2252 8208 2304
rect 8260 2252 8266 2304
rect 8478 2252 8484 2304
rect 8536 2292 8542 2304
rect 8772 2292 8800 2459
rect 9416 2428 9444 2459
rect 9674 2456 9680 2508
rect 9732 2456 9738 2508
rect 10336 2505 10364 2604
rect 10594 2592 10600 2644
rect 10652 2592 10658 2644
rect 13817 2635 13875 2641
rect 13817 2601 13829 2635
rect 13863 2632 13875 2635
rect 13863 2604 14780 2632
rect 13863 2601 13875 2604
rect 13817 2595 13875 2601
rect 13446 2564 13452 2576
rect 12544 2536 13452 2564
rect 12544 2508 12572 2536
rect 13446 2524 13452 2536
rect 13504 2564 13510 2576
rect 14752 2564 14780 2604
rect 15286 2592 15292 2644
rect 15344 2632 15350 2644
rect 15473 2635 15531 2641
rect 15473 2632 15485 2635
rect 15344 2604 15485 2632
rect 15344 2592 15350 2604
rect 15473 2601 15485 2604
rect 15519 2601 15531 2635
rect 15473 2595 15531 2601
rect 15654 2592 15660 2644
rect 15712 2592 15718 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 16761 2635 16819 2641
rect 16761 2632 16773 2635
rect 16632 2604 16773 2632
rect 16632 2592 16638 2604
rect 16761 2601 16773 2604
rect 16807 2601 16819 2635
rect 16761 2595 16819 2601
rect 17129 2635 17187 2641
rect 17129 2601 17141 2635
rect 17175 2632 17187 2635
rect 17310 2632 17316 2644
rect 17175 2604 17316 2632
rect 17175 2601 17187 2604
rect 17129 2595 17187 2601
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17589 2635 17647 2641
rect 17589 2601 17601 2635
rect 17635 2632 17647 2635
rect 17862 2632 17868 2644
rect 17635 2604 17868 2632
rect 17635 2601 17647 2604
rect 17589 2595 17647 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 15672 2564 15700 2592
rect 16485 2567 16543 2573
rect 16485 2564 16497 2567
rect 13504 2536 13952 2564
rect 14752 2536 15700 2564
rect 16316 2536 16497 2564
rect 13504 2524 13510 2536
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 10045 2499 10103 2505
rect 9815 2468 9996 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 9416 2400 9628 2428
rect 9600 2304 9628 2400
rect 9968 2360 9996 2468
rect 10045 2465 10057 2499
rect 10091 2496 10103 2499
rect 10321 2499 10379 2505
rect 10091 2468 10272 2496
rect 10091 2465 10103 2468
rect 10045 2459 10103 2465
rect 10244 2440 10272 2468
rect 10321 2465 10333 2499
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 10413 2499 10471 2505
rect 10413 2465 10425 2499
rect 10459 2496 10471 2499
rect 10870 2496 10876 2508
rect 10459 2468 10876 2496
rect 10459 2465 10471 2468
rect 10413 2459 10471 2465
rect 10226 2388 10232 2440
rect 10284 2388 10290 2440
rect 10428 2360 10456 2459
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 10965 2499 11023 2505
rect 10965 2465 10977 2499
rect 11011 2465 11023 2499
rect 10965 2459 11023 2465
rect 9968 2332 10456 2360
rect 8536 2264 8800 2292
rect 8849 2295 8907 2301
rect 8536 2252 8542 2264
rect 8849 2261 8861 2295
rect 8895 2292 8907 2295
rect 8938 2292 8944 2304
rect 8895 2264 8944 2292
rect 8895 2261 8907 2264
rect 8849 2255 8907 2261
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 9122 2252 9128 2304
rect 9180 2252 9186 2304
rect 9582 2252 9588 2304
rect 9640 2252 9646 2304
rect 9950 2252 9956 2304
rect 10008 2252 10014 2304
rect 10134 2252 10140 2304
rect 10192 2292 10198 2304
rect 10980 2292 11008 2459
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 11112 2468 11437 2496
rect 11112 2456 11118 2468
rect 11425 2465 11437 2468
rect 11471 2496 11483 2499
rect 12437 2499 12495 2505
rect 11471 2468 12020 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11992 2304 12020 2468
rect 12437 2465 12449 2499
rect 12483 2496 12495 2499
rect 12526 2496 12532 2508
rect 12483 2468 12532 2496
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 12526 2456 12532 2468
rect 12584 2456 12590 2508
rect 12710 2505 12716 2508
rect 12704 2496 12716 2505
rect 12671 2468 12716 2496
rect 12704 2459 12716 2468
rect 12710 2456 12716 2459
rect 12768 2456 12774 2508
rect 13924 2505 13952 2536
rect 13909 2499 13967 2505
rect 13909 2465 13921 2499
rect 13955 2465 13967 2499
rect 13909 2459 13967 2465
rect 13998 2456 14004 2508
rect 14056 2496 14062 2508
rect 14165 2499 14223 2505
rect 14165 2496 14177 2499
rect 14056 2468 14177 2496
rect 14056 2456 14062 2468
rect 14165 2465 14177 2468
rect 14211 2465 14223 2499
rect 14165 2459 14223 2465
rect 15565 2499 15623 2505
rect 15565 2465 15577 2499
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 15580 2428 15608 2459
rect 15654 2456 15660 2508
rect 15712 2456 15718 2508
rect 16114 2456 16120 2508
rect 16172 2496 16178 2508
rect 16316 2505 16344 2536
rect 16485 2533 16497 2536
rect 16531 2533 16543 2567
rect 16485 2527 16543 2533
rect 17770 2524 17776 2576
rect 17828 2524 17834 2576
rect 16301 2499 16359 2505
rect 16301 2496 16313 2499
rect 16172 2468 16313 2496
rect 16172 2456 16178 2468
rect 16301 2465 16313 2468
rect 16347 2465 16359 2499
rect 16301 2459 16359 2465
rect 16393 2499 16451 2505
rect 16393 2465 16405 2499
rect 16439 2465 16451 2499
rect 16393 2459 16451 2465
rect 16669 2499 16727 2505
rect 16669 2465 16681 2499
rect 16715 2465 16727 2499
rect 16669 2459 16727 2465
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2496 17095 2499
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17083 2468 17693 2496
rect 17083 2465 17095 2468
rect 17037 2459 17095 2465
rect 17681 2465 17693 2468
rect 17727 2496 17739 2499
rect 17788 2496 17816 2524
rect 17727 2468 17816 2496
rect 17727 2465 17739 2468
rect 17681 2459 17739 2465
rect 16408 2428 16436 2459
rect 15580 2400 16436 2428
rect 15764 2304 15792 2400
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 16684 2360 16712 2459
rect 16448 2332 16712 2360
rect 16448 2320 16454 2332
rect 10192 2264 11008 2292
rect 10192 2252 10198 2264
rect 11330 2252 11336 2304
rect 11388 2252 11394 2304
rect 11974 2252 11980 2304
rect 12032 2252 12038 2304
rect 14274 2252 14280 2304
rect 14332 2292 14338 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 14332 2264 15301 2292
rect 14332 2252 14338 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 15746 2252 15752 2304
rect 15804 2252 15810 2304
rect 15930 2252 15936 2304
rect 15988 2292 15994 2304
rect 16209 2295 16267 2301
rect 16209 2292 16221 2295
rect 15988 2264 16221 2292
rect 15988 2252 15994 2264
rect 16209 2261 16221 2264
rect 16255 2261 16267 2295
rect 16209 2255 16267 2261
rect 19058 2252 19064 2304
rect 19116 2252 19122 2304
rect 552 2202 19412 2224
rect 552 2150 2755 2202
rect 2807 2150 2819 2202
rect 2871 2150 2883 2202
rect 2935 2150 2947 2202
rect 2999 2150 3011 2202
rect 3063 2150 7470 2202
rect 7522 2150 7534 2202
rect 7586 2150 7598 2202
rect 7650 2150 7662 2202
rect 7714 2150 7726 2202
rect 7778 2150 12185 2202
rect 12237 2150 12249 2202
rect 12301 2150 12313 2202
rect 12365 2150 12377 2202
rect 12429 2150 12441 2202
rect 12493 2150 16900 2202
rect 16952 2150 16964 2202
rect 17016 2150 17028 2202
rect 17080 2150 17092 2202
rect 17144 2150 17156 2202
rect 17208 2150 19412 2202
rect 552 2128 19412 2150
rect 1210 2048 1216 2100
rect 1268 2048 1274 2100
rect 1305 2091 1363 2097
rect 1305 2057 1317 2091
rect 1351 2088 1363 2091
rect 1394 2088 1400 2100
rect 1351 2060 1400 2088
rect 1351 2057 1363 2060
rect 1305 2051 1363 2057
rect 1394 2048 1400 2060
rect 1452 2048 1458 2100
rect 1857 2091 1915 2097
rect 1857 2057 1869 2091
rect 1903 2088 1915 2091
rect 2498 2088 2504 2100
rect 1903 2060 2504 2088
rect 1903 2057 1915 2060
rect 1857 2051 1915 2057
rect 2498 2048 2504 2060
rect 2556 2088 2562 2100
rect 2774 2088 2780 2100
rect 2556 2060 2780 2088
rect 2556 2048 2562 2060
rect 2774 2048 2780 2060
rect 2832 2048 2838 2100
rect 2961 2091 3019 2097
rect 2961 2057 2973 2091
rect 3007 2088 3019 2091
rect 3510 2088 3516 2100
rect 3007 2060 3516 2088
rect 3007 2057 3019 2060
rect 2961 2051 3019 2057
rect 3510 2048 3516 2060
rect 3568 2048 3574 2100
rect 4154 2088 4160 2100
rect 3804 2060 4160 2088
rect 1228 1952 1256 2048
rect 1136 1924 1256 1952
rect 1136 1893 1164 1924
rect 1121 1887 1179 1893
rect 1121 1853 1133 1887
rect 1167 1853 1179 1887
rect 1121 1847 1179 1853
rect 1210 1844 1216 1896
rect 1268 1844 1274 1896
rect 1412 1884 1440 2048
rect 3421 2023 3479 2029
rect 3421 1989 3433 2023
rect 3467 2020 3479 2023
rect 3804 2020 3832 2060
rect 4154 2048 4160 2060
rect 4212 2048 4218 2100
rect 7006 2048 7012 2100
rect 7064 2088 7070 2100
rect 7466 2088 7472 2100
rect 7064 2060 7472 2088
rect 7064 2048 7070 2060
rect 7466 2048 7472 2060
rect 7524 2048 7530 2100
rect 7561 2091 7619 2097
rect 7561 2057 7573 2091
rect 7607 2088 7619 2091
rect 8202 2088 8208 2100
rect 7607 2060 8208 2088
rect 7607 2057 7619 2060
rect 7561 2051 7619 2057
rect 8202 2048 8208 2060
rect 8260 2048 8266 2100
rect 8570 2048 8576 2100
rect 8628 2088 8634 2100
rect 8628 2060 9996 2088
rect 8628 2048 8634 2060
rect 3467 1992 3832 2020
rect 3467 1989 3479 1992
rect 3421 1983 3479 1989
rect 2222 1952 2228 1964
rect 2056 1924 2228 1952
rect 2056 1893 2084 1924
rect 2222 1912 2228 1924
rect 2280 1952 2286 1964
rect 2406 1952 2412 1964
rect 2280 1924 2412 1952
rect 2280 1912 2286 1924
rect 2406 1912 2412 1924
rect 2464 1912 2470 1964
rect 3234 1952 3240 1964
rect 2516 1924 3240 1952
rect 2516 1893 2544 1924
rect 3234 1912 3240 1924
rect 3292 1912 3298 1964
rect 3694 1952 3700 1964
rect 3344 1924 3700 1952
rect 1489 1887 1547 1893
rect 1489 1884 1501 1887
rect 1412 1856 1501 1884
rect 1489 1853 1501 1856
rect 1535 1853 1547 1887
rect 1489 1847 1547 1853
rect 1949 1887 2007 1893
rect 1949 1853 1961 1887
rect 1995 1884 2007 1887
rect 2041 1887 2099 1893
rect 2041 1884 2053 1887
rect 1995 1856 2053 1884
rect 1995 1853 2007 1856
rect 1949 1847 2007 1853
rect 2041 1853 2053 1856
rect 2087 1853 2099 1887
rect 2041 1847 2099 1853
rect 2501 1887 2559 1893
rect 2501 1853 2513 1887
rect 2547 1853 2559 1887
rect 2501 1847 2559 1853
rect 2590 1844 2596 1896
rect 2648 1844 2654 1896
rect 2685 1887 2743 1893
rect 2685 1853 2697 1887
rect 2731 1853 2743 1887
rect 2685 1847 2743 1853
rect 1581 1819 1639 1825
rect 1581 1785 1593 1819
rect 1627 1816 1639 1819
rect 2608 1816 2636 1844
rect 1627 1788 2636 1816
rect 2700 1816 2728 1847
rect 2774 1844 2780 1896
rect 2832 1886 2838 1896
rect 3344 1893 3372 1924
rect 3694 1912 3700 1924
rect 3752 1912 3758 1964
rect 2869 1887 2927 1893
rect 2869 1886 2881 1887
rect 2832 1858 2881 1886
rect 2832 1844 2838 1858
rect 2869 1853 2881 1858
rect 2915 1853 2927 1887
rect 2869 1847 2927 1853
rect 3329 1887 3387 1893
rect 3329 1853 3341 1887
rect 3375 1853 3387 1887
rect 3329 1847 3387 1853
rect 3344 1816 3372 1847
rect 3510 1844 3516 1896
rect 3568 1844 3574 1896
rect 3605 1887 3663 1893
rect 3605 1853 3617 1887
rect 3651 1884 3663 1887
rect 3804 1884 3832 1992
rect 7285 2023 7343 2029
rect 7285 1989 7297 2023
rect 7331 2020 7343 2023
rect 8478 2020 8484 2032
rect 7331 1992 8484 2020
rect 7331 1989 7343 1992
rect 7285 1983 7343 1989
rect 6914 1912 6920 1964
rect 6972 1952 6978 1964
rect 6972 1924 7512 1952
rect 6972 1912 6978 1924
rect 3651 1856 3832 1884
rect 3651 1853 3663 1856
rect 3605 1847 3663 1853
rect 3878 1844 3884 1896
rect 3936 1884 3942 1896
rect 5626 1893 5632 1896
rect 5353 1887 5411 1893
rect 5353 1884 5365 1887
rect 3936 1856 5365 1884
rect 3936 1844 3942 1856
rect 5353 1853 5365 1856
rect 5399 1853 5411 1887
rect 5620 1884 5632 1893
rect 5587 1856 5632 1884
rect 5353 1847 5411 1853
rect 5620 1847 5632 1856
rect 5626 1844 5632 1847
rect 5684 1844 5690 1896
rect 5902 1844 5908 1896
rect 5960 1844 5966 1896
rect 7101 1887 7159 1893
rect 7101 1853 7113 1887
rect 7147 1884 7159 1887
rect 7190 1884 7196 1896
rect 7147 1856 7196 1884
rect 7147 1853 7159 1856
rect 7101 1847 7159 1853
rect 7190 1844 7196 1856
rect 7248 1844 7254 1896
rect 7484 1893 7512 1924
rect 7558 1912 7564 1964
rect 7616 1952 7622 1964
rect 7834 1952 7840 1964
rect 7616 1924 7840 1952
rect 7616 1912 7622 1924
rect 7760 1893 7788 1924
rect 7834 1912 7840 1924
rect 7892 1912 7898 1964
rect 8220 1893 8248 1992
rect 8478 1980 8484 1992
rect 8536 1980 8542 2032
rect 9968 2020 9996 2060
rect 10226 2048 10232 2100
rect 10284 2088 10290 2100
rect 10413 2091 10471 2097
rect 10413 2088 10425 2091
rect 10284 2060 10425 2088
rect 10284 2048 10290 2060
rect 10413 2057 10425 2060
rect 10459 2057 10471 2091
rect 10413 2051 10471 2057
rect 10689 2091 10747 2097
rect 10689 2057 10701 2091
rect 10735 2088 10747 2091
rect 11330 2088 11336 2100
rect 10735 2060 11336 2088
rect 10735 2057 10747 2060
rect 10689 2051 10747 2057
rect 11330 2048 11336 2060
rect 11388 2048 11394 2100
rect 12066 2048 12072 2100
rect 12124 2088 12130 2100
rect 12345 2091 12403 2097
rect 12345 2088 12357 2091
rect 12124 2060 12357 2088
rect 12124 2048 12130 2060
rect 12345 2057 12357 2060
rect 12391 2057 12403 2091
rect 12345 2051 12403 2057
rect 12529 2091 12587 2097
rect 12529 2057 12541 2091
rect 12575 2088 12587 2091
rect 12710 2088 12716 2100
rect 12575 2060 12716 2088
rect 12575 2057 12587 2060
rect 12529 2051 12587 2057
rect 12710 2048 12716 2060
rect 12768 2088 12774 2100
rect 12805 2091 12863 2097
rect 12805 2088 12817 2091
rect 12768 2060 12817 2088
rect 12768 2048 12774 2060
rect 12805 2057 12817 2060
rect 12851 2057 12863 2091
rect 12805 2051 12863 2057
rect 13262 2048 13268 2100
rect 13320 2088 13326 2100
rect 14553 2091 14611 2097
rect 14553 2088 14565 2091
rect 13320 2060 14565 2088
rect 13320 2048 13326 2060
rect 14553 2057 14565 2060
rect 14599 2088 14611 2091
rect 15654 2088 15660 2100
rect 14599 2060 15660 2088
rect 14599 2057 14611 2060
rect 14553 2051 14611 2057
rect 10134 2020 10140 2032
rect 9968 1992 10140 2020
rect 10134 1980 10140 1992
rect 10192 1980 10198 2032
rect 11974 1980 11980 2032
rect 12032 2020 12038 2032
rect 13998 2020 14004 2032
rect 12032 1992 14004 2020
rect 12032 1980 12038 1992
rect 9030 1952 9036 1964
rect 8404 1924 9036 1952
rect 8404 1896 8432 1924
rect 9030 1912 9036 1924
rect 9088 1912 9094 1964
rect 10778 1912 10784 1964
rect 10836 1952 10842 1964
rect 10965 1955 11023 1961
rect 10965 1952 10977 1955
rect 10836 1924 10977 1952
rect 10836 1912 10842 1924
rect 10965 1921 10977 1924
rect 11011 1921 11023 1955
rect 10965 1915 11023 1921
rect 7469 1887 7527 1893
rect 7469 1853 7481 1887
rect 7515 1853 7527 1887
rect 7469 1847 7527 1853
rect 7745 1887 7803 1893
rect 7745 1853 7757 1887
rect 7791 1853 7803 1887
rect 7745 1847 7803 1853
rect 8205 1887 8263 1893
rect 8205 1853 8217 1887
rect 8251 1853 8263 1887
rect 8205 1847 8263 1853
rect 8386 1844 8392 1896
rect 8444 1844 8450 1896
rect 8481 1887 8539 1893
rect 8481 1853 8493 1887
rect 8527 1884 8539 1887
rect 8757 1887 8815 1893
rect 8757 1884 8769 1887
rect 8527 1856 8769 1884
rect 8527 1853 8539 1856
rect 8481 1847 8539 1853
rect 8757 1853 8769 1856
rect 8803 1853 8815 1887
rect 9674 1884 9680 1896
rect 8757 1847 8815 1853
rect 8864 1856 9680 1884
rect 2700 1788 3372 1816
rect 3528 1816 3556 1844
rect 4126 1819 4184 1825
rect 4126 1816 4138 1819
rect 3528 1788 4138 1816
rect 1627 1785 1639 1788
rect 1581 1779 1639 1785
rect 4126 1785 4138 1788
rect 4172 1785 4184 1819
rect 4126 1779 4184 1785
rect 4430 1776 4436 1828
rect 4488 1816 4494 1828
rect 5920 1816 5948 1844
rect 7837 1819 7895 1825
rect 4488 1788 5948 1816
rect 6104 1788 7788 1816
rect 4488 1776 4494 1788
rect 1029 1751 1087 1757
rect 1029 1717 1041 1751
rect 1075 1748 1087 1751
rect 1486 1748 1492 1760
rect 1075 1720 1492 1748
rect 1075 1717 1087 1720
rect 1029 1711 1087 1717
rect 1486 1708 1492 1720
rect 1544 1708 1550 1760
rect 2133 1751 2191 1757
rect 2133 1717 2145 1751
rect 2179 1748 2191 1751
rect 2409 1751 2467 1757
rect 2409 1748 2421 1751
rect 2179 1720 2421 1748
rect 2179 1717 2191 1720
rect 2133 1711 2191 1717
rect 2409 1717 2421 1720
rect 2455 1748 2467 1751
rect 2682 1748 2688 1760
rect 2455 1720 2688 1748
rect 2455 1717 2467 1720
rect 2409 1711 2467 1717
rect 2682 1708 2688 1720
rect 2740 1708 2746 1760
rect 3697 1751 3755 1757
rect 3697 1717 3709 1751
rect 3743 1748 3755 1751
rect 4890 1748 4896 1760
rect 3743 1720 4896 1748
rect 3743 1717 3755 1720
rect 3697 1711 3755 1717
rect 4890 1708 4896 1720
rect 4948 1708 4954 1760
rect 5261 1751 5319 1757
rect 5261 1717 5273 1751
rect 5307 1748 5319 1751
rect 6104 1748 6132 1788
rect 5307 1720 6132 1748
rect 6733 1751 6791 1757
rect 5307 1717 5319 1720
rect 5261 1711 5319 1717
rect 6733 1717 6745 1751
rect 6779 1748 6791 1751
rect 7374 1748 7380 1760
rect 6779 1720 7380 1748
rect 6779 1717 6791 1720
rect 6733 1711 6791 1717
rect 7374 1708 7380 1720
rect 7432 1708 7438 1760
rect 7760 1748 7788 1788
rect 7837 1785 7849 1819
rect 7883 1816 7895 1819
rect 8113 1819 8171 1825
rect 8113 1816 8125 1819
rect 7883 1788 8125 1816
rect 7883 1785 7895 1788
rect 7837 1779 7895 1785
rect 8113 1785 8125 1788
rect 8159 1816 8171 1819
rect 8496 1816 8524 1847
rect 8864 1816 8892 1856
rect 9674 1844 9680 1856
rect 9732 1844 9738 1896
rect 12452 1893 12480 1992
rect 13998 1980 14004 1992
rect 14056 1980 14062 2032
rect 13648 1924 13860 1952
rect 10597 1887 10655 1893
rect 10597 1853 10609 1887
rect 10643 1853 10655 1887
rect 10597 1847 10655 1853
rect 12437 1887 12495 1893
rect 12437 1853 12449 1887
rect 12483 1853 12495 1887
rect 12437 1847 12495 1853
rect 12897 1887 12955 1893
rect 12897 1853 12909 1887
rect 12943 1853 12955 1887
rect 12897 1847 12955 1853
rect 8159 1788 8524 1816
rect 8588 1788 8892 1816
rect 8159 1785 8171 1788
rect 8113 1779 8171 1785
rect 8588 1748 8616 1788
rect 8938 1776 8944 1828
rect 8996 1816 9002 1828
rect 9278 1819 9336 1825
rect 9278 1816 9290 1819
rect 8996 1788 9290 1816
rect 8996 1776 9002 1788
rect 9278 1785 9290 1788
rect 9324 1816 9336 1819
rect 10318 1816 10324 1828
rect 9324 1788 10324 1816
rect 9324 1785 9336 1788
rect 9278 1779 9336 1785
rect 10318 1776 10324 1788
rect 10376 1776 10382 1828
rect 10612 1760 10640 1847
rect 11232 1819 11290 1825
rect 11232 1785 11244 1819
rect 11278 1816 11290 1819
rect 11422 1816 11428 1828
rect 11278 1788 11428 1816
rect 11278 1785 11290 1788
rect 11232 1779 11290 1785
rect 11422 1776 11428 1788
rect 11480 1776 11486 1828
rect 12912 1816 12940 1847
rect 13078 1844 13084 1896
rect 13136 1884 13142 1896
rect 13648 1893 13676 1924
rect 13832 1893 13860 1924
rect 13357 1887 13415 1893
rect 13357 1884 13369 1887
rect 13136 1856 13369 1884
rect 13136 1844 13142 1856
rect 13357 1853 13369 1856
rect 13403 1884 13415 1887
rect 13633 1887 13691 1893
rect 13633 1884 13645 1887
rect 13403 1856 13645 1884
rect 13403 1853 13415 1856
rect 13357 1847 13415 1853
rect 13633 1853 13645 1856
rect 13679 1853 13691 1887
rect 13633 1847 13691 1853
rect 13725 1887 13783 1893
rect 13725 1853 13737 1887
rect 13771 1853 13783 1887
rect 13725 1847 13783 1853
rect 13817 1887 13875 1893
rect 13817 1853 13829 1887
rect 13863 1853 13875 1887
rect 13817 1847 13875 1853
rect 14093 1887 14151 1893
rect 14093 1853 14105 1887
rect 14139 1884 14151 1887
rect 14182 1884 14188 1896
rect 14139 1856 14188 1884
rect 14139 1853 14151 1856
rect 14093 1847 14151 1853
rect 13740 1816 13768 1847
rect 14108 1816 14136 1847
rect 14182 1844 14188 1856
rect 14240 1844 14246 1896
rect 14461 1887 14519 1893
rect 14461 1853 14473 1887
rect 14507 1853 14519 1887
rect 14568 1884 14596 2051
rect 15654 2048 15660 2060
rect 15712 2048 15718 2100
rect 16666 2048 16672 2100
rect 16724 2048 16730 2100
rect 17954 2048 17960 2100
rect 18012 2088 18018 2100
rect 18141 2091 18199 2097
rect 18141 2088 18153 2091
rect 18012 2060 18153 2088
rect 18012 2048 18018 2060
rect 18141 2057 18153 2060
rect 18187 2057 18199 2091
rect 18141 2051 18199 2057
rect 18506 1912 18512 1964
rect 18564 1912 18570 1964
rect 15013 1897 15071 1903
rect 15013 1896 15025 1897
rect 15059 1896 15071 1897
rect 14737 1887 14795 1893
rect 14737 1884 14749 1887
rect 14568 1856 14749 1884
rect 14461 1847 14519 1853
rect 14737 1853 14749 1856
rect 14783 1853 14795 1887
rect 14737 1847 14795 1853
rect 14476 1816 14504 1847
rect 15010 1844 15016 1896
rect 15068 1894 15074 1896
rect 15068 1866 15103 1894
rect 15068 1844 15074 1866
rect 15286 1844 15292 1896
rect 15344 1884 15350 1896
rect 16482 1884 16488 1896
rect 15344 1856 16488 1884
rect 15344 1844 15350 1856
rect 16482 1844 16488 1856
rect 16540 1884 16546 1896
rect 16761 1887 16819 1893
rect 16761 1884 16773 1887
rect 16540 1856 16773 1884
rect 16540 1844 16546 1856
rect 16761 1853 16773 1856
rect 16807 1884 16819 1887
rect 18524 1884 18552 1912
rect 16807 1856 18552 1884
rect 16807 1853 16819 1856
rect 16761 1847 16819 1853
rect 19058 1844 19064 1896
rect 19116 1844 19122 1896
rect 15194 1816 15200 1828
rect 12176 1788 13216 1816
rect 13740 1788 14136 1816
rect 14200 1788 15200 1816
rect 12176 1760 12204 1788
rect 13188 1760 13216 1788
rect 7760 1720 8616 1748
rect 8849 1751 8907 1757
rect 8849 1717 8861 1751
rect 8895 1748 8907 1751
rect 10410 1748 10416 1760
rect 8895 1720 10416 1748
rect 8895 1717 8907 1720
rect 8849 1711 8907 1717
rect 10410 1708 10416 1720
rect 10468 1708 10474 1760
rect 10594 1708 10600 1760
rect 10652 1708 10658 1760
rect 12158 1708 12164 1760
rect 12216 1708 12222 1760
rect 13170 1708 13176 1760
rect 13228 1708 13234 1760
rect 13906 1708 13912 1760
rect 13964 1708 13970 1760
rect 14200 1757 14228 1788
rect 15194 1776 15200 1788
rect 15252 1776 15258 1828
rect 15556 1819 15614 1825
rect 15556 1785 15568 1819
rect 15602 1816 15614 1819
rect 15746 1816 15752 1828
rect 15602 1788 15752 1816
rect 15602 1785 15614 1788
rect 15556 1779 15614 1785
rect 15746 1776 15752 1788
rect 15804 1816 15810 1828
rect 15804 1788 16252 1816
rect 15804 1776 15810 1788
rect 16224 1760 16252 1788
rect 16298 1776 16304 1828
rect 16356 1816 16362 1828
rect 16574 1816 16580 1828
rect 16356 1788 16580 1816
rect 16356 1776 16362 1788
rect 16574 1776 16580 1788
rect 16632 1816 16638 1828
rect 17006 1819 17064 1825
rect 17006 1816 17018 1819
rect 16632 1788 17018 1816
rect 16632 1776 16638 1788
rect 17006 1785 17018 1788
rect 17052 1785 17064 1819
rect 17006 1779 17064 1785
rect 14185 1751 14243 1757
rect 14185 1717 14197 1751
rect 14231 1717 14243 1751
rect 14185 1711 14243 1717
rect 14829 1751 14887 1757
rect 14829 1717 14841 1751
rect 14875 1748 14887 1751
rect 15105 1751 15163 1757
rect 15105 1748 15117 1751
rect 14875 1720 15117 1748
rect 14875 1717 14887 1720
rect 14829 1711 14887 1717
rect 15105 1717 15117 1720
rect 15151 1748 15163 1751
rect 15654 1748 15660 1760
rect 15151 1720 15660 1748
rect 15151 1717 15163 1720
rect 15105 1711 15163 1717
rect 15654 1708 15660 1720
rect 15712 1708 15718 1760
rect 16206 1708 16212 1760
rect 16264 1708 16270 1760
rect 552 1658 19571 1680
rect 552 1606 5112 1658
rect 5164 1606 5176 1658
rect 5228 1606 5240 1658
rect 5292 1606 5304 1658
rect 5356 1606 5368 1658
rect 5420 1606 9827 1658
rect 9879 1606 9891 1658
rect 9943 1606 9955 1658
rect 10007 1606 10019 1658
rect 10071 1606 10083 1658
rect 10135 1606 14542 1658
rect 14594 1606 14606 1658
rect 14658 1606 14670 1658
rect 14722 1606 14734 1658
rect 14786 1606 14798 1658
rect 14850 1606 19257 1658
rect 19309 1606 19321 1658
rect 19373 1606 19385 1658
rect 19437 1606 19449 1658
rect 19501 1606 19513 1658
rect 19565 1606 19571 1658
rect 552 1584 19571 1606
rect 1394 1504 1400 1556
rect 1452 1504 1458 1556
rect 1486 1504 1492 1556
rect 1544 1504 1550 1556
rect 3053 1547 3111 1553
rect 3053 1513 3065 1547
rect 3099 1544 3111 1547
rect 4430 1544 4436 1556
rect 3099 1516 4436 1544
rect 3099 1513 3111 1516
rect 3053 1507 3111 1513
rect 4430 1504 4436 1516
rect 4488 1504 4494 1556
rect 4798 1504 4804 1556
rect 4856 1504 4862 1556
rect 4982 1504 4988 1556
rect 5040 1504 5046 1556
rect 5261 1547 5319 1553
rect 5261 1513 5273 1547
rect 5307 1544 5319 1547
rect 5534 1544 5540 1556
rect 5307 1516 5540 1544
rect 5307 1513 5319 1516
rect 5261 1507 5319 1513
rect 5534 1504 5540 1516
rect 5592 1544 5598 1556
rect 5592 1516 5764 1544
rect 5592 1504 5598 1516
rect 1412 1417 1440 1504
rect 1504 1476 1532 1504
rect 1918 1479 1976 1485
rect 1918 1476 1930 1479
rect 1504 1448 1930 1476
rect 1918 1445 1930 1448
rect 1964 1476 1976 1479
rect 2038 1476 2044 1488
rect 1964 1448 2044 1476
rect 1964 1445 1976 1448
rect 1918 1439 1976 1445
rect 2038 1436 2044 1448
rect 2096 1436 2102 1488
rect 3234 1436 3240 1488
rect 3292 1476 3298 1488
rect 3666 1479 3724 1485
rect 3666 1476 3678 1479
rect 3292 1448 3678 1476
rect 3292 1436 3298 1448
rect 3666 1445 3678 1448
rect 3712 1445 3724 1479
rect 3666 1439 3724 1445
rect 3878 1436 3884 1488
rect 3936 1436 3942 1488
rect 5000 1476 5028 1504
rect 5000 1448 5488 1476
rect 1397 1411 1455 1417
rect 1397 1377 1409 1411
rect 1443 1377 1455 1411
rect 2056 1408 2084 1436
rect 3145 1411 3203 1417
rect 3145 1408 3157 1411
rect 2056 1380 3157 1408
rect 1397 1371 1455 1377
rect 3145 1377 3157 1380
rect 3191 1377 3203 1411
rect 3145 1371 3203 1377
rect 1670 1300 1676 1352
rect 1728 1300 1734 1352
rect 3252 1349 3280 1436
rect 3896 1408 3924 1436
rect 3436 1380 3924 1408
rect 5077 1411 5135 1417
rect 3436 1349 3464 1380
rect 5077 1377 5089 1411
rect 5123 1377 5135 1411
rect 5077 1371 5135 1377
rect 3237 1343 3295 1349
rect 3237 1309 3249 1343
rect 3283 1309 3295 1343
rect 3237 1303 3295 1309
rect 3421 1343 3479 1349
rect 3421 1309 3433 1343
rect 3467 1309 3479 1343
rect 5092 1340 5120 1371
rect 5166 1368 5172 1420
rect 5224 1368 5230 1420
rect 5350 1408 5356 1420
rect 5267 1380 5356 1408
rect 5267 1340 5295 1380
rect 5350 1368 5356 1380
rect 5408 1368 5414 1420
rect 5460 1417 5488 1448
rect 5445 1411 5503 1417
rect 5445 1377 5457 1411
rect 5491 1377 5503 1411
rect 5736 1408 5764 1516
rect 5810 1504 5816 1556
rect 5868 1544 5874 1556
rect 5905 1547 5963 1553
rect 5905 1544 5917 1547
rect 5868 1516 5917 1544
rect 5868 1504 5874 1516
rect 5905 1513 5917 1516
rect 5951 1513 5963 1547
rect 5905 1507 5963 1513
rect 6457 1547 6515 1553
rect 6457 1513 6469 1547
rect 6503 1544 6515 1547
rect 6503 1516 7144 1544
rect 6503 1513 6515 1516
rect 6457 1507 6515 1513
rect 6181 1479 6239 1485
rect 6181 1445 6193 1479
rect 6227 1476 6239 1479
rect 6914 1476 6920 1488
rect 6227 1448 6920 1476
rect 6227 1445 6239 1448
rect 6181 1439 6239 1445
rect 6914 1436 6920 1448
rect 6972 1436 6978 1488
rect 5997 1411 6055 1417
rect 5997 1408 6009 1411
rect 5736 1380 6009 1408
rect 5445 1371 5503 1377
rect 5997 1377 6009 1380
rect 6043 1408 6055 1411
rect 6089 1411 6147 1417
rect 6089 1408 6101 1411
rect 6043 1380 6101 1408
rect 6043 1377 6055 1380
rect 5997 1371 6055 1377
rect 6089 1377 6101 1380
rect 6135 1377 6147 1411
rect 6089 1371 6147 1377
rect 6362 1368 6368 1420
rect 6420 1368 6426 1420
rect 6641 1411 6699 1417
rect 6641 1408 6653 1411
rect 6472 1380 6653 1408
rect 5092 1312 5295 1340
rect 5537 1343 5595 1349
rect 3421 1303 3479 1309
rect 5537 1309 5549 1343
rect 5583 1340 5595 1343
rect 6472 1340 6500 1380
rect 6641 1377 6653 1380
rect 6687 1377 6699 1411
rect 6641 1371 6699 1377
rect 6733 1411 6791 1417
rect 6733 1377 6745 1411
rect 6779 1408 6791 1411
rect 7006 1408 7012 1420
rect 6779 1380 7012 1408
rect 6779 1377 6791 1380
rect 6733 1371 6791 1377
rect 7006 1368 7012 1380
rect 7064 1368 7070 1420
rect 7116 1408 7144 1516
rect 8294 1504 8300 1556
rect 8352 1504 8358 1556
rect 8478 1504 8484 1556
rect 8536 1504 8542 1556
rect 8754 1504 8760 1556
rect 8812 1504 8818 1556
rect 9122 1504 9128 1556
rect 9180 1504 9186 1556
rect 9582 1504 9588 1556
rect 9640 1544 9646 1556
rect 9769 1547 9827 1553
rect 9769 1544 9781 1547
rect 9640 1516 9781 1544
rect 9640 1504 9646 1516
rect 9769 1513 9781 1516
rect 9815 1513 9827 1547
rect 9769 1507 9827 1513
rect 10410 1504 10416 1556
rect 10468 1544 10474 1556
rect 10468 1516 11008 1544
rect 10468 1504 10474 1516
rect 8496 1476 8524 1504
rect 8634 1479 8692 1485
rect 8634 1476 8646 1479
rect 8496 1448 8646 1476
rect 8634 1445 8646 1448
rect 8680 1445 8692 1479
rect 8634 1439 8692 1445
rect 7190 1417 7196 1420
rect 7184 1408 7196 1417
rect 7116 1380 7196 1408
rect 7184 1371 7196 1380
rect 7190 1368 7196 1371
rect 7248 1368 7254 1420
rect 8772 1408 8800 1504
rect 9140 1476 9168 1504
rect 9953 1479 10011 1485
rect 9953 1476 9965 1479
rect 9140 1448 9965 1476
rect 9953 1445 9965 1448
rect 9999 1476 10011 1479
rect 9999 1448 10640 1476
rect 9999 1445 10011 1448
rect 9953 1439 10011 1445
rect 10612 1420 10640 1448
rect 10045 1411 10103 1417
rect 10045 1408 10057 1411
rect 8772 1380 10057 1408
rect 10045 1377 10057 1380
rect 10091 1377 10103 1411
rect 10045 1371 10103 1377
rect 10318 1368 10324 1420
rect 10376 1408 10382 1420
rect 10505 1411 10563 1417
rect 10505 1408 10517 1411
rect 10376 1380 10517 1408
rect 10376 1368 10382 1380
rect 10505 1377 10517 1380
rect 10551 1377 10563 1411
rect 10505 1371 10563 1377
rect 5583 1312 6500 1340
rect 5583 1309 5595 1312
rect 5537 1303 5595 1309
rect 1688 1204 1716 1300
rect 2774 1232 2780 1284
rect 2832 1272 2838 1284
rect 3326 1272 3332 1284
rect 2832 1244 3332 1272
rect 2832 1232 2838 1244
rect 3326 1232 3332 1244
rect 3384 1232 3390 1284
rect 3436 1204 3464 1303
rect 6104 1284 6132 1312
rect 6546 1300 6552 1352
rect 6604 1340 6610 1352
rect 6917 1343 6975 1349
rect 6917 1340 6929 1343
rect 6604 1312 6929 1340
rect 6604 1300 6610 1312
rect 6917 1309 6929 1312
rect 6963 1309 6975 1343
rect 8386 1340 8392 1352
rect 6917 1303 6975 1309
rect 8220 1312 8392 1340
rect 6086 1232 6092 1284
rect 6144 1232 6150 1284
rect 1688 1176 3464 1204
rect 6932 1204 6960 1303
rect 8220 1204 8248 1312
rect 8386 1300 8392 1312
rect 8444 1300 8450 1352
rect 10520 1340 10548 1371
rect 10594 1368 10600 1420
rect 10652 1368 10658 1420
rect 10980 1417 11008 1516
rect 11054 1504 11060 1556
rect 11112 1504 11118 1556
rect 11330 1504 11336 1556
rect 11388 1504 11394 1556
rect 11422 1504 11428 1556
rect 11480 1544 11486 1556
rect 11885 1547 11943 1553
rect 11885 1544 11897 1547
rect 11480 1516 11897 1544
rect 11480 1504 11486 1516
rect 11885 1513 11897 1516
rect 11931 1544 11943 1547
rect 11931 1516 12480 1544
rect 11931 1513 11943 1516
rect 11885 1507 11943 1513
rect 11348 1476 11376 1504
rect 11348 1448 12388 1476
rect 10965 1411 11023 1417
rect 10965 1377 10977 1411
rect 11011 1398 11023 1411
rect 11011 1377 11100 1398
rect 10965 1371 11100 1377
rect 10980 1370 11100 1371
rect 10689 1343 10747 1349
rect 10689 1340 10701 1343
rect 10520 1312 10701 1340
rect 10689 1309 10701 1312
rect 10735 1309 10747 1343
rect 11072 1340 11100 1370
rect 11238 1368 11244 1420
rect 11296 1368 11302 1420
rect 11333 1411 11391 1417
rect 11333 1377 11345 1411
rect 11379 1408 11391 1411
rect 11422 1408 11428 1420
rect 11379 1380 11428 1408
rect 11379 1377 11391 1380
rect 11333 1371 11391 1377
rect 11422 1368 11428 1380
rect 11480 1368 11486 1420
rect 11992 1417 12020 1448
rect 11517 1411 11575 1417
rect 11517 1377 11529 1411
rect 11563 1377 11575 1411
rect 11517 1371 11575 1377
rect 11609 1411 11667 1417
rect 11609 1377 11621 1411
rect 11655 1408 11667 1411
rect 11977 1411 12035 1417
rect 11655 1380 11928 1408
rect 11655 1377 11667 1380
rect 11609 1371 11667 1377
rect 11532 1340 11560 1371
rect 11072 1312 11560 1340
rect 11900 1340 11928 1380
rect 11977 1377 11989 1411
rect 12023 1377 12035 1411
rect 12158 1408 12164 1420
rect 11977 1371 12035 1377
rect 12084 1380 12164 1408
rect 12084 1340 12112 1380
rect 12158 1368 12164 1380
rect 12216 1368 12222 1420
rect 12360 1417 12388 1448
rect 12253 1411 12311 1417
rect 12253 1377 12265 1411
rect 12299 1377 12311 1411
rect 12253 1371 12311 1377
rect 12345 1411 12403 1417
rect 12345 1377 12357 1411
rect 12391 1377 12403 1411
rect 12345 1371 12403 1377
rect 12452 1408 12480 1516
rect 12710 1504 12716 1556
rect 12768 1504 12774 1556
rect 13265 1547 13323 1553
rect 13265 1513 13277 1547
rect 13311 1544 13323 1547
rect 14182 1544 14188 1556
rect 13311 1516 14188 1544
rect 13311 1513 13323 1516
rect 13265 1507 13323 1513
rect 14182 1504 14188 1516
rect 14240 1504 14246 1556
rect 14829 1547 14887 1553
rect 14829 1513 14841 1547
rect 14875 1544 14887 1547
rect 14918 1544 14924 1556
rect 14875 1516 14924 1544
rect 14875 1513 14887 1516
rect 14829 1507 14887 1513
rect 14918 1504 14924 1516
rect 14976 1504 14982 1556
rect 15194 1504 15200 1556
rect 15252 1544 15258 1556
rect 15289 1547 15347 1553
rect 15289 1544 15301 1547
rect 15252 1516 15301 1544
rect 15252 1504 15258 1516
rect 15289 1513 15301 1516
rect 15335 1513 15347 1547
rect 15289 1507 15347 1513
rect 15565 1547 15623 1553
rect 15565 1513 15577 1547
rect 15611 1544 15623 1547
rect 16114 1544 16120 1556
rect 15611 1516 16120 1544
rect 15611 1513 15623 1516
rect 15565 1507 15623 1513
rect 12621 1411 12679 1417
rect 12621 1408 12633 1411
rect 12452 1380 12633 1408
rect 11900 1312 12112 1340
rect 12268 1340 12296 1371
rect 12452 1340 12480 1380
rect 12621 1377 12633 1380
rect 12667 1377 12679 1411
rect 12728 1408 12756 1504
rect 13906 1436 13912 1488
rect 13964 1476 13970 1488
rect 15010 1476 15016 1488
rect 13964 1448 15016 1476
rect 13964 1436 13970 1448
rect 12897 1411 12955 1417
rect 12897 1408 12909 1411
rect 12728 1380 12909 1408
rect 12621 1371 12679 1377
rect 12897 1377 12909 1380
rect 12943 1377 12955 1411
rect 12897 1371 12955 1377
rect 13170 1368 13176 1420
rect 13228 1368 13234 1420
rect 13446 1368 13452 1420
rect 13504 1368 13510 1420
rect 13538 1368 13544 1420
rect 13596 1408 13602 1420
rect 14936 1417 14964 1448
rect 15010 1436 15016 1448
rect 15068 1436 15074 1488
rect 15304 1476 15332 1507
rect 16114 1504 16120 1516
rect 16172 1504 16178 1556
rect 16206 1504 16212 1556
rect 16264 1504 16270 1556
rect 17865 1547 17923 1553
rect 17865 1513 17877 1547
rect 17911 1544 17923 1547
rect 18230 1544 18236 1556
rect 17911 1516 18236 1544
rect 17911 1513 17923 1516
rect 17865 1507 17923 1513
rect 18230 1504 18236 1516
rect 18288 1504 18294 1556
rect 15304 1448 15792 1476
rect 13705 1411 13763 1417
rect 13705 1408 13717 1411
rect 13596 1380 13717 1408
rect 13596 1368 13602 1380
rect 13705 1377 13717 1380
rect 13751 1377 13763 1411
rect 13705 1371 13763 1377
rect 14921 1411 14979 1417
rect 14921 1377 14933 1411
rect 14967 1377 14979 1411
rect 15381 1411 15439 1417
rect 15381 1408 15393 1411
rect 14921 1371 14979 1377
rect 15028 1380 15393 1408
rect 12268 1312 12480 1340
rect 12713 1343 12771 1349
rect 10689 1303 10747 1309
rect 12713 1309 12725 1343
rect 12759 1340 12771 1343
rect 13556 1340 13584 1368
rect 12759 1312 13584 1340
rect 12759 1309 12771 1312
rect 12713 1303 12771 1309
rect 6932 1176 8248 1204
rect 10704 1204 10732 1303
rect 12437 1275 12495 1281
rect 12437 1241 12449 1275
rect 12483 1272 12495 1275
rect 12989 1275 13047 1281
rect 12989 1272 13001 1275
rect 12483 1244 13001 1272
rect 12483 1241 12495 1244
rect 12437 1235 12495 1241
rect 12989 1241 13001 1244
rect 13035 1272 13047 1275
rect 13170 1272 13176 1284
rect 13035 1244 13176 1272
rect 13035 1241 13047 1244
rect 12989 1235 13047 1241
rect 13170 1232 13176 1244
rect 13228 1232 13234 1284
rect 11238 1204 11244 1216
rect 10704 1176 11244 1204
rect 11238 1164 11244 1176
rect 11296 1164 11302 1216
rect 14458 1164 14464 1216
rect 14516 1204 14522 1216
rect 15028 1213 15056 1380
rect 15381 1377 15393 1380
rect 15427 1408 15439 1411
rect 15427 1380 15608 1408
rect 15427 1377 15439 1380
rect 15381 1371 15439 1377
rect 15580 1272 15608 1380
rect 15654 1368 15660 1420
rect 15712 1368 15718 1420
rect 15764 1417 15792 1448
rect 15749 1411 15807 1417
rect 15749 1377 15761 1411
rect 15795 1377 15807 1411
rect 15749 1371 15807 1377
rect 15841 1411 15899 1417
rect 15841 1377 15853 1411
rect 15887 1408 15899 1411
rect 16301 1411 16359 1417
rect 16301 1408 16313 1411
rect 15887 1380 16313 1408
rect 15887 1377 15899 1380
rect 15841 1371 15899 1377
rect 16301 1377 16313 1380
rect 16347 1408 16359 1411
rect 16390 1408 16396 1420
rect 16347 1380 16396 1408
rect 16347 1377 16359 1380
rect 16301 1371 16359 1377
rect 16390 1368 16396 1380
rect 16448 1368 16454 1420
rect 16482 1368 16488 1420
rect 16540 1368 16546 1420
rect 16574 1368 16580 1420
rect 16632 1408 16638 1420
rect 16741 1411 16799 1417
rect 16741 1408 16753 1411
rect 16632 1380 16753 1408
rect 16632 1368 16638 1380
rect 16741 1377 16753 1380
rect 16787 1377 16799 1411
rect 16741 1371 16799 1377
rect 15672 1340 15700 1368
rect 16114 1340 16120 1352
rect 15672 1312 16120 1340
rect 16114 1300 16120 1312
rect 16172 1300 16178 1352
rect 16592 1340 16620 1368
rect 16500 1312 16620 1340
rect 16500 1272 16528 1312
rect 15580 1244 16528 1272
rect 15013 1207 15071 1213
rect 15013 1204 15025 1207
rect 14516 1176 15025 1204
rect 14516 1164 14522 1176
rect 15013 1173 15025 1176
rect 15059 1173 15071 1207
rect 15013 1167 15071 1173
rect 552 1114 19412 1136
rect 552 1062 2755 1114
rect 2807 1062 2819 1114
rect 2871 1062 2883 1114
rect 2935 1062 2947 1114
rect 2999 1062 3011 1114
rect 3063 1062 7470 1114
rect 7522 1062 7534 1114
rect 7586 1062 7598 1114
rect 7650 1062 7662 1114
rect 7714 1062 7726 1114
rect 7778 1062 12185 1114
rect 12237 1062 12249 1114
rect 12301 1062 12313 1114
rect 12365 1062 12377 1114
rect 12429 1062 12441 1114
rect 12493 1062 16900 1114
rect 16952 1062 16964 1114
rect 17016 1062 17028 1114
rect 17080 1062 17092 1114
rect 17144 1062 17156 1114
rect 17208 1062 19412 1114
rect 552 1040 19412 1062
rect 2222 960 2228 1012
rect 2280 960 2286 1012
rect 4157 1003 4215 1009
rect 4157 969 4169 1003
rect 4203 1000 4215 1003
rect 4890 1000 4896 1012
rect 4203 972 4896 1000
rect 4203 969 4215 972
rect 4157 963 4215 969
rect 4890 960 4896 972
rect 4948 960 4954 1012
rect 7190 960 7196 1012
rect 7248 960 7254 1012
rect 10597 1003 10655 1009
rect 10597 969 10609 1003
rect 10643 1000 10655 1003
rect 11146 1000 11152 1012
rect 10643 972 11152 1000
rect 10643 969 10655 972
rect 10597 963 10655 969
rect 11146 960 11152 972
rect 11204 960 11210 1012
rect 11882 960 11888 1012
rect 11940 1000 11946 1012
rect 13173 1003 13231 1009
rect 13173 1000 13185 1003
rect 11940 972 13185 1000
rect 11940 960 11946 972
rect 13173 969 13185 972
rect 13219 969 13231 1003
rect 13173 963 13231 969
rect 13538 960 13544 1012
rect 13596 1000 13602 1012
rect 13633 1003 13691 1009
rect 13633 1000 13645 1003
rect 13596 972 13645 1000
rect 13596 960 13602 972
rect 13633 969 13645 972
rect 13679 969 13691 1003
rect 13633 963 13691 969
rect 1946 892 1952 944
rect 2004 932 2010 944
rect 2409 935 2467 941
rect 2409 932 2421 935
rect 2004 904 2421 932
rect 2004 892 2010 904
rect 2409 901 2421 904
rect 2455 901 2467 935
rect 2409 895 2467 901
rect 11790 892 11796 944
rect 11848 932 11854 944
rect 11977 935 12035 941
rect 11977 932 11989 935
rect 11848 904 11989 932
rect 11848 892 11854 904
rect 11977 901 11989 904
rect 12023 901 12035 935
rect 11977 895 12035 901
rect 12894 892 12900 944
rect 12952 892 12958 944
rect 2038 824 2044 876
rect 2096 864 2102 876
rect 13648 864 13676 963
rect 13906 960 13912 1012
rect 13964 960 13970 1012
rect 14182 960 14188 1012
rect 14240 960 14246 1012
rect 14458 960 14464 1012
rect 14516 960 14522 1012
rect 15657 1003 15715 1009
rect 15657 969 15669 1003
rect 15703 1000 15715 1003
rect 15930 1000 15936 1012
rect 15703 972 15936 1000
rect 15703 969 15715 972
rect 15657 963 15715 969
rect 15930 960 15936 972
rect 15988 960 15994 1012
rect 16209 1003 16267 1009
rect 16209 969 16221 1003
rect 16255 1000 16267 1003
rect 16298 1000 16304 1012
rect 16255 972 16304 1000
rect 16255 969 16267 972
rect 16209 963 16267 969
rect 16298 960 16304 972
rect 16356 1000 16362 1012
rect 16485 1003 16543 1009
rect 16485 1000 16497 1003
rect 16356 972 16497 1000
rect 16356 960 16362 972
rect 16485 969 16497 972
rect 16531 969 16543 1003
rect 16485 963 16543 969
rect 2096 836 2360 864
rect 13648 836 14320 864
rect 2096 824 2102 836
rect 842 756 848 808
rect 900 756 906 808
rect 1302 756 1308 808
rect 1360 796 1366 808
rect 2332 805 2360 836
rect 1397 799 1455 805
rect 1397 796 1409 799
rect 1360 768 1409 796
rect 1360 756 1366 768
rect 1397 765 1409 768
rect 1443 765 1455 799
rect 1397 759 1455 765
rect 2317 799 2375 805
rect 2317 765 2329 799
rect 2363 765 2375 799
rect 2317 759 2375 765
rect 3602 756 3608 808
rect 3660 796 3666 808
rect 4065 799 4123 805
rect 4065 796 4077 799
rect 3660 768 4077 796
rect 3660 756 3666 768
rect 4065 765 4077 768
rect 4111 765 4123 799
rect 4065 759 4123 765
rect 6914 756 6920 808
rect 6972 796 6978 808
rect 7285 799 7343 805
rect 7285 796 7297 799
rect 6972 768 7297 796
rect 6972 756 6978 768
rect 7285 765 7297 768
rect 7331 765 7343 799
rect 7285 759 7343 765
rect 10410 756 10416 808
rect 10468 756 10474 808
rect 13170 756 13176 808
rect 13228 796 13234 808
rect 14292 805 14320 836
rect 13725 799 13783 805
rect 13725 796 13737 799
rect 13228 768 13737 796
rect 13228 756 13234 768
rect 13725 765 13737 768
rect 13771 796 13783 799
rect 13817 799 13875 805
rect 13817 796 13829 799
rect 13771 768 13829 796
rect 13771 765 13783 768
rect 13725 759 13783 765
rect 13817 765 13829 768
rect 13863 765 13875 799
rect 13817 759 13875 765
rect 14277 799 14335 805
rect 14277 765 14289 799
rect 14323 796 14335 799
rect 14369 799 14427 805
rect 14369 796 14381 799
rect 14323 768 14381 796
rect 14323 765 14335 768
rect 14277 759 14335 765
rect 14369 765 14381 768
rect 14415 765 14427 799
rect 14369 759 14427 765
rect 15749 799 15807 805
rect 15749 765 15761 799
rect 15795 765 15807 799
rect 15749 759 15807 765
rect 11790 688 11796 740
rect 11848 688 11854 740
rect 12250 688 12256 740
rect 12308 728 12314 740
rect 12713 731 12771 737
rect 12713 728 12725 731
rect 12308 700 12725 728
rect 12308 688 12314 700
rect 12713 697 12725 700
rect 12759 697 12771 731
rect 12713 691 12771 697
rect 13078 688 13084 740
rect 13136 688 13142 740
rect 15764 728 15792 759
rect 16114 756 16120 808
rect 16172 756 16178 808
rect 16298 756 16304 808
rect 16356 756 16362 808
rect 16574 756 16580 808
rect 16632 756 16638 808
rect 18506 756 18512 808
rect 18564 756 18570 808
rect 19058 756 19064 808
rect 19116 756 19122 808
rect 16316 728 16344 756
rect 15764 700 16344 728
rect 552 570 19571 592
rect 552 518 5112 570
rect 5164 518 5176 570
rect 5228 518 5240 570
rect 5292 518 5304 570
rect 5356 518 5368 570
rect 5420 518 9827 570
rect 9879 518 9891 570
rect 9943 518 9955 570
rect 10007 518 10019 570
rect 10071 518 10083 570
rect 10135 518 14542 570
rect 14594 518 14606 570
rect 14658 518 14670 570
rect 14722 518 14734 570
rect 14786 518 14798 570
rect 14850 518 19257 570
rect 19309 518 19321 570
rect 19373 518 19385 570
rect 19437 518 19449 570
rect 19501 518 19513 570
rect 19565 518 19571 570
rect 552 496 19571 518
<< via1 >>
rect 5112 19014 5164 19066
rect 5176 19014 5228 19066
rect 5240 19014 5292 19066
rect 5304 19014 5356 19066
rect 5368 19014 5420 19066
rect 9827 19014 9879 19066
rect 9891 19014 9943 19066
rect 9955 19014 10007 19066
rect 10019 19014 10071 19066
rect 10083 19014 10135 19066
rect 14542 19014 14594 19066
rect 14606 19014 14658 19066
rect 14670 19014 14722 19066
rect 14734 19014 14786 19066
rect 14798 19014 14850 19066
rect 19257 19014 19309 19066
rect 19321 19014 19373 19066
rect 19385 19014 19437 19066
rect 19449 19014 19501 19066
rect 19513 19014 19565 19066
rect 13544 18912 13596 18964
rect 15384 18912 15436 18964
rect 10416 18844 10468 18896
rect 756 18776 808 18828
rect 1124 18751 1176 18760
rect 1124 18717 1133 18751
rect 1133 18717 1167 18751
rect 1167 18717 1176 18751
rect 1124 18708 1176 18717
rect 11980 18776 12032 18828
rect 12992 18819 13044 18828
rect 12992 18785 13001 18819
rect 13001 18785 13035 18819
rect 13035 18785 13044 18819
rect 12992 18776 13044 18785
rect 848 18615 900 18624
rect 848 18581 857 18615
rect 857 18581 891 18615
rect 891 18581 900 18615
rect 848 18572 900 18581
rect 11428 18572 11480 18624
rect 12532 18572 12584 18624
rect 14004 18708 14056 18760
rect 14188 18776 14240 18828
rect 18512 18819 18564 18828
rect 18512 18785 18521 18819
rect 18521 18785 18555 18819
rect 18555 18785 18564 18819
rect 18512 18776 18564 18785
rect 13912 18615 13964 18624
rect 13912 18581 13921 18615
rect 13921 18581 13955 18615
rect 13955 18581 13964 18615
rect 13912 18572 13964 18581
rect 14372 18572 14424 18624
rect 19064 18615 19116 18624
rect 19064 18581 19073 18615
rect 19073 18581 19107 18615
rect 19107 18581 19116 18615
rect 19064 18572 19116 18581
rect 2755 18470 2807 18522
rect 2819 18470 2871 18522
rect 2883 18470 2935 18522
rect 2947 18470 2999 18522
rect 3011 18470 3063 18522
rect 7470 18470 7522 18522
rect 7534 18470 7586 18522
rect 7598 18470 7650 18522
rect 7662 18470 7714 18522
rect 7726 18470 7778 18522
rect 12185 18470 12237 18522
rect 12249 18470 12301 18522
rect 12313 18470 12365 18522
rect 12377 18470 12429 18522
rect 12441 18470 12493 18522
rect 16900 18470 16952 18522
rect 16964 18470 17016 18522
rect 17028 18470 17080 18522
rect 17092 18470 17144 18522
rect 17156 18470 17208 18522
rect 10416 18411 10468 18420
rect 10416 18377 10425 18411
rect 10425 18377 10459 18411
rect 10459 18377 10468 18411
rect 10416 18368 10468 18377
rect 10508 18368 10560 18420
rect 11428 18368 11480 18420
rect 12532 18411 12584 18420
rect 12532 18377 12541 18411
rect 12541 18377 12575 18411
rect 12575 18377 12584 18411
rect 12532 18368 12584 18377
rect 2412 18232 2464 18284
rect 848 18207 900 18216
rect 848 18173 857 18207
rect 857 18173 891 18207
rect 891 18173 900 18207
rect 848 18164 900 18173
rect 2688 18207 2740 18216
rect 2688 18173 2697 18207
rect 2697 18173 2731 18207
rect 2731 18173 2740 18207
rect 2688 18164 2740 18173
rect 3792 18096 3844 18148
rect 4160 18096 4212 18148
rect 2596 18071 2648 18080
rect 2596 18037 2605 18071
rect 2605 18037 2639 18071
rect 2639 18037 2648 18071
rect 2596 18028 2648 18037
rect 5724 18028 5776 18080
rect 6092 18071 6144 18080
rect 6092 18037 6101 18071
rect 6101 18037 6135 18071
rect 6135 18037 6144 18071
rect 6092 18028 6144 18037
rect 6276 18028 6328 18080
rect 8392 18164 8444 18216
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 8484 18096 8536 18148
rect 11796 18207 11848 18216
rect 11796 18173 11805 18207
rect 11805 18173 11839 18207
rect 11839 18173 11848 18207
rect 11796 18164 11848 18173
rect 14464 18164 14516 18216
rect 15292 18164 15344 18216
rect 18052 18207 18104 18216
rect 13912 18096 13964 18148
rect 14832 18139 14884 18148
rect 14832 18105 14861 18139
rect 14861 18105 14884 18139
rect 14832 18096 14884 18105
rect 9588 18028 9640 18080
rect 10140 18028 10192 18080
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 10692 18028 10744 18080
rect 11336 18028 11388 18080
rect 12992 18028 13044 18080
rect 13360 18028 13412 18080
rect 13728 18071 13780 18080
rect 13728 18037 13737 18071
rect 13737 18037 13771 18071
rect 13771 18037 13780 18071
rect 13728 18028 13780 18037
rect 15384 18096 15436 18148
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 19064 18207 19116 18216
rect 19064 18173 19073 18207
rect 19073 18173 19107 18207
rect 19107 18173 19116 18207
rect 19064 18164 19116 18173
rect 18236 18096 18288 18148
rect 16580 18071 16632 18080
rect 16580 18037 16589 18071
rect 16589 18037 16623 18071
rect 16623 18037 16632 18071
rect 16580 18028 16632 18037
rect 16672 18071 16724 18080
rect 16672 18037 16681 18071
rect 16681 18037 16715 18071
rect 16715 18037 16724 18071
rect 16672 18028 16724 18037
rect 5112 17926 5164 17978
rect 5176 17926 5228 17978
rect 5240 17926 5292 17978
rect 5304 17926 5356 17978
rect 5368 17926 5420 17978
rect 9827 17926 9879 17978
rect 9891 17926 9943 17978
rect 9955 17926 10007 17978
rect 10019 17926 10071 17978
rect 10083 17926 10135 17978
rect 14542 17926 14594 17978
rect 14606 17926 14658 17978
rect 14670 17926 14722 17978
rect 14734 17926 14786 17978
rect 14798 17926 14850 17978
rect 19257 17926 19309 17978
rect 19321 17926 19373 17978
rect 19385 17926 19437 17978
rect 19449 17926 19501 17978
rect 19513 17926 19565 17978
rect 4344 17824 4396 17876
rect 9864 17824 9916 17876
rect 2596 17756 2648 17808
rect 2320 17731 2372 17740
rect 2320 17697 2329 17731
rect 2329 17697 2363 17731
rect 2363 17697 2372 17731
rect 2320 17688 2372 17697
rect 4160 17731 4212 17740
rect 4160 17697 4169 17731
rect 4169 17697 4203 17731
rect 4203 17697 4212 17731
rect 4160 17688 4212 17697
rect 6276 17756 6328 17808
rect 9404 17756 9456 17808
rect 4436 17731 4488 17740
rect 4436 17697 4470 17731
rect 4470 17697 4488 17731
rect 4436 17688 4488 17697
rect 1492 17620 1544 17672
rect 1584 17620 1636 17672
rect 2412 17663 2464 17672
rect 2412 17629 2421 17663
rect 2421 17629 2455 17663
rect 2455 17629 2464 17663
rect 2412 17620 2464 17629
rect 6552 17731 6604 17740
rect 6552 17697 6561 17731
rect 6561 17697 6595 17731
rect 6595 17697 6604 17731
rect 6552 17688 6604 17697
rect 8116 17688 8168 17740
rect 8392 17688 8444 17740
rect 9680 17688 9732 17740
rect 10232 17756 10284 17808
rect 11244 17824 11296 17876
rect 13728 17824 13780 17876
rect 13912 17824 13964 17876
rect 18236 17824 18288 17876
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 1860 17484 1912 17536
rect 2228 17527 2280 17536
rect 2228 17493 2237 17527
rect 2237 17493 2271 17527
rect 2271 17493 2280 17527
rect 2228 17484 2280 17493
rect 4068 17484 4120 17536
rect 6276 17552 6328 17604
rect 6736 17527 6788 17536
rect 6736 17493 6745 17527
rect 6745 17493 6779 17527
rect 6779 17493 6788 17527
rect 6736 17484 6788 17493
rect 6828 17527 6880 17536
rect 6828 17493 6837 17527
rect 6837 17493 6871 17527
rect 6871 17493 6880 17527
rect 6828 17484 6880 17493
rect 10324 17552 10376 17604
rect 9772 17527 9824 17536
rect 9772 17493 9781 17527
rect 9781 17493 9815 17527
rect 9815 17493 9824 17527
rect 9772 17484 9824 17493
rect 9864 17484 9916 17536
rect 11152 17731 11204 17740
rect 11152 17697 11161 17731
rect 11161 17697 11195 17731
rect 11195 17697 11204 17731
rect 11152 17688 11204 17697
rect 11244 17731 11296 17740
rect 11244 17697 11253 17731
rect 11253 17697 11287 17731
rect 11287 17697 11296 17731
rect 11244 17688 11296 17697
rect 18052 17756 18104 17808
rect 11888 17688 11940 17740
rect 12532 17688 12584 17740
rect 13360 17731 13412 17740
rect 13360 17697 13369 17731
rect 13369 17697 13403 17731
rect 13403 17697 13412 17731
rect 13360 17688 13412 17697
rect 13728 17731 13780 17740
rect 13728 17697 13737 17731
rect 13737 17697 13771 17731
rect 13771 17697 13780 17731
rect 13728 17688 13780 17697
rect 14004 17731 14056 17740
rect 14004 17697 14013 17731
rect 14013 17697 14047 17731
rect 14047 17697 14056 17731
rect 14004 17688 14056 17697
rect 14280 17731 14332 17740
rect 14280 17697 14289 17731
rect 14289 17697 14323 17731
rect 14323 17697 14332 17731
rect 14280 17688 14332 17697
rect 14372 17688 14424 17740
rect 15108 17688 15160 17740
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 14464 17620 14516 17672
rect 16580 17688 16632 17740
rect 18788 17688 18840 17740
rect 11428 17552 11480 17604
rect 14188 17552 14240 17604
rect 10692 17527 10744 17536
rect 10692 17493 10701 17527
rect 10701 17493 10735 17527
rect 10735 17493 10744 17527
rect 10692 17484 10744 17493
rect 11520 17527 11572 17536
rect 11520 17493 11529 17527
rect 11529 17493 11563 17527
rect 11563 17493 11572 17527
rect 11520 17484 11572 17493
rect 12900 17484 12952 17536
rect 14556 17484 14608 17536
rect 16304 17552 16356 17604
rect 16672 17552 16724 17604
rect 16120 17527 16172 17536
rect 16120 17493 16129 17527
rect 16129 17493 16163 17527
rect 16163 17493 16172 17527
rect 16120 17484 16172 17493
rect 16764 17484 16816 17536
rect 17224 17484 17276 17536
rect 18696 17527 18748 17536
rect 18696 17493 18705 17527
rect 18705 17493 18739 17527
rect 18739 17493 18748 17527
rect 18696 17484 18748 17493
rect 2755 17382 2807 17434
rect 2819 17382 2871 17434
rect 2883 17382 2935 17434
rect 2947 17382 2999 17434
rect 3011 17382 3063 17434
rect 7470 17382 7522 17434
rect 7534 17382 7586 17434
rect 7598 17382 7650 17434
rect 7662 17382 7714 17434
rect 7726 17382 7778 17434
rect 12185 17382 12237 17434
rect 12249 17382 12301 17434
rect 12313 17382 12365 17434
rect 12377 17382 12429 17434
rect 12441 17382 12493 17434
rect 16900 17382 16952 17434
rect 16964 17382 17016 17434
rect 17028 17382 17080 17434
rect 17092 17382 17144 17434
rect 17156 17382 17208 17434
rect 2228 17280 2280 17332
rect 4344 17280 4396 17332
rect 4436 17280 4488 17332
rect 6828 17280 6880 17332
rect 8484 17323 8536 17332
rect 8484 17289 8493 17323
rect 8493 17289 8527 17323
rect 8527 17289 8536 17323
rect 8484 17280 8536 17289
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 9588 17323 9640 17332
rect 9588 17289 9597 17323
rect 9597 17289 9631 17323
rect 9631 17289 9640 17323
rect 9588 17280 9640 17289
rect 10140 17280 10192 17332
rect 11152 17280 11204 17332
rect 11428 17323 11480 17332
rect 11428 17289 11437 17323
rect 11437 17289 11471 17323
rect 11471 17289 11480 17323
rect 11428 17280 11480 17289
rect 11796 17280 11848 17332
rect 11980 17323 12032 17332
rect 11980 17289 11989 17323
rect 11989 17289 12023 17323
rect 12023 17289 12032 17323
rect 11980 17280 12032 17289
rect 13728 17280 13780 17332
rect 14280 17280 14332 17332
rect 14556 17280 14608 17332
rect 15108 17280 15160 17332
rect 1584 17187 1636 17196
rect 1584 17153 1593 17187
rect 1593 17153 1627 17187
rect 1627 17153 1636 17187
rect 1584 17144 1636 17153
rect 848 17119 900 17128
rect 848 17085 857 17119
rect 857 17085 891 17119
rect 891 17085 900 17119
rect 848 17076 900 17085
rect 1492 17119 1544 17128
rect 1492 17085 1501 17119
rect 1501 17085 1535 17119
rect 1535 17085 1544 17119
rect 1492 17076 1544 17085
rect 1860 17119 1912 17128
rect 1860 17085 1894 17119
rect 1894 17085 1912 17119
rect 1860 17076 1912 17085
rect 4160 17144 4212 17196
rect 2320 16940 2372 16992
rect 3148 17008 3200 17060
rect 4252 17076 4304 17128
rect 4344 17119 4396 17128
rect 4344 17085 4353 17119
rect 4353 17085 4387 17119
rect 4387 17085 4396 17119
rect 4344 17076 4396 17085
rect 3884 17008 3936 17060
rect 4804 17119 4856 17128
rect 4804 17085 4813 17119
rect 4813 17085 4847 17119
rect 4847 17085 4856 17119
rect 4804 17076 4856 17085
rect 4988 17008 5040 17060
rect 3700 16983 3752 16992
rect 3700 16949 3709 16983
rect 3709 16949 3743 16983
rect 3743 16949 3752 16983
rect 3700 16940 3752 16949
rect 3792 16940 3844 16992
rect 4068 16940 4120 16992
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 7932 17076 7984 17085
rect 8116 17076 8168 17128
rect 9312 17144 9364 17196
rect 7748 17051 7800 17060
rect 7748 17017 7757 17051
rect 7757 17017 7791 17051
rect 7791 17017 7800 17051
rect 9496 17076 9548 17128
rect 9588 17076 9640 17128
rect 10692 17119 10744 17128
rect 10692 17085 10701 17119
rect 10701 17085 10735 17119
rect 10735 17085 10744 17119
rect 10692 17076 10744 17085
rect 10876 17076 10928 17128
rect 11612 17144 11664 17196
rect 7748 17008 7800 17017
rect 8116 16983 8168 16992
rect 8116 16949 8125 16983
rect 8125 16949 8159 16983
rect 8159 16949 8168 16983
rect 8116 16940 8168 16949
rect 11060 17008 11112 17060
rect 11428 17076 11480 17128
rect 14188 17212 14240 17264
rect 13544 17144 13596 17196
rect 13912 17144 13964 17196
rect 15108 17144 15160 17196
rect 14924 17076 14976 17128
rect 15568 17280 15620 17332
rect 16764 17280 16816 17332
rect 18696 17280 18748 17332
rect 18788 17323 18840 17332
rect 18788 17289 18797 17323
rect 18797 17289 18831 17323
rect 18831 17289 18840 17323
rect 18788 17280 18840 17289
rect 15384 17119 15436 17128
rect 15384 17085 15393 17119
rect 15393 17085 15427 17119
rect 15427 17085 15436 17119
rect 15384 17076 15436 17085
rect 16764 17119 16816 17128
rect 16764 17085 16773 17119
rect 16773 17085 16807 17119
rect 16807 17085 16816 17119
rect 16764 17076 16816 17085
rect 9312 16940 9364 16992
rect 11888 16940 11940 16992
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 15200 16940 15252 16992
rect 16672 16940 16724 16992
rect 16948 16940 17000 16992
rect 17316 17008 17368 17060
rect 17776 17119 17828 17128
rect 17776 17085 17785 17119
rect 17785 17085 17819 17119
rect 17819 17085 17828 17119
rect 17776 17076 17828 17085
rect 17960 17076 18012 17128
rect 18696 17121 18748 17128
rect 18696 17087 18705 17121
rect 18705 17087 18739 17121
rect 18739 17087 18748 17121
rect 18696 17076 18748 17087
rect 17868 16940 17920 16992
rect 18236 16983 18288 16992
rect 18236 16949 18245 16983
rect 18245 16949 18279 16983
rect 18279 16949 18288 16983
rect 18236 16940 18288 16949
rect 5112 16838 5164 16890
rect 5176 16838 5228 16890
rect 5240 16838 5292 16890
rect 5304 16838 5356 16890
rect 5368 16838 5420 16890
rect 9827 16838 9879 16890
rect 9891 16838 9943 16890
rect 9955 16838 10007 16890
rect 10019 16838 10071 16890
rect 10083 16838 10135 16890
rect 14542 16838 14594 16890
rect 14606 16838 14658 16890
rect 14670 16838 14722 16890
rect 14734 16838 14786 16890
rect 14798 16838 14850 16890
rect 19257 16838 19309 16890
rect 19321 16838 19373 16890
rect 19385 16838 19437 16890
rect 19449 16838 19501 16890
rect 19513 16838 19565 16890
rect 1400 16736 1452 16788
rect 1860 16736 1912 16788
rect 2228 16736 2280 16788
rect 2320 16736 2372 16788
rect 2780 16736 2832 16788
rect 3148 16736 3200 16788
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 2596 16668 2648 16720
rect 1860 16439 1912 16448
rect 1860 16405 1869 16439
rect 1869 16405 1903 16439
rect 1903 16405 1912 16439
rect 1860 16396 1912 16405
rect 2412 16396 2464 16448
rect 3700 16736 3752 16788
rect 3884 16736 3936 16788
rect 4804 16736 4856 16788
rect 4988 16736 5040 16788
rect 6092 16736 6144 16788
rect 4344 16668 4396 16720
rect 3240 16532 3292 16584
rect 4068 16600 4120 16652
rect 4988 16643 5040 16652
rect 4988 16609 4997 16643
rect 4997 16609 5031 16643
rect 5031 16609 5040 16643
rect 4988 16600 5040 16609
rect 5540 16600 5592 16652
rect 5724 16600 5776 16652
rect 6000 16643 6052 16652
rect 6000 16609 6017 16643
rect 6017 16609 6051 16643
rect 6051 16609 6052 16643
rect 6000 16600 6052 16609
rect 6276 16643 6328 16652
rect 6276 16609 6285 16643
rect 6285 16609 6319 16643
rect 6319 16609 6328 16643
rect 6276 16600 6328 16609
rect 6552 16736 6604 16788
rect 7932 16736 7984 16788
rect 10784 16736 10836 16788
rect 10876 16736 10928 16788
rect 11060 16779 11112 16788
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 11612 16779 11664 16788
rect 11612 16745 11621 16779
rect 11621 16745 11655 16779
rect 11655 16745 11664 16779
rect 11612 16736 11664 16745
rect 7748 16600 7800 16652
rect 5908 16575 5960 16584
rect 4252 16464 4304 16516
rect 5908 16541 5917 16575
rect 5917 16541 5951 16575
rect 5951 16541 5960 16575
rect 5908 16532 5960 16541
rect 3792 16396 3844 16448
rect 6644 16439 6696 16448
rect 6644 16405 6653 16439
rect 6653 16405 6687 16439
rect 6687 16405 6696 16439
rect 6644 16396 6696 16405
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 8208 16600 8260 16652
rect 13912 16668 13964 16720
rect 14648 16668 14700 16720
rect 11428 16643 11480 16652
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 11612 16532 11664 16584
rect 11060 16464 11112 16516
rect 11980 16643 12032 16652
rect 11980 16609 11989 16643
rect 11989 16609 12023 16643
rect 12023 16609 12032 16643
rect 11980 16600 12032 16609
rect 14096 16643 14148 16652
rect 14096 16609 14105 16643
rect 14105 16609 14139 16643
rect 14139 16609 14148 16643
rect 14924 16736 14976 16788
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 16948 16779 17000 16788
rect 16948 16745 16957 16779
rect 16957 16745 16991 16779
rect 16991 16745 17000 16779
rect 16948 16736 17000 16745
rect 18236 16736 18288 16788
rect 14832 16668 14884 16720
rect 15568 16668 15620 16720
rect 14096 16600 14148 16609
rect 15016 16643 15068 16652
rect 15016 16609 15025 16643
rect 15025 16609 15059 16643
rect 15059 16609 15068 16643
rect 15016 16600 15068 16609
rect 15108 16643 15160 16652
rect 15108 16609 15117 16643
rect 15117 16609 15151 16643
rect 15151 16609 15160 16643
rect 15108 16600 15160 16609
rect 18052 16668 18104 16720
rect 17500 16600 17552 16652
rect 17868 16600 17920 16652
rect 18604 16643 18656 16652
rect 18604 16609 18613 16643
rect 18613 16609 18647 16643
rect 18647 16609 18656 16643
rect 18604 16600 18656 16609
rect 19064 16643 19116 16652
rect 19064 16609 19073 16643
rect 19073 16609 19107 16643
rect 19107 16609 19116 16643
rect 19064 16600 19116 16609
rect 17224 16532 17276 16584
rect 13176 16464 13228 16516
rect 17316 16464 17368 16516
rect 8392 16396 8444 16448
rect 11152 16396 11204 16448
rect 11888 16396 11940 16448
rect 14004 16439 14056 16448
rect 14004 16405 14013 16439
rect 14013 16405 14047 16439
rect 14047 16405 14056 16439
rect 14004 16396 14056 16405
rect 14280 16396 14332 16448
rect 14832 16396 14884 16448
rect 15108 16396 15160 16448
rect 17224 16396 17276 16448
rect 18696 16439 18748 16448
rect 18696 16405 18705 16439
rect 18705 16405 18739 16439
rect 18739 16405 18748 16439
rect 18696 16396 18748 16405
rect 2755 16294 2807 16346
rect 2819 16294 2871 16346
rect 2883 16294 2935 16346
rect 2947 16294 2999 16346
rect 3011 16294 3063 16346
rect 7470 16294 7522 16346
rect 7534 16294 7586 16346
rect 7598 16294 7650 16346
rect 7662 16294 7714 16346
rect 7726 16294 7778 16346
rect 12185 16294 12237 16346
rect 12249 16294 12301 16346
rect 12313 16294 12365 16346
rect 12377 16294 12429 16346
rect 12441 16294 12493 16346
rect 16900 16294 16952 16346
rect 16964 16294 17016 16346
rect 17028 16294 17080 16346
rect 17092 16294 17144 16346
rect 17156 16294 17208 16346
rect 4988 16192 5040 16244
rect 5540 16192 5592 16244
rect 1584 16124 1636 16176
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 1860 16031 1912 16040
rect 1860 15997 1869 16031
rect 1869 15997 1903 16031
rect 1903 15997 1912 16031
rect 1860 15988 1912 15997
rect 2504 16056 2556 16108
rect 5908 16192 5960 16244
rect 3240 16031 3292 16040
rect 3240 15997 3249 16031
rect 3249 15997 3283 16031
rect 3283 15997 3292 16031
rect 3240 15988 3292 15997
rect 3608 15988 3660 16040
rect 6000 16056 6052 16108
rect 8208 16192 8260 16244
rect 9312 16192 9364 16244
rect 3516 15920 3568 15972
rect 6828 15920 6880 15972
rect 7564 15920 7616 15972
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 11152 16192 11204 16244
rect 14004 16192 14056 16244
rect 15292 16192 15344 16244
rect 11336 16124 11388 16176
rect 11520 16124 11572 16176
rect 17500 16192 17552 16244
rect 9128 15920 9180 15972
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 11152 16031 11204 16040
rect 11152 15997 11161 16031
rect 11161 15997 11195 16031
rect 11195 15997 11204 16031
rect 11152 15988 11204 15997
rect 11612 15988 11664 16040
rect 12348 15988 12400 16040
rect 13176 15988 13228 16040
rect 13912 16031 13964 16040
rect 13912 15997 13921 16031
rect 13921 15997 13955 16031
rect 13955 15997 13964 16031
rect 13912 15988 13964 15997
rect 17868 16235 17920 16244
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 17776 16124 17828 16176
rect 18420 16167 18472 16176
rect 18420 16133 18429 16167
rect 18429 16133 18463 16167
rect 18463 16133 18472 16167
rect 18420 16124 18472 16133
rect 17224 15988 17276 16040
rect 17776 15988 17828 16040
rect 17868 15988 17920 16040
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 2228 15852 2280 15904
rect 2320 15895 2372 15904
rect 2320 15861 2329 15895
rect 2329 15861 2363 15895
rect 2363 15861 2372 15895
rect 2320 15852 2372 15861
rect 2412 15852 2464 15904
rect 5448 15852 5500 15904
rect 6276 15852 6328 15904
rect 7840 15895 7892 15904
rect 7840 15861 7849 15895
rect 7849 15861 7883 15895
rect 7883 15861 7892 15895
rect 7840 15852 7892 15861
rect 15200 15920 15252 15972
rect 11152 15852 11204 15904
rect 11428 15852 11480 15904
rect 12072 15852 12124 15904
rect 12164 15852 12216 15904
rect 13176 15852 13228 15904
rect 13544 15852 13596 15904
rect 14096 15852 14148 15904
rect 17316 15852 17368 15904
rect 17960 15852 18012 15904
rect 18604 15852 18656 15904
rect 5112 15750 5164 15802
rect 5176 15750 5228 15802
rect 5240 15750 5292 15802
rect 5304 15750 5356 15802
rect 5368 15750 5420 15802
rect 9827 15750 9879 15802
rect 9891 15750 9943 15802
rect 9955 15750 10007 15802
rect 10019 15750 10071 15802
rect 10083 15750 10135 15802
rect 14542 15750 14594 15802
rect 14606 15750 14658 15802
rect 14670 15750 14722 15802
rect 14734 15750 14786 15802
rect 14798 15750 14850 15802
rect 19257 15750 19309 15802
rect 19321 15750 19373 15802
rect 19385 15750 19437 15802
rect 19449 15750 19501 15802
rect 19513 15750 19565 15802
rect 1768 15648 1820 15700
rect 5540 15691 5592 15700
rect 5540 15657 5549 15691
rect 5549 15657 5583 15691
rect 5583 15657 5592 15691
rect 5540 15648 5592 15657
rect 1492 15555 1544 15564
rect 1492 15521 1501 15555
rect 1501 15521 1535 15555
rect 1535 15521 1544 15555
rect 2228 15580 2280 15632
rect 2504 15580 2556 15632
rect 1492 15512 1544 15521
rect 2412 15555 2464 15564
rect 2412 15521 2421 15555
rect 2421 15521 2455 15555
rect 2455 15521 2464 15555
rect 2412 15512 2464 15521
rect 3332 15512 3384 15564
rect 3608 15512 3660 15564
rect 4160 15512 4212 15564
rect 2320 15444 2372 15496
rect 2044 15376 2096 15428
rect 7564 15691 7616 15700
rect 7564 15657 7573 15691
rect 7573 15657 7607 15691
rect 7607 15657 7616 15691
rect 7564 15648 7616 15657
rect 7840 15648 7892 15700
rect 11060 15691 11112 15700
rect 11060 15657 11069 15691
rect 11069 15657 11103 15691
rect 11103 15657 11112 15691
rect 11060 15648 11112 15657
rect 6460 15555 6512 15564
rect 6460 15521 6469 15555
rect 6469 15521 6503 15555
rect 6503 15521 6512 15555
rect 6460 15512 6512 15521
rect 6552 15444 6604 15496
rect 7288 15512 7340 15564
rect 7380 15555 7432 15564
rect 7380 15521 7389 15555
rect 7389 15521 7423 15555
rect 7423 15521 7432 15555
rect 7380 15512 7432 15521
rect 11520 15623 11572 15632
rect 11520 15589 11529 15623
rect 11529 15589 11563 15623
rect 11563 15589 11572 15623
rect 11520 15580 11572 15589
rect 11980 15648 12032 15700
rect 12072 15691 12124 15700
rect 12072 15657 12081 15691
rect 12081 15657 12115 15691
rect 12115 15657 12124 15691
rect 12072 15648 12124 15657
rect 12348 15691 12400 15700
rect 12348 15657 12357 15691
rect 12357 15657 12391 15691
rect 12391 15657 12400 15691
rect 12348 15648 12400 15657
rect 13176 15648 13228 15700
rect 11612 15555 11664 15564
rect 11612 15521 11621 15555
rect 11621 15521 11655 15555
rect 11655 15521 11664 15555
rect 11612 15512 11664 15521
rect 11888 15512 11940 15564
rect 12072 15512 12124 15564
rect 12716 15555 12768 15564
rect 12716 15521 12725 15555
rect 12725 15521 12759 15555
rect 12759 15521 12768 15555
rect 12716 15512 12768 15521
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 12808 15444 12860 15496
rect 14004 15648 14056 15700
rect 17316 15691 17368 15700
rect 17316 15657 17325 15691
rect 17325 15657 17359 15691
rect 17359 15657 17368 15691
rect 17316 15648 17368 15657
rect 17500 15648 17552 15700
rect 18420 15648 18472 15700
rect 13544 15555 13596 15564
rect 13544 15521 13553 15555
rect 13553 15521 13587 15555
rect 13587 15521 13596 15555
rect 13544 15512 13596 15521
rect 14096 15555 14148 15564
rect 14096 15521 14105 15555
rect 14105 15521 14139 15555
rect 14139 15521 14148 15555
rect 14096 15512 14148 15521
rect 14924 15580 14976 15632
rect 14464 15512 14516 15564
rect 15108 15512 15160 15564
rect 18236 15580 18288 15632
rect 1676 15351 1728 15360
rect 1676 15317 1685 15351
rect 1685 15317 1719 15351
rect 1719 15317 1728 15351
rect 1676 15308 1728 15317
rect 2228 15351 2280 15360
rect 2228 15317 2237 15351
rect 2237 15317 2271 15351
rect 2271 15317 2280 15351
rect 2228 15308 2280 15317
rect 5356 15308 5408 15360
rect 6276 15376 6328 15428
rect 10692 15376 10744 15428
rect 8300 15308 8352 15360
rect 11796 15351 11848 15360
rect 11796 15317 11805 15351
rect 11805 15317 11839 15351
rect 11839 15317 11848 15351
rect 11796 15308 11848 15317
rect 12532 15308 12584 15360
rect 13544 15308 13596 15360
rect 18696 15555 18748 15564
rect 18696 15521 18705 15555
rect 18705 15521 18739 15555
rect 18739 15521 18748 15555
rect 18696 15512 18748 15521
rect 18880 15555 18932 15564
rect 18880 15521 18889 15555
rect 18889 15521 18923 15555
rect 18923 15521 18932 15555
rect 18880 15512 18932 15521
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 16580 15308 16632 15360
rect 17408 15308 17460 15360
rect 17868 15351 17920 15360
rect 17868 15317 17877 15351
rect 17877 15317 17911 15351
rect 17911 15317 17920 15351
rect 17868 15308 17920 15317
rect 18328 15351 18380 15360
rect 18328 15317 18337 15351
rect 18337 15317 18371 15351
rect 18371 15317 18380 15351
rect 18328 15308 18380 15317
rect 2755 15206 2807 15258
rect 2819 15206 2871 15258
rect 2883 15206 2935 15258
rect 2947 15206 2999 15258
rect 3011 15206 3063 15258
rect 7470 15206 7522 15258
rect 7534 15206 7586 15258
rect 7598 15206 7650 15258
rect 7662 15206 7714 15258
rect 7726 15206 7778 15258
rect 12185 15206 12237 15258
rect 12249 15206 12301 15258
rect 12313 15206 12365 15258
rect 12377 15206 12429 15258
rect 12441 15206 12493 15258
rect 16900 15206 16952 15258
rect 16964 15206 17016 15258
rect 17028 15206 17080 15258
rect 17092 15206 17144 15258
rect 17156 15206 17208 15258
rect 6552 15104 6604 15156
rect 7380 15104 7432 15156
rect 9404 15104 9456 15156
rect 2412 15036 2464 15088
rect 1492 14943 1544 14952
rect 1492 14909 1526 14943
rect 1526 14909 1544 14943
rect 1492 14900 1544 14909
rect 2320 14900 2372 14952
rect 2872 14832 2924 14884
rect 3332 14900 3384 14952
rect 3516 14875 3568 14884
rect 3516 14841 3550 14875
rect 3550 14841 3568 14875
rect 3516 14832 3568 14841
rect 5356 14875 5408 14884
rect 5356 14841 5390 14875
rect 5390 14841 5408 14875
rect 5356 14832 5408 14841
rect 5908 14832 5960 14884
rect 7564 14943 7616 14952
rect 7564 14909 7573 14943
rect 7573 14909 7607 14943
rect 7607 14909 7616 14943
rect 7564 14900 7616 14909
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 8208 14900 8260 14952
rect 8576 14900 8628 14952
rect 2596 14764 2648 14816
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 6276 14764 6328 14816
rect 6368 14764 6420 14816
rect 9036 14900 9088 14952
rect 9588 15036 9640 15088
rect 9404 14900 9456 14952
rect 9588 14900 9640 14952
rect 10416 15104 10468 15156
rect 11612 15104 11664 15156
rect 12256 15104 12308 15156
rect 12624 15104 12676 15156
rect 12716 15104 12768 15156
rect 12808 15104 12860 15156
rect 14280 15104 14332 15156
rect 12072 15036 12124 15088
rect 10692 14900 10744 14952
rect 11060 14943 11112 14952
rect 11060 14909 11078 14943
rect 11078 14909 11112 14943
rect 11060 14900 11112 14909
rect 12808 14968 12860 15020
rect 12532 14900 12584 14952
rect 14280 14900 14332 14952
rect 13912 14832 13964 14884
rect 7380 14764 7432 14816
rect 8944 14764 8996 14816
rect 9588 14764 9640 14816
rect 10600 14764 10652 14816
rect 11612 14807 11664 14816
rect 11612 14773 11621 14807
rect 11621 14773 11655 14807
rect 11655 14773 11664 14807
rect 11612 14764 11664 14773
rect 12072 14807 12124 14816
rect 12072 14773 12081 14807
rect 12081 14773 12115 14807
rect 12115 14773 12124 14807
rect 12072 14764 12124 14773
rect 12532 14764 12584 14816
rect 13268 14764 13320 14816
rect 14004 14764 14056 14816
rect 15108 14900 15160 14952
rect 17592 14943 17644 14952
rect 17592 14909 17610 14943
rect 17610 14909 17644 14943
rect 17592 14900 17644 14909
rect 17776 14900 17828 14952
rect 18696 15104 18748 15156
rect 18880 15104 18932 15156
rect 18972 14900 19024 14952
rect 14464 14832 14516 14884
rect 18604 14832 18656 14884
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 16396 14764 16448 14773
rect 16488 14807 16540 14816
rect 16488 14773 16497 14807
rect 16497 14773 16531 14807
rect 16531 14773 16540 14807
rect 16488 14764 16540 14773
rect 18236 14764 18288 14816
rect 18696 14764 18748 14816
rect 5112 14662 5164 14714
rect 5176 14662 5228 14714
rect 5240 14662 5292 14714
rect 5304 14662 5356 14714
rect 5368 14662 5420 14714
rect 9827 14662 9879 14714
rect 9891 14662 9943 14714
rect 9955 14662 10007 14714
rect 10019 14662 10071 14714
rect 10083 14662 10135 14714
rect 14542 14662 14594 14714
rect 14606 14662 14658 14714
rect 14670 14662 14722 14714
rect 14734 14662 14786 14714
rect 14798 14662 14850 14714
rect 19257 14662 19309 14714
rect 19321 14662 19373 14714
rect 19385 14662 19437 14714
rect 19449 14662 19501 14714
rect 19513 14662 19565 14714
rect 1584 14560 1636 14612
rect 2596 14560 2648 14612
rect 5908 14603 5960 14612
rect 5908 14569 5917 14603
rect 5917 14569 5951 14603
rect 5951 14569 5960 14603
rect 5908 14560 5960 14569
rect 2044 14492 2096 14544
rect 1676 14424 1728 14476
rect 2872 14492 2924 14544
rect 2228 14424 2280 14476
rect 5908 14424 5960 14476
rect 6460 14560 6512 14612
rect 7564 14560 7616 14612
rect 6276 14288 6328 14340
rect 9588 14560 9640 14612
rect 12072 14560 12124 14612
rect 7932 14492 7984 14544
rect 11060 14492 11112 14544
rect 15200 14560 15252 14612
rect 8852 14424 8904 14476
rect 9036 14467 9088 14476
rect 9036 14433 9070 14467
rect 9070 14433 9088 14467
rect 9036 14424 9088 14433
rect 10692 14424 10744 14476
rect 8392 14356 8444 14408
rect 11612 14424 11664 14476
rect 12256 14424 12308 14476
rect 18420 14492 18472 14544
rect 18972 14535 19024 14544
rect 18972 14501 18981 14535
rect 18981 14501 19015 14535
rect 19015 14501 19024 14535
rect 18972 14492 19024 14501
rect 13912 14467 13964 14476
rect 13912 14433 13946 14467
rect 13946 14433 13964 14467
rect 13912 14424 13964 14433
rect 14280 14424 14332 14476
rect 14464 14424 14516 14476
rect 15660 14424 15712 14476
rect 16212 14424 16264 14476
rect 12532 14399 12584 14408
rect 7840 14288 7892 14340
rect 8668 14288 8720 14340
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 15476 14356 15528 14408
rect 16120 14356 16172 14408
rect 1400 14263 1452 14272
rect 1400 14229 1409 14263
rect 1409 14229 1443 14263
rect 1443 14229 1452 14263
rect 1400 14220 1452 14229
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 4436 14220 4488 14272
rect 6644 14220 6696 14272
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 7288 14220 7340 14229
rect 8576 14220 8628 14272
rect 9128 14220 9180 14272
rect 15936 14288 15988 14340
rect 16580 14424 16632 14476
rect 18696 14424 18748 14476
rect 18880 14467 18932 14476
rect 18880 14433 18889 14467
rect 18889 14433 18923 14467
rect 18923 14433 18932 14467
rect 18880 14424 18932 14433
rect 10232 14220 10284 14272
rect 11336 14220 11388 14272
rect 15016 14263 15068 14272
rect 15016 14229 15025 14263
rect 15025 14229 15059 14263
rect 15059 14229 15068 14263
rect 15016 14220 15068 14229
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 18512 14220 18564 14272
rect 2755 14118 2807 14170
rect 2819 14118 2871 14170
rect 2883 14118 2935 14170
rect 2947 14118 2999 14170
rect 3011 14118 3063 14170
rect 7470 14118 7522 14170
rect 7534 14118 7586 14170
rect 7598 14118 7650 14170
rect 7662 14118 7714 14170
rect 7726 14118 7778 14170
rect 12185 14118 12237 14170
rect 12249 14118 12301 14170
rect 12313 14118 12365 14170
rect 12377 14118 12429 14170
rect 12441 14118 12493 14170
rect 16900 14118 16952 14170
rect 16964 14118 17016 14170
rect 17028 14118 17080 14170
rect 17092 14118 17144 14170
rect 17156 14118 17208 14170
rect 1400 14016 1452 14068
rect 1768 14016 1820 14068
rect 1952 14016 2004 14068
rect 2596 14016 2648 14068
rect 6552 14016 6604 14068
rect 7840 14016 7892 14068
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 12992 14016 13044 14068
rect 1584 13812 1636 13864
rect 2136 13880 2188 13932
rect 7748 13948 7800 14000
rect 8208 13948 8260 14000
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 3332 13880 3384 13932
rect 7288 13880 7340 13932
rect 5632 13855 5684 13864
rect 5632 13821 5641 13855
rect 5641 13821 5675 13855
rect 5675 13821 5684 13855
rect 5632 13812 5684 13821
rect 5908 13855 5960 13864
rect 5908 13821 5942 13855
rect 5942 13821 5960 13855
rect 5908 13812 5960 13821
rect 7380 13812 7432 13864
rect 8024 13812 8076 13864
rect 8576 13855 8628 13864
rect 8576 13821 8585 13855
rect 8585 13821 8619 13855
rect 8619 13821 8628 13855
rect 8576 13812 8628 13821
rect 8944 13880 8996 13932
rect 13268 14016 13320 14068
rect 15016 14016 15068 14068
rect 17408 14016 17460 14068
rect 18880 14016 18932 14068
rect 9128 13855 9180 13864
rect 9128 13821 9137 13855
rect 9137 13821 9171 13855
rect 9171 13821 9180 13855
rect 9128 13812 9180 13821
rect 14280 13880 14332 13932
rect 14464 13923 14516 13932
rect 14464 13889 14473 13923
rect 14473 13889 14507 13923
rect 14507 13889 14516 13923
rect 14464 13880 14516 13889
rect 3240 13744 3292 13796
rect 6276 13744 6328 13796
rect 15016 13812 15068 13864
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 16488 13812 16540 13864
rect 16212 13744 16264 13796
rect 2504 13676 2556 13728
rect 2596 13676 2648 13728
rect 3148 13676 3200 13728
rect 4528 13676 4580 13728
rect 7012 13719 7064 13728
rect 7012 13685 7021 13719
rect 7021 13685 7055 13719
rect 7055 13685 7064 13719
rect 7012 13676 7064 13685
rect 7656 13676 7708 13728
rect 9036 13676 9088 13728
rect 13728 13676 13780 13728
rect 13820 13676 13872 13728
rect 15292 13719 15344 13728
rect 15292 13685 15301 13719
rect 15301 13685 15335 13719
rect 15335 13685 15344 13719
rect 15292 13676 15344 13685
rect 16028 13676 16080 13728
rect 16580 13676 16632 13728
rect 17776 13812 17828 13864
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 18604 13812 18656 13864
rect 18788 13744 18840 13796
rect 18144 13676 18196 13728
rect 18972 13676 19024 13728
rect 5112 13574 5164 13626
rect 5176 13574 5228 13626
rect 5240 13574 5292 13626
rect 5304 13574 5356 13626
rect 5368 13574 5420 13626
rect 9827 13574 9879 13626
rect 9891 13574 9943 13626
rect 9955 13574 10007 13626
rect 10019 13574 10071 13626
rect 10083 13574 10135 13626
rect 14542 13574 14594 13626
rect 14606 13574 14658 13626
rect 14670 13574 14722 13626
rect 14734 13574 14786 13626
rect 14798 13574 14850 13626
rect 19257 13574 19309 13626
rect 19321 13574 19373 13626
rect 19385 13574 19437 13626
rect 19449 13574 19501 13626
rect 19513 13574 19565 13626
rect 6092 13472 6144 13524
rect 7380 13472 7432 13524
rect 1584 13404 1636 13456
rect 3240 13404 3292 13456
rect 3332 13447 3384 13456
rect 3332 13413 3341 13447
rect 3341 13413 3375 13447
rect 3375 13413 3384 13447
rect 3332 13404 3384 13413
rect 4160 13447 4212 13456
rect 4160 13413 4169 13447
rect 4169 13413 4203 13447
rect 4203 13413 4212 13447
rect 4160 13404 4212 13413
rect 7932 13404 7984 13456
rect 8576 13404 8628 13456
rect 12716 13404 12768 13456
rect 1216 13336 1268 13388
rect 2504 13336 2556 13388
rect 4528 13379 4580 13388
rect 3240 13268 3292 13320
rect 4528 13345 4562 13379
rect 4562 13345 4580 13379
rect 4528 13336 4580 13345
rect 4896 13336 4948 13388
rect 4252 13311 4304 13320
rect 4252 13277 4261 13311
rect 4261 13277 4295 13311
rect 4295 13277 4304 13311
rect 4252 13268 4304 13277
rect 6092 13379 6144 13388
rect 6092 13345 6101 13379
rect 6101 13345 6135 13379
rect 6135 13345 6144 13379
rect 6092 13336 6144 13345
rect 6276 13336 6328 13388
rect 6368 13379 6420 13388
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 6552 13336 6604 13388
rect 7012 13336 7064 13388
rect 7656 13379 7708 13388
rect 7656 13345 7665 13379
rect 7665 13345 7699 13379
rect 7699 13345 7708 13379
rect 7656 13336 7708 13345
rect 3516 13200 3568 13252
rect 2596 13132 2648 13184
rect 6368 13132 6420 13184
rect 6736 13268 6788 13320
rect 8668 13379 8720 13388
rect 8668 13345 8677 13379
rect 8677 13345 8711 13379
rect 8711 13345 8720 13379
rect 8668 13336 8720 13345
rect 10600 13336 10652 13388
rect 12532 13268 12584 13320
rect 8576 13132 8628 13184
rect 10048 13175 10100 13184
rect 10048 13141 10057 13175
rect 10057 13141 10091 13175
rect 10091 13141 10100 13175
rect 10048 13132 10100 13141
rect 10968 13175 11020 13184
rect 10968 13141 10977 13175
rect 10977 13141 11011 13175
rect 11011 13141 11020 13175
rect 10968 13132 11020 13141
rect 13084 13336 13136 13388
rect 13820 13472 13872 13524
rect 14280 13515 14332 13524
rect 14280 13481 14289 13515
rect 14289 13481 14323 13515
rect 14323 13481 14332 13515
rect 14280 13472 14332 13481
rect 16120 13472 16172 13524
rect 16212 13472 16264 13524
rect 13544 13379 13596 13388
rect 13544 13345 13553 13379
rect 13553 13345 13587 13379
rect 13587 13345 13596 13379
rect 13544 13336 13596 13345
rect 13820 13379 13872 13388
rect 13820 13345 13829 13379
rect 13829 13345 13863 13379
rect 13863 13345 13872 13379
rect 13820 13336 13872 13345
rect 15200 13404 15252 13456
rect 17224 13404 17276 13456
rect 12992 13200 13044 13252
rect 16028 13336 16080 13388
rect 18604 13379 18656 13388
rect 18604 13345 18613 13379
rect 18613 13345 18647 13379
rect 18647 13345 18656 13379
rect 18604 13336 18656 13345
rect 17776 13268 17828 13320
rect 13360 13132 13412 13184
rect 13820 13132 13872 13184
rect 14188 13132 14240 13184
rect 14556 13175 14608 13184
rect 14556 13141 14565 13175
rect 14565 13141 14599 13175
rect 14599 13141 14608 13175
rect 14556 13132 14608 13141
rect 16488 13132 16540 13184
rect 2755 13030 2807 13082
rect 2819 13030 2871 13082
rect 2883 13030 2935 13082
rect 2947 13030 2999 13082
rect 3011 13030 3063 13082
rect 7470 13030 7522 13082
rect 7534 13030 7586 13082
rect 7598 13030 7650 13082
rect 7662 13030 7714 13082
rect 7726 13030 7778 13082
rect 12185 13030 12237 13082
rect 12249 13030 12301 13082
rect 12313 13030 12365 13082
rect 12377 13030 12429 13082
rect 12441 13030 12493 13082
rect 16900 13030 16952 13082
rect 16964 13030 17016 13082
rect 17028 13030 17080 13082
rect 17092 13030 17144 13082
rect 17156 13030 17208 13082
rect 3976 12928 4028 12980
rect 2596 12860 2648 12912
rect 3240 12792 3292 12844
rect 3148 12656 3200 12708
rect 4252 12792 4304 12844
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 5632 12928 5684 12980
rect 6828 12928 6880 12980
rect 8116 12928 8168 12980
rect 4712 12792 4764 12801
rect 4160 12724 4212 12776
rect 4528 12724 4580 12776
rect 7380 12792 7432 12844
rect 7104 12767 7156 12776
rect 7104 12733 7113 12767
rect 7113 12733 7147 12767
rect 7147 12733 7156 12767
rect 7104 12724 7156 12733
rect 10048 12860 10100 12912
rect 10140 12860 10192 12912
rect 2504 12588 2556 12640
rect 3884 12588 3936 12640
rect 4252 12588 4304 12640
rect 5448 12656 5500 12708
rect 8024 12767 8076 12776
rect 8024 12733 8033 12767
rect 8033 12733 8067 12767
rect 8067 12733 8076 12767
rect 8024 12724 8076 12733
rect 8760 12767 8812 12776
rect 8760 12733 8769 12767
rect 8769 12733 8803 12767
rect 8803 12733 8812 12767
rect 9312 12792 9364 12844
rect 8760 12724 8812 12733
rect 9220 12724 9272 12776
rect 10416 12792 10468 12844
rect 12900 12860 12952 12912
rect 13360 12860 13412 12912
rect 11152 12792 11204 12844
rect 13820 12928 13872 12980
rect 13912 12971 13964 12980
rect 13912 12937 13921 12971
rect 13921 12937 13955 12971
rect 13955 12937 13964 12971
rect 13912 12928 13964 12937
rect 17592 12928 17644 12980
rect 18328 12971 18380 12980
rect 18328 12937 18337 12971
rect 18337 12937 18371 12971
rect 18371 12937 18380 12971
rect 18328 12928 18380 12937
rect 18696 12928 18748 12980
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 8668 12699 8720 12708
rect 8668 12665 8677 12699
rect 8677 12665 8711 12699
rect 8711 12665 8720 12699
rect 8668 12656 8720 12665
rect 9496 12588 9548 12640
rect 10876 12767 10928 12776
rect 10876 12733 10885 12767
rect 10885 12733 10919 12767
rect 10919 12733 10928 12767
rect 10876 12724 10928 12733
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 10692 12656 10744 12708
rect 11612 12588 11664 12640
rect 11796 12588 11848 12640
rect 12072 12588 12124 12640
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 13544 12724 13596 12776
rect 14556 12860 14608 12912
rect 14372 12792 14424 12844
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 13820 12767 13872 12776
rect 13820 12733 13829 12767
rect 13829 12733 13863 12767
rect 13863 12733 13872 12767
rect 13820 12724 13872 12733
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 14464 12724 14516 12776
rect 14832 12724 14884 12776
rect 16212 12656 16264 12708
rect 17224 12767 17276 12776
rect 17224 12733 17233 12767
rect 17233 12733 17267 12767
rect 17267 12733 17276 12767
rect 17224 12724 17276 12733
rect 18420 12767 18472 12776
rect 18420 12733 18429 12767
rect 18429 12733 18463 12767
rect 18463 12733 18472 12767
rect 18420 12724 18472 12733
rect 18880 12767 18932 12776
rect 18880 12733 18889 12767
rect 18889 12733 18923 12767
rect 18923 12733 18932 12767
rect 18880 12724 18932 12733
rect 13912 12588 13964 12640
rect 15752 12631 15804 12640
rect 15752 12597 15761 12631
rect 15761 12597 15795 12631
rect 15795 12597 15804 12631
rect 15752 12588 15804 12597
rect 18880 12588 18932 12640
rect 5112 12486 5164 12538
rect 5176 12486 5228 12538
rect 5240 12486 5292 12538
rect 5304 12486 5356 12538
rect 5368 12486 5420 12538
rect 9827 12486 9879 12538
rect 9891 12486 9943 12538
rect 9955 12486 10007 12538
rect 10019 12486 10071 12538
rect 10083 12486 10135 12538
rect 14542 12486 14594 12538
rect 14606 12486 14658 12538
rect 14670 12486 14722 12538
rect 14734 12486 14786 12538
rect 14798 12486 14850 12538
rect 19257 12486 19309 12538
rect 19321 12486 19373 12538
rect 19385 12486 19437 12538
rect 19449 12486 19501 12538
rect 19513 12486 19565 12538
rect 1308 12316 1360 12368
rect 2412 12316 2464 12368
rect 2596 12291 2648 12300
rect 2596 12257 2605 12291
rect 2605 12257 2639 12291
rect 2639 12257 2648 12291
rect 2596 12248 2648 12257
rect 1216 12044 1268 12096
rect 2412 12044 2464 12096
rect 3608 12384 3660 12436
rect 5448 12384 5500 12436
rect 3516 12359 3568 12368
rect 3516 12325 3525 12359
rect 3525 12325 3559 12359
rect 3559 12325 3568 12359
rect 3516 12316 3568 12325
rect 3516 12180 3568 12232
rect 3884 12248 3936 12300
rect 3976 12248 4028 12300
rect 4712 12316 4764 12368
rect 4896 12180 4948 12232
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 5632 12248 5684 12300
rect 6736 12316 6788 12368
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 4252 12112 4304 12164
rect 4436 12112 4488 12164
rect 3608 12044 3660 12096
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 4712 12087 4764 12096
rect 4712 12053 4721 12087
rect 4721 12053 4755 12087
rect 4755 12053 4764 12087
rect 4712 12044 4764 12053
rect 4804 12044 4856 12096
rect 7196 12180 7248 12232
rect 9220 12427 9272 12436
rect 9220 12393 9229 12427
rect 9229 12393 9263 12427
rect 9263 12393 9272 12427
rect 9220 12384 9272 12393
rect 10876 12384 10928 12436
rect 10324 12316 10376 12368
rect 10508 12359 10560 12368
rect 10508 12325 10517 12359
rect 10517 12325 10551 12359
rect 10551 12325 10560 12359
rect 10508 12316 10560 12325
rect 9496 12248 9548 12300
rect 9584 12180 9636 12232
rect 9772 12248 9824 12300
rect 12532 12316 12584 12368
rect 10048 12180 10100 12232
rect 10324 12180 10376 12232
rect 10784 12180 10836 12232
rect 12808 12248 12860 12300
rect 14280 12359 14332 12368
rect 14280 12325 14289 12359
rect 14289 12325 14323 12359
rect 14323 12325 14332 12359
rect 14280 12316 14332 12325
rect 14096 12291 14148 12300
rect 14096 12257 14105 12291
rect 14105 12257 14139 12291
rect 14139 12257 14148 12291
rect 14096 12248 14148 12257
rect 16028 12316 16080 12368
rect 15752 12248 15804 12300
rect 17592 12427 17644 12436
rect 17592 12393 17601 12427
rect 17601 12393 17635 12427
rect 17635 12393 17644 12427
rect 17592 12384 17644 12393
rect 5724 12044 5776 12096
rect 8208 12044 8260 12096
rect 10140 12044 10192 12096
rect 11152 12044 11204 12096
rect 12532 12044 12584 12096
rect 13636 12044 13688 12096
rect 16212 12180 16264 12232
rect 14372 12112 14424 12164
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 17316 12248 17368 12257
rect 18696 12291 18748 12300
rect 18696 12257 18714 12291
rect 18714 12257 18748 12291
rect 18696 12248 18748 12257
rect 18880 12248 18932 12300
rect 16580 12223 16632 12232
rect 16580 12189 16589 12223
rect 16589 12189 16623 12223
rect 16623 12189 16632 12223
rect 16580 12180 16632 12189
rect 15108 12044 15160 12096
rect 15660 12044 15712 12096
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 15844 12044 15896 12096
rect 2755 11942 2807 11994
rect 2819 11942 2871 11994
rect 2883 11942 2935 11994
rect 2947 11942 2999 11994
rect 3011 11942 3063 11994
rect 7470 11942 7522 11994
rect 7534 11942 7586 11994
rect 7598 11942 7650 11994
rect 7662 11942 7714 11994
rect 7726 11942 7778 11994
rect 12185 11942 12237 11994
rect 12249 11942 12301 11994
rect 12313 11942 12365 11994
rect 12377 11942 12429 11994
rect 12441 11942 12493 11994
rect 16900 11942 16952 11994
rect 16964 11942 17016 11994
rect 17028 11942 17080 11994
rect 17092 11942 17144 11994
rect 17156 11942 17208 11994
rect 2596 11840 2648 11892
rect 3884 11883 3936 11892
rect 3884 11849 3893 11883
rect 3893 11849 3927 11883
rect 3927 11849 3936 11883
rect 3884 11840 3936 11849
rect 11244 11840 11296 11892
rect 11704 11883 11756 11892
rect 11704 11849 11713 11883
rect 11713 11849 11747 11883
rect 11747 11849 11756 11883
rect 11704 11840 11756 11849
rect 12532 11840 12584 11892
rect 12900 11840 12952 11892
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 14280 11840 14332 11892
rect 16028 11840 16080 11892
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 18420 11840 18472 11849
rect 18788 11883 18840 11892
rect 18788 11849 18797 11883
rect 18797 11849 18831 11883
rect 18831 11849 18840 11883
rect 18788 11840 18840 11849
rect 2504 11772 2556 11824
rect 4712 11772 4764 11824
rect 1768 11636 1820 11688
rect 4436 11704 4488 11756
rect 3976 11679 4028 11688
rect 1400 11568 1452 11620
rect 3976 11645 3985 11679
rect 3985 11645 4019 11679
rect 4019 11645 4028 11679
rect 3976 11636 4028 11645
rect 4804 11636 4856 11688
rect 5724 11704 5776 11756
rect 5080 11636 5132 11688
rect 4712 11611 4764 11620
rect 4712 11577 4721 11611
rect 4721 11577 4755 11611
rect 4755 11577 4764 11611
rect 4712 11568 4764 11577
rect 4988 11611 5040 11620
rect 4988 11577 4997 11611
rect 4997 11577 5031 11611
rect 5031 11577 5040 11611
rect 4988 11568 5040 11577
rect 7564 11636 7616 11688
rect 10048 11704 10100 11756
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 9220 11636 9272 11688
rect 9588 11679 9640 11688
rect 9588 11645 9617 11679
rect 9617 11645 9640 11679
rect 9588 11636 9640 11645
rect 9864 11679 9916 11688
rect 9864 11645 9873 11679
rect 9873 11645 9907 11679
rect 9907 11645 9916 11679
rect 9864 11636 9916 11645
rect 10416 11636 10468 11688
rect 10508 11636 10560 11688
rect 9496 11568 9548 11620
rect 10876 11611 10928 11620
rect 10876 11577 10885 11611
rect 10885 11577 10919 11611
rect 10919 11577 10928 11611
rect 10876 11568 10928 11577
rect 1216 11500 1268 11552
rect 3332 11500 3384 11552
rect 5816 11543 5868 11552
rect 5816 11509 5825 11543
rect 5825 11509 5859 11543
rect 5859 11509 5868 11543
rect 5816 11500 5868 11509
rect 6092 11543 6144 11552
rect 6092 11509 6101 11543
rect 6101 11509 6135 11543
rect 6135 11509 6144 11543
rect 6092 11500 6144 11509
rect 8024 11500 8076 11552
rect 9312 11500 9364 11552
rect 9404 11500 9456 11552
rect 13636 11747 13688 11756
rect 11612 11636 11664 11688
rect 12532 11636 12584 11688
rect 13636 11713 13645 11747
rect 13645 11713 13679 11747
rect 13679 11713 13688 11747
rect 13636 11704 13688 11713
rect 14096 11704 14148 11756
rect 12808 11568 12860 11620
rect 13820 11568 13872 11620
rect 14464 11636 14516 11688
rect 15660 11704 15712 11756
rect 15752 11704 15804 11756
rect 15476 11679 15528 11688
rect 15476 11645 15485 11679
rect 15485 11645 15519 11679
rect 15519 11645 15528 11679
rect 15476 11636 15528 11645
rect 16304 11679 16356 11688
rect 16304 11645 16313 11679
rect 16313 11645 16347 11679
rect 16347 11645 16356 11679
rect 16304 11636 16356 11645
rect 16488 11636 16540 11688
rect 13728 11500 13780 11552
rect 14372 11500 14424 11552
rect 14924 11500 14976 11552
rect 18420 11636 18472 11688
rect 18604 11636 18656 11688
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 17684 11543 17736 11552
rect 17684 11509 17693 11543
rect 17693 11509 17727 11543
rect 17727 11509 17736 11543
rect 17684 11500 17736 11509
rect 18144 11543 18196 11552
rect 18144 11509 18153 11543
rect 18153 11509 18187 11543
rect 18187 11509 18196 11543
rect 18144 11500 18196 11509
rect 18512 11500 18564 11552
rect 5112 11398 5164 11450
rect 5176 11398 5228 11450
rect 5240 11398 5292 11450
rect 5304 11398 5356 11450
rect 5368 11398 5420 11450
rect 9827 11398 9879 11450
rect 9891 11398 9943 11450
rect 9955 11398 10007 11450
rect 10019 11398 10071 11450
rect 10083 11398 10135 11450
rect 14542 11398 14594 11450
rect 14606 11398 14658 11450
rect 14670 11398 14722 11450
rect 14734 11398 14786 11450
rect 14798 11398 14850 11450
rect 19257 11398 19309 11450
rect 19321 11398 19373 11450
rect 19385 11398 19437 11450
rect 19449 11398 19501 11450
rect 19513 11398 19565 11450
rect 1308 11339 1360 11348
rect 1308 11305 1317 11339
rect 1317 11305 1351 11339
rect 1351 11305 1360 11339
rect 1308 11296 1360 11305
rect 1400 11228 1452 11280
rect 1216 11092 1268 11144
rect 3240 11228 3292 11280
rect 1768 11203 1820 11212
rect 1768 11169 1802 11203
rect 1802 11169 1820 11203
rect 1768 11160 1820 11169
rect 4344 11228 4396 11280
rect 7564 11339 7616 11348
rect 7564 11305 7573 11339
rect 7573 11305 7607 11339
rect 7607 11305 7616 11339
rect 7564 11296 7616 11305
rect 3976 11160 4028 11212
rect 4712 11160 4764 11212
rect 4988 11160 5040 11212
rect 5816 11160 5868 11212
rect 8116 11228 8168 11280
rect 9588 11296 9640 11348
rect 10508 11339 10560 11348
rect 10508 11305 10517 11339
rect 10517 11305 10551 11339
rect 10551 11305 10560 11339
rect 10508 11296 10560 11305
rect 14096 11296 14148 11348
rect 15200 11296 15252 11348
rect 7748 11160 7800 11212
rect 9496 11203 9548 11212
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 9496 11160 9548 11169
rect 9772 11203 9824 11212
rect 9772 11169 9781 11203
rect 9781 11169 9815 11203
rect 9815 11169 9824 11203
rect 9772 11160 9824 11169
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 3148 10956 3200 11008
rect 5448 10956 5500 11008
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 6000 10956 6052 10965
rect 6368 10956 6420 11008
rect 9404 10956 9456 11008
rect 9864 11024 9916 11076
rect 11612 11160 11664 11212
rect 14464 11228 14516 11280
rect 11796 11203 11848 11212
rect 11796 11169 11805 11203
rect 11805 11169 11839 11203
rect 11839 11169 11848 11203
rect 11796 11160 11848 11169
rect 13820 11203 13872 11212
rect 13820 11169 13838 11203
rect 13838 11169 13872 11203
rect 13820 11160 13872 11169
rect 13084 11092 13136 11144
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 14556 11203 14608 11212
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 14556 11160 14608 11169
rect 15568 11228 15620 11280
rect 16304 11296 16356 11348
rect 15476 11160 15528 11212
rect 16212 11203 16264 11212
rect 16212 11169 16221 11203
rect 16221 11169 16255 11203
rect 16255 11169 16264 11203
rect 16212 11160 16264 11169
rect 17684 11160 17736 11212
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 19064 11203 19116 11212
rect 19064 11169 19073 11203
rect 19073 11169 19107 11203
rect 19107 11169 19116 11203
rect 19064 11160 19116 11169
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 12072 10956 12124 11008
rect 13360 10956 13412 11008
rect 14924 10956 14976 11008
rect 15292 10999 15344 11008
rect 15292 10965 15301 10999
rect 15301 10965 15335 10999
rect 15335 10965 15344 10999
rect 15292 10956 15344 10965
rect 15660 10956 15712 11008
rect 18144 10956 18196 11008
rect 18696 10956 18748 11008
rect 2755 10854 2807 10906
rect 2819 10854 2871 10906
rect 2883 10854 2935 10906
rect 2947 10854 2999 10906
rect 3011 10854 3063 10906
rect 7470 10854 7522 10906
rect 7534 10854 7586 10906
rect 7598 10854 7650 10906
rect 7662 10854 7714 10906
rect 7726 10854 7778 10906
rect 12185 10854 12237 10906
rect 12249 10854 12301 10906
rect 12313 10854 12365 10906
rect 12377 10854 12429 10906
rect 12441 10854 12493 10906
rect 16900 10854 16952 10906
rect 16964 10854 17016 10906
rect 17028 10854 17080 10906
rect 17092 10854 17144 10906
rect 17156 10854 17208 10906
rect 2412 10548 2464 10600
rect 2504 10591 2556 10600
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 3516 10752 3568 10804
rect 6460 10795 6512 10804
rect 6460 10761 6469 10795
rect 6469 10761 6503 10795
rect 6503 10761 6512 10795
rect 6460 10752 6512 10761
rect 7196 10752 7248 10804
rect 9680 10795 9732 10804
rect 9680 10761 9689 10795
rect 9689 10761 9723 10795
rect 9723 10761 9732 10795
rect 9680 10752 9732 10761
rect 10048 10752 10100 10804
rect 11244 10752 11296 10804
rect 11796 10752 11848 10804
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 4988 10616 5040 10668
rect 3056 10548 3108 10600
rect 3148 10548 3200 10600
rect 3332 10548 3384 10600
rect 8024 10616 8076 10668
rect 8116 10616 8168 10668
rect 5632 10548 5684 10600
rect 6368 10548 6420 10600
rect 5632 10412 5684 10464
rect 6000 10412 6052 10464
rect 9680 10548 9732 10600
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 10508 10684 10560 10736
rect 9772 10480 9824 10532
rect 7748 10412 7800 10464
rect 10324 10548 10376 10600
rect 10968 10616 11020 10668
rect 10784 10548 10836 10600
rect 11428 10591 11480 10600
rect 11428 10557 11437 10591
rect 11437 10557 11471 10591
rect 11471 10557 11480 10591
rect 11428 10548 11480 10557
rect 11796 10616 11848 10668
rect 13912 10795 13964 10804
rect 13912 10761 13921 10795
rect 13921 10761 13955 10795
rect 13955 10761 13964 10795
rect 13912 10752 13964 10761
rect 14280 10752 14332 10804
rect 14556 10795 14608 10804
rect 14556 10761 14565 10795
rect 14565 10761 14599 10795
rect 14599 10761 14608 10795
rect 14556 10752 14608 10761
rect 18236 10752 18288 10804
rect 12072 10616 12124 10668
rect 10968 10480 11020 10532
rect 11244 10412 11296 10464
rect 12164 10591 12216 10600
rect 12164 10557 12173 10591
rect 12173 10557 12207 10591
rect 12207 10557 12216 10591
rect 12164 10548 12216 10557
rect 15292 10684 15344 10736
rect 15108 10548 15160 10600
rect 11980 10523 12032 10532
rect 11980 10489 11989 10523
rect 11989 10489 12023 10523
rect 12023 10489 12032 10523
rect 11980 10480 12032 10489
rect 15568 10523 15620 10532
rect 12624 10412 12676 10464
rect 15568 10489 15602 10523
rect 15602 10489 15620 10523
rect 15568 10480 15620 10489
rect 17684 10480 17736 10532
rect 18696 10591 18748 10600
rect 18696 10557 18705 10591
rect 18705 10557 18739 10591
rect 18739 10557 18748 10591
rect 18696 10548 18748 10557
rect 18880 10548 18932 10600
rect 18788 10523 18840 10532
rect 18788 10489 18797 10523
rect 18797 10489 18831 10523
rect 18831 10489 18840 10523
rect 18788 10480 18840 10489
rect 16212 10412 16264 10464
rect 16396 10412 16448 10464
rect 16764 10455 16816 10464
rect 16764 10421 16773 10455
rect 16773 10421 16807 10455
rect 16807 10421 16816 10455
rect 16764 10412 16816 10421
rect 5112 10310 5164 10362
rect 5176 10310 5228 10362
rect 5240 10310 5292 10362
rect 5304 10310 5356 10362
rect 5368 10310 5420 10362
rect 9827 10310 9879 10362
rect 9891 10310 9943 10362
rect 9955 10310 10007 10362
rect 10019 10310 10071 10362
rect 10083 10310 10135 10362
rect 14542 10310 14594 10362
rect 14606 10310 14658 10362
rect 14670 10310 14722 10362
rect 14734 10310 14786 10362
rect 14798 10310 14850 10362
rect 19257 10310 19309 10362
rect 19321 10310 19373 10362
rect 19385 10310 19437 10362
rect 19449 10310 19501 10362
rect 19513 10310 19565 10362
rect 5632 10208 5684 10260
rect 1584 10140 1636 10192
rect 3424 10140 3476 10192
rect 10692 10208 10744 10260
rect 11060 10208 11112 10260
rect 12072 10208 12124 10260
rect 14096 10208 14148 10260
rect 1216 10115 1268 10124
rect 1216 10081 1225 10115
rect 1225 10081 1259 10115
rect 1259 10081 1268 10115
rect 1216 10072 1268 10081
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 6000 10115 6052 10124
rect 6000 10081 6009 10115
rect 6009 10081 6043 10115
rect 6043 10081 6052 10115
rect 6000 10072 6052 10081
rect 6736 10115 6788 10124
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 6828 10072 6880 10124
rect 7564 10072 7616 10124
rect 6184 10004 6236 10056
rect 7748 10004 7800 10056
rect 9588 10047 9640 10056
rect 9588 10013 9597 10047
rect 9597 10013 9631 10047
rect 9631 10013 9640 10047
rect 9588 10004 9640 10013
rect 14464 10115 14516 10124
rect 18236 10140 18288 10192
rect 14464 10081 14482 10115
rect 14482 10081 14516 10115
rect 14464 10072 14516 10081
rect 15108 10072 15160 10124
rect 15844 10072 15896 10124
rect 16672 10115 16724 10124
rect 16672 10081 16681 10115
rect 16681 10081 16715 10115
rect 16715 10081 16724 10115
rect 16672 10072 16724 10081
rect 18880 10115 18932 10124
rect 18880 10081 18889 10115
rect 18889 10081 18923 10115
rect 18923 10081 18932 10115
rect 18880 10072 18932 10081
rect 10600 10004 10652 10056
rect 11980 10004 12032 10056
rect 5908 9911 5960 9920
rect 5908 9877 5917 9911
rect 5917 9877 5951 9911
rect 5951 9877 5960 9911
rect 5908 9868 5960 9877
rect 6184 9911 6236 9920
rect 6184 9877 6193 9911
rect 6193 9877 6227 9911
rect 6227 9877 6236 9911
rect 6184 9868 6236 9877
rect 11060 9936 11112 9988
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 16580 10047 16632 10056
rect 16580 10013 16589 10047
rect 16589 10013 16623 10047
rect 16623 10013 16632 10047
rect 16580 10004 16632 10013
rect 17316 10004 17368 10056
rect 10232 9868 10284 9920
rect 11980 9868 12032 9920
rect 12164 9868 12216 9920
rect 12532 9868 12584 9920
rect 15108 9868 15160 9920
rect 17500 9911 17552 9920
rect 17500 9877 17509 9911
rect 17509 9877 17543 9911
rect 17543 9877 17552 9911
rect 17500 9868 17552 9877
rect 2755 9766 2807 9818
rect 2819 9766 2871 9818
rect 2883 9766 2935 9818
rect 2947 9766 2999 9818
rect 3011 9766 3063 9818
rect 7470 9766 7522 9818
rect 7534 9766 7586 9818
rect 7598 9766 7650 9818
rect 7662 9766 7714 9818
rect 7726 9766 7778 9818
rect 12185 9766 12237 9818
rect 12249 9766 12301 9818
rect 12313 9766 12365 9818
rect 12377 9766 12429 9818
rect 12441 9766 12493 9818
rect 16900 9766 16952 9818
rect 16964 9766 17016 9818
rect 17028 9766 17080 9818
rect 17092 9766 17144 9818
rect 17156 9766 17208 9818
rect 2504 9664 2556 9716
rect 1032 9503 1084 9512
rect 1032 9469 1041 9503
rect 1041 9469 1075 9503
rect 1075 9469 1084 9503
rect 1032 9460 1084 9469
rect 4620 9460 4672 9512
rect 4804 9460 4856 9512
rect 6000 9596 6052 9648
rect 6828 9664 6880 9716
rect 9220 9664 9272 9716
rect 11796 9664 11848 9716
rect 13728 9664 13780 9716
rect 17776 9664 17828 9716
rect 18972 9664 19024 9716
rect 6552 9528 6604 9580
rect 13820 9596 13872 9648
rect 1124 9392 1176 9444
rect 5540 9460 5592 9512
rect 5724 9460 5776 9512
rect 6184 9503 6236 9512
rect 5264 9435 5316 9444
rect 5264 9401 5273 9435
rect 5273 9401 5307 9435
rect 5307 9401 5316 9435
rect 5264 9392 5316 9401
rect 4896 9324 4948 9376
rect 5448 9324 5500 9376
rect 5724 9324 5776 9376
rect 6184 9469 6193 9503
rect 6193 9469 6227 9503
rect 6227 9469 6236 9503
rect 6184 9460 6236 9469
rect 6736 9460 6788 9512
rect 7656 9460 7708 9512
rect 9128 9460 9180 9512
rect 10416 9460 10468 9512
rect 10692 9460 10744 9512
rect 11060 9503 11112 9512
rect 11060 9469 11069 9503
rect 11069 9469 11103 9503
rect 11103 9469 11112 9503
rect 11060 9460 11112 9469
rect 11336 9503 11388 9512
rect 11336 9469 11345 9503
rect 11345 9469 11379 9503
rect 11379 9469 11388 9503
rect 11336 9460 11388 9469
rect 11428 9503 11480 9512
rect 11428 9469 11437 9503
rect 11437 9469 11471 9503
rect 11471 9469 11480 9503
rect 11428 9460 11480 9469
rect 11612 9460 11664 9512
rect 12256 9503 12308 9512
rect 12256 9469 12265 9503
rect 12265 9469 12299 9503
rect 12299 9469 12308 9503
rect 12256 9460 12308 9469
rect 6184 9324 6236 9376
rect 10416 9367 10468 9376
rect 10416 9333 10425 9367
rect 10425 9333 10459 9367
rect 10459 9333 10468 9367
rect 10416 9324 10468 9333
rect 10784 9392 10836 9444
rect 11796 9392 11848 9444
rect 11980 9392 12032 9444
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 12716 9460 12768 9512
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 14280 9460 14332 9512
rect 13820 9392 13872 9444
rect 16672 9528 16724 9580
rect 17040 9503 17092 9512
rect 17040 9469 17049 9503
rect 17049 9469 17083 9503
rect 17083 9469 17092 9503
rect 17040 9460 17092 9469
rect 18788 9528 18840 9580
rect 13636 9324 13688 9376
rect 14004 9324 14056 9376
rect 14280 9367 14332 9376
rect 14280 9333 14289 9367
rect 14289 9333 14323 9367
rect 14323 9333 14332 9367
rect 14280 9324 14332 9333
rect 14464 9367 14516 9376
rect 14464 9333 14473 9367
rect 14473 9333 14507 9367
rect 14507 9333 14516 9367
rect 14464 9324 14516 9333
rect 15292 9392 15344 9444
rect 16764 9392 16816 9444
rect 15936 9324 15988 9376
rect 18236 9324 18288 9376
rect 5112 9222 5164 9274
rect 5176 9222 5228 9274
rect 5240 9222 5292 9274
rect 5304 9222 5356 9274
rect 5368 9222 5420 9274
rect 9827 9222 9879 9274
rect 9891 9222 9943 9274
rect 9955 9222 10007 9274
rect 10019 9222 10071 9274
rect 10083 9222 10135 9274
rect 14542 9222 14594 9274
rect 14606 9222 14658 9274
rect 14670 9222 14722 9274
rect 14734 9222 14786 9274
rect 14798 9222 14850 9274
rect 19257 9222 19309 9274
rect 19321 9222 19373 9274
rect 19385 9222 19437 9274
rect 19449 9222 19501 9274
rect 19513 9222 19565 9274
rect 1584 9120 1636 9172
rect 1952 9120 2004 9172
rect 3148 9120 3200 9172
rect 1032 8984 1084 9036
rect 1124 8984 1176 9036
rect 1492 8916 1544 8968
rect 1676 8984 1728 9036
rect 4160 9052 4212 9104
rect 4804 9120 4856 9172
rect 5540 9120 5592 9172
rect 5908 9120 5960 9172
rect 7196 9120 7248 9172
rect 9036 9120 9088 9172
rect 2596 8916 2648 8968
rect 4528 9027 4580 9036
rect 4528 8993 4537 9027
rect 4537 8993 4571 9027
rect 4571 8993 4580 9027
rect 4528 8984 4580 8993
rect 4804 9027 4856 9036
rect 4804 8993 4813 9027
rect 4813 8993 4847 9027
rect 4847 8993 4856 9027
rect 4804 8984 4856 8993
rect 4712 8916 4764 8968
rect 5356 9027 5408 9036
rect 5356 8993 5365 9027
rect 5365 8993 5399 9027
rect 5399 8993 5408 9027
rect 5356 8984 5408 8993
rect 5632 9027 5684 9036
rect 5632 8993 5641 9027
rect 5641 8993 5675 9027
rect 5675 8993 5684 9027
rect 5632 8984 5684 8993
rect 6276 8984 6328 9036
rect 7932 9052 7984 9104
rect 7104 8984 7156 9036
rect 7656 8984 7708 9036
rect 8760 8984 8812 9036
rect 9220 9027 9272 9036
rect 9220 8993 9229 9027
rect 9229 8993 9263 9027
rect 9263 8993 9272 9027
rect 9220 8984 9272 8993
rect 9588 9163 9640 9172
rect 9588 9129 9597 9163
rect 9597 9129 9631 9163
rect 9631 9129 9640 9163
rect 9588 9120 9640 9129
rect 11152 9120 11204 9172
rect 11336 9120 11388 9172
rect 11704 9120 11756 9172
rect 12532 9120 12584 9172
rect 12624 9120 12676 9172
rect 10324 8984 10376 9036
rect 5172 8848 5224 8900
rect 5448 8848 5500 8900
rect 9404 8848 9456 8900
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 5540 8780 5592 8832
rect 6000 8780 6052 8832
rect 6276 8780 6328 8832
rect 8852 8780 8904 8832
rect 9220 8780 9272 8832
rect 10416 8848 10468 8900
rect 10692 8984 10744 9036
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 11428 9052 11480 9104
rect 11520 8984 11572 9036
rect 11612 9027 11664 9036
rect 11612 8993 11621 9027
rect 11621 8993 11655 9027
rect 11655 8993 11664 9027
rect 11612 8984 11664 8993
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 11980 8984 12032 9036
rect 12440 9052 12492 9104
rect 12348 9027 12400 9036
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 14096 9120 14148 9172
rect 14280 9120 14332 9172
rect 14464 9120 14516 9172
rect 13544 9052 13596 9104
rect 13268 8984 13320 9036
rect 11060 8916 11112 8968
rect 13820 9027 13872 9036
rect 13820 8993 13829 9027
rect 13829 8993 13863 9027
rect 13863 8993 13872 9027
rect 13820 8984 13872 8993
rect 14096 8984 14148 9036
rect 13176 8848 13228 8900
rect 13728 8916 13780 8968
rect 14004 8916 14056 8968
rect 14280 8916 14332 8968
rect 15200 9052 15252 9104
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 16212 9120 16264 9172
rect 18512 9120 18564 9172
rect 17040 9052 17092 9104
rect 17316 9052 17368 9104
rect 16672 9027 16724 9036
rect 16672 8993 16681 9027
rect 16681 8993 16715 9027
rect 16715 8993 16724 9027
rect 16672 8984 16724 8993
rect 17868 8984 17920 9036
rect 18420 9027 18472 9036
rect 18420 8993 18429 9027
rect 18429 8993 18463 9027
rect 18463 8993 18472 9027
rect 18420 8984 18472 8993
rect 18512 9027 18564 9036
rect 18512 8993 18521 9027
rect 18521 8993 18555 9027
rect 18555 8993 18564 9027
rect 18512 8984 18564 8993
rect 15844 8916 15896 8968
rect 15936 8959 15988 8968
rect 15936 8925 15945 8959
rect 15945 8925 15979 8959
rect 15979 8925 15988 8959
rect 15936 8916 15988 8925
rect 12624 8780 12676 8832
rect 18696 8780 18748 8832
rect 2755 8678 2807 8730
rect 2819 8678 2871 8730
rect 2883 8678 2935 8730
rect 2947 8678 2999 8730
rect 3011 8678 3063 8730
rect 7470 8678 7522 8730
rect 7534 8678 7586 8730
rect 7598 8678 7650 8730
rect 7662 8678 7714 8730
rect 7726 8678 7778 8730
rect 12185 8678 12237 8730
rect 12249 8678 12301 8730
rect 12313 8678 12365 8730
rect 12377 8678 12429 8730
rect 12441 8678 12493 8730
rect 16900 8678 16952 8730
rect 16964 8678 17016 8730
rect 17028 8678 17080 8730
rect 17092 8678 17144 8730
rect 17156 8678 17208 8730
rect 1400 8576 1452 8628
rect 4712 8576 4764 8628
rect 5632 8576 5684 8628
rect 6000 8576 6052 8628
rect 8576 8576 8628 8628
rect 1032 8372 1084 8424
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 2596 8440 2648 8492
rect 1124 8304 1176 8356
rect 4620 8415 4672 8424
rect 4620 8381 4629 8415
rect 4629 8381 4663 8415
rect 4663 8381 4672 8415
rect 4620 8372 4672 8381
rect 1216 8236 1268 8288
rect 2044 8236 2096 8288
rect 4712 8236 4764 8288
rect 5172 8415 5224 8424
rect 5172 8381 5181 8415
rect 5181 8381 5215 8415
rect 5215 8381 5224 8415
rect 5172 8372 5224 8381
rect 9404 8576 9456 8628
rect 9588 8576 9640 8628
rect 11060 8576 11112 8628
rect 11612 8576 11664 8628
rect 11980 8576 12032 8628
rect 9312 8508 9364 8560
rect 9772 8551 9824 8560
rect 9772 8517 9781 8551
rect 9781 8517 9815 8551
rect 9815 8517 9824 8551
rect 9772 8508 9824 8517
rect 11336 8508 11388 8560
rect 17500 8576 17552 8628
rect 17776 8576 17828 8628
rect 5540 8372 5592 8424
rect 5908 8372 5960 8424
rect 6276 8415 6328 8424
rect 6276 8381 6310 8415
rect 6310 8381 6328 8415
rect 6276 8372 6328 8381
rect 7840 8372 7892 8424
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 11060 8440 11112 8492
rect 8668 8347 8720 8356
rect 8668 8313 8677 8347
rect 8677 8313 8711 8347
rect 8711 8313 8720 8347
rect 8668 8304 8720 8313
rect 5448 8236 5500 8288
rect 8484 8236 8536 8288
rect 8852 8372 8904 8424
rect 9220 8415 9272 8424
rect 9220 8381 9229 8415
rect 9229 8381 9263 8415
rect 9263 8381 9272 8415
rect 9220 8372 9272 8381
rect 9312 8415 9364 8424
rect 9312 8381 9321 8415
rect 9321 8381 9355 8415
rect 9355 8381 9364 8415
rect 9312 8372 9364 8381
rect 10140 8279 10192 8288
rect 10140 8245 10149 8279
rect 10149 8245 10183 8279
rect 10183 8245 10192 8279
rect 10140 8236 10192 8245
rect 10692 8304 10744 8356
rect 11244 8415 11296 8424
rect 11244 8381 11253 8415
rect 11253 8381 11287 8415
rect 11287 8381 11296 8415
rect 11244 8372 11296 8381
rect 16028 8508 16080 8560
rect 17316 8508 17368 8560
rect 12164 8483 12216 8492
rect 12164 8449 12173 8483
rect 12173 8449 12207 8483
rect 12207 8449 12216 8483
rect 12164 8440 12216 8449
rect 13084 8440 13136 8492
rect 11612 8415 11664 8424
rect 11612 8381 11645 8415
rect 11645 8381 11664 8415
rect 11612 8372 11664 8381
rect 11796 8372 11848 8424
rect 11888 8372 11940 8424
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 12532 8415 12584 8424
rect 12532 8381 12541 8415
rect 12541 8381 12575 8415
rect 12575 8381 12584 8415
rect 12532 8372 12584 8381
rect 13268 8372 13320 8424
rect 15476 8440 15528 8492
rect 13636 8372 13688 8424
rect 14188 8372 14240 8424
rect 14924 8372 14976 8424
rect 15200 8372 15252 8424
rect 16028 8415 16080 8424
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 16028 8372 16080 8381
rect 16304 8415 16356 8424
rect 16304 8381 16313 8415
rect 16313 8381 16347 8415
rect 16347 8381 16356 8415
rect 16304 8372 16356 8381
rect 16672 8440 16724 8492
rect 17684 8440 17736 8492
rect 17960 8440 18012 8492
rect 18144 8440 18196 8492
rect 17868 8415 17920 8424
rect 17868 8381 17877 8415
rect 17877 8381 17911 8415
rect 17911 8381 17920 8415
rect 17868 8372 17920 8381
rect 18236 8415 18288 8424
rect 18236 8381 18245 8415
rect 18245 8381 18279 8415
rect 18279 8381 18288 8415
rect 18236 8372 18288 8381
rect 10416 8236 10468 8288
rect 10968 8236 11020 8288
rect 11428 8236 11480 8288
rect 11980 8236 12032 8288
rect 12164 8236 12216 8288
rect 14004 8304 14056 8356
rect 15568 8304 15620 8356
rect 16672 8347 16724 8356
rect 16672 8313 16681 8347
rect 16681 8313 16715 8347
rect 16715 8313 16724 8347
rect 16672 8304 16724 8313
rect 17960 8347 18012 8356
rect 17960 8313 17969 8347
rect 17969 8313 18003 8347
rect 18003 8313 18012 8347
rect 17960 8304 18012 8313
rect 18052 8347 18104 8356
rect 18052 8313 18061 8347
rect 18061 8313 18095 8347
rect 18095 8313 18104 8347
rect 18052 8304 18104 8313
rect 18512 8304 18564 8356
rect 13820 8236 13872 8288
rect 13912 8236 13964 8288
rect 14464 8236 14516 8288
rect 14924 8279 14976 8288
rect 14924 8245 14933 8279
rect 14933 8245 14967 8279
rect 14967 8245 14976 8279
rect 14924 8236 14976 8245
rect 16396 8236 16448 8288
rect 18696 8236 18748 8288
rect 5112 8134 5164 8186
rect 5176 8134 5228 8186
rect 5240 8134 5292 8186
rect 5304 8134 5356 8186
rect 5368 8134 5420 8186
rect 9827 8134 9879 8186
rect 9891 8134 9943 8186
rect 9955 8134 10007 8186
rect 10019 8134 10071 8186
rect 10083 8134 10135 8186
rect 14542 8134 14594 8186
rect 14606 8134 14658 8186
rect 14670 8134 14722 8186
rect 14734 8134 14786 8186
rect 14798 8134 14850 8186
rect 19257 8134 19309 8186
rect 19321 8134 19373 8186
rect 19385 8134 19437 8186
rect 19449 8134 19501 8186
rect 19513 8134 19565 8186
rect 1216 8075 1268 8084
rect 1216 8041 1225 8075
rect 1225 8041 1259 8075
rect 1259 8041 1268 8075
rect 1216 8032 1268 8041
rect 1676 8032 1728 8084
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 1584 7896 1636 7948
rect 3332 8032 3384 8084
rect 4620 8032 4672 8084
rect 4528 7964 4580 8016
rect 940 7803 992 7812
rect 940 7769 949 7803
rect 949 7769 983 7803
rect 983 7769 992 7803
rect 940 7760 992 7769
rect 1308 7760 1360 7812
rect 2044 7828 2096 7880
rect 3148 7939 3200 7948
rect 3148 7905 3157 7939
rect 3157 7905 3191 7939
rect 3191 7905 3200 7939
rect 3148 7896 3200 7905
rect 5540 8032 5592 8084
rect 5724 8032 5776 8084
rect 7288 8007 7340 8016
rect 7288 7973 7322 8007
rect 7322 7973 7340 8007
rect 7288 7964 7340 7973
rect 9036 8032 9088 8084
rect 9404 8032 9456 8084
rect 9588 8032 9640 8084
rect 10048 8032 10100 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 11060 7964 11112 8016
rect 11336 7964 11388 8016
rect 3240 7828 3292 7880
rect 4528 7828 4580 7880
rect 4712 7828 4764 7880
rect 5448 7939 5500 7948
rect 5448 7905 5457 7939
rect 5457 7905 5491 7939
rect 5491 7905 5500 7939
rect 5448 7896 5500 7905
rect 7104 7896 7156 7948
rect 8944 7939 8996 7948
rect 8944 7905 8953 7939
rect 8953 7905 8987 7939
rect 8987 7905 8996 7939
rect 8944 7896 8996 7905
rect 2136 7760 2188 7812
rect 4068 7760 4120 7812
rect 4344 7692 4396 7744
rect 4528 7735 4580 7744
rect 4528 7701 4537 7735
rect 4537 7701 4571 7735
rect 4571 7701 4580 7735
rect 4528 7692 4580 7701
rect 4896 7760 4948 7812
rect 8852 7828 8904 7880
rect 10048 7939 10100 7948
rect 10048 7905 10057 7939
rect 10057 7905 10091 7939
rect 10091 7905 10100 7939
rect 10048 7896 10100 7905
rect 6276 7760 6328 7812
rect 9128 7760 9180 7812
rect 9496 7760 9548 7812
rect 9588 7760 9640 7812
rect 9956 7828 10008 7880
rect 10416 7896 10468 7948
rect 10968 7828 11020 7880
rect 11704 7896 11756 7948
rect 11888 7896 11940 7948
rect 12348 8075 12400 8084
rect 12348 8041 12357 8075
rect 12357 8041 12391 8075
rect 12391 8041 12400 8075
rect 12348 8032 12400 8041
rect 12624 8032 12676 8084
rect 12164 7964 12216 8016
rect 12440 7964 12492 8016
rect 13084 8032 13136 8084
rect 14924 8032 14976 8084
rect 15108 8032 15160 8084
rect 11336 7760 11388 7812
rect 11796 7828 11848 7880
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 12808 7896 12860 7905
rect 13084 7939 13136 7948
rect 13084 7905 13093 7939
rect 13093 7905 13127 7939
rect 13127 7905 13136 7939
rect 13084 7896 13136 7905
rect 13452 7828 13504 7880
rect 14004 7896 14056 7948
rect 14188 7896 14240 7948
rect 13912 7871 13964 7880
rect 13912 7837 13921 7871
rect 13921 7837 13955 7871
rect 13955 7837 13964 7871
rect 13912 7828 13964 7837
rect 12256 7760 12308 7812
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 10784 7692 10836 7744
rect 11152 7692 11204 7744
rect 11520 7692 11572 7744
rect 11704 7692 11756 7744
rect 12164 7692 12216 7744
rect 12716 7760 12768 7812
rect 13268 7760 13320 7812
rect 14004 7735 14056 7744
rect 14004 7701 14013 7735
rect 14013 7701 14047 7735
rect 14047 7701 14056 7735
rect 14004 7692 14056 7701
rect 16580 8075 16632 8084
rect 16580 8041 16589 8075
rect 16589 8041 16623 8075
rect 16623 8041 16632 8075
rect 16580 8032 16632 8041
rect 14556 7896 14608 7948
rect 14924 7939 14976 7948
rect 14924 7905 14933 7939
rect 14933 7905 14967 7939
rect 14967 7905 14976 7939
rect 14924 7896 14976 7905
rect 15016 7828 15068 7880
rect 15568 7939 15620 7948
rect 15568 7905 15577 7939
rect 15577 7905 15611 7939
rect 15611 7905 15620 7939
rect 15568 7896 15620 7905
rect 15660 7939 15712 7948
rect 15660 7905 15669 7939
rect 15669 7905 15703 7939
rect 15703 7905 15712 7939
rect 15660 7896 15712 7905
rect 17316 7964 17368 8016
rect 18972 7964 19024 8016
rect 16212 7896 16264 7948
rect 17224 7939 17276 7948
rect 17224 7905 17233 7939
rect 17233 7905 17267 7939
rect 17267 7905 17276 7939
rect 17224 7896 17276 7905
rect 17684 7896 17736 7948
rect 18512 7896 18564 7948
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 15844 7760 15896 7812
rect 18052 7760 18104 7812
rect 15384 7692 15436 7744
rect 16396 7735 16448 7744
rect 16396 7701 16405 7735
rect 16405 7701 16439 7735
rect 16439 7701 16448 7735
rect 16396 7692 16448 7701
rect 2755 7590 2807 7642
rect 2819 7590 2871 7642
rect 2883 7590 2935 7642
rect 2947 7590 2999 7642
rect 3011 7590 3063 7642
rect 7470 7590 7522 7642
rect 7534 7590 7586 7642
rect 7598 7590 7650 7642
rect 7662 7590 7714 7642
rect 7726 7590 7778 7642
rect 12185 7590 12237 7642
rect 12249 7590 12301 7642
rect 12313 7590 12365 7642
rect 12377 7590 12429 7642
rect 12441 7590 12493 7642
rect 16900 7590 16952 7642
rect 16964 7590 17016 7642
rect 17028 7590 17080 7642
rect 17092 7590 17144 7642
rect 17156 7590 17208 7642
rect 1032 7531 1084 7540
rect 1032 7497 1041 7531
rect 1041 7497 1075 7531
rect 1075 7497 1084 7531
rect 1032 7488 1084 7497
rect 1584 7488 1636 7540
rect 2136 7531 2188 7540
rect 2136 7497 2145 7531
rect 2145 7497 2179 7531
rect 2179 7497 2188 7531
rect 2136 7488 2188 7497
rect 2596 7488 2648 7540
rect 2872 7488 2924 7540
rect 3332 7488 3384 7540
rect 2596 7284 2648 7336
rect 4528 7420 4580 7472
rect 4068 7352 4120 7404
rect 4160 7352 4212 7404
rect 5908 7488 5960 7540
rect 8208 7488 8260 7540
rect 10508 7488 10560 7540
rect 11244 7488 11296 7540
rect 11336 7488 11388 7540
rect 12440 7488 12492 7540
rect 12716 7488 12768 7540
rect 13728 7488 13780 7540
rect 14004 7488 14056 7540
rect 14188 7488 14240 7540
rect 4896 7327 4948 7336
rect 4896 7293 4905 7327
rect 4905 7293 4939 7327
rect 4939 7293 4948 7327
rect 4896 7284 4948 7293
rect 5632 7284 5684 7336
rect 6000 7284 6052 7336
rect 2044 7148 2096 7200
rect 3240 7216 3292 7268
rect 4988 7216 5040 7268
rect 5448 7216 5500 7268
rect 2872 7148 2924 7200
rect 3148 7148 3200 7200
rect 4896 7148 4948 7200
rect 6552 7284 6604 7336
rect 7104 7352 7156 7404
rect 8484 7352 8536 7404
rect 6460 7148 6512 7200
rect 10416 7420 10468 7472
rect 8024 7148 8076 7200
rect 8576 7191 8628 7200
rect 8576 7157 8585 7191
rect 8585 7157 8619 7191
rect 8619 7157 8628 7191
rect 8576 7148 8628 7157
rect 8852 7216 8904 7268
rect 9036 7216 9088 7268
rect 10048 7284 10100 7336
rect 10232 7284 10284 7336
rect 12900 7420 12952 7472
rect 11796 7352 11848 7404
rect 11980 7352 12032 7404
rect 9588 7191 9640 7200
rect 9588 7157 9597 7191
rect 9597 7157 9631 7191
rect 9631 7157 9640 7191
rect 9588 7148 9640 7157
rect 9956 7216 10008 7268
rect 10968 7284 11020 7336
rect 11244 7327 11296 7336
rect 11244 7293 11253 7327
rect 11253 7293 11287 7327
rect 11287 7293 11296 7327
rect 11244 7284 11296 7293
rect 11520 7284 11572 7336
rect 11152 7216 11204 7268
rect 9864 7148 9916 7200
rect 10416 7148 10468 7200
rect 11704 7327 11756 7336
rect 11704 7293 11713 7327
rect 11713 7293 11747 7327
rect 11747 7293 11756 7327
rect 11704 7284 11756 7293
rect 11888 7284 11940 7336
rect 12532 7352 12584 7404
rect 12992 7352 13044 7404
rect 13268 7352 13320 7404
rect 14556 7420 14608 7472
rect 14924 7420 14976 7472
rect 14188 7352 14240 7404
rect 15200 7488 15252 7540
rect 16304 7531 16356 7540
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 18512 7488 18564 7540
rect 18880 7531 18932 7540
rect 18880 7497 18889 7531
rect 18889 7497 18923 7531
rect 18923 7497 18932 7531
rect 18880 7488 18932 7497
rect 15844 7352 15896 7404
rect 18696 7352 18748 7404
rect 12532 7148 12584 7200
rect 12808 7148 12860 7200
rect 13820 7216 13872 7268
rect 14464 7216 14516 7268
rect 16304 7284 16356 7336
rect 17224 7284 17276 7336
rect 17684 7284 17736 7336
rect 17868 7327 17920 7336
rect 17868 7293 17877 7327
rect 17877 7293 17911 7327
rect 17911 7293 17920 7327
rect 17868 7284 17920 7293
rect 18604 7148 18656 7200
rect 5112 7046 5164 7098
rect 5176 7046 5228 7098
rect 5240 7046 5292 7098
rect 5304 7046 5356 7098
rect 5368 7046 5420 7098
rect 9827 7046 9879 7098
rect 9891 7046 9943 7098
rect 9955 7046 10007 7098
rect 10019 7046 10071 7098
rect 10083 7046 10135 7098
rect 14542 7046 14594 7098
rect 14606 7046 14658 7098
rect 14670 7046 14722 7098
rect 14734 7046 14786 7098
rect 14798 7046 14850 7098
rect 19257 7046 19309 7098
rect 19321 7046 19373 7098
rect 19385 7046 19437 7098
rect 19449 7046 19501 7098
rect 19513 7046 19565 7098
rect 3240 6944 3292 6996
rect 4068 6944 4120 6996
rect 5172 6944 5224 6996
rect 1124 6851 1176 6860
rect 1124 6817 1133 6851
rect 1133 6817 1167 6851
rect 1167 6817 1176 6851
rect 1124 6808 1176 6817
rect 1216 6808 1268 6860
rect 1492 6808 1544 6860
rect 2596 6808 2648 6860
rect 8392 6944 8444 6996
rect 4896 6876 4948 6928
rect 940 6672 992 6724
rect 1400 6672 1452 6724
rect 3516 6672 3568 6724
rect 1124 6604 1176 6656
rect 1584 6604 1636 6656
rect 3148 6604 3200 6656
rect 4160 6851 4212 6860
rect 4160 6817 4169 6851
rect 4169 6817 4203 6851
rect 4203 6817 4212 6851
rect 4160 6808 4212 6817
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 6184 6851 6236 6860
rect 6184 6817 6218 6851
rect 6218 6817 6236 6851
rect 6184 6808 6236 6817
rect 8024 6876 8076 6928
rect 9680 6876 9732 6928
rect 4436 6604 4488 6656
rect 5448 6604 5500 6656
rect 5540 6647 5592 6656
rect 5540 6613 5549 6647
rect 5549 6613 5583 6647
rect 5583 6613 5592 6647
rect 5540 6604 5592 6613
rect 6920 6740 6972 6792
rect 7380 6808 7432 6860
rect 8392 6851 8444 6860
rect 8392 6817 8401 6851
rect 8401 6817 8435 6851
rect 8435 6817 8444 6851
rect 8392 6808 8444 6817
rect 8484 6808 8536 6860
rect 8944 6808 8996 6860
rect 9128 6808 9180 6860
rect 9404 6851 9456 6860
rect 9404 6817 9413 6851
rect 9413 6817 9447 6851
rect 9447 6817 9456 6851
rect 9404 6808 9456 6817
rect 7104 6672 7156 6724
rect 9588 6740 9640 6792
rect 9220 6672 9272 6724
rect 10232 6851 10284 6860
rect 10232 6817 10241 6851
rect 10241 6817 10275 6851
rect 10275 6817 10284 6851
rect 10232 6808 10284 6817
rect 10968 6808 11020 6860
rect 11704 6876 11756 6928
rect 11244 6740 11296 6792
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 9404 6604 9456 6656
rect 11152 6604 11204 6656
rect 11244 6604 11296 6656
rect 12624 6944 12676 6996
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 12808 6808 12860 6860
rect 12900 6808 12952 6860
rect 13268 6808 13320 6860
rect 11888 6740 11940 6792
rect 11980 6740 12032 6792
rect 12716 6740 12768 6792
rect 13912 6944 13964 6996
rect 17500 6987 17552 6996
rect 17500 6953 17509 6987
rect 17509 6953 17543 6987
rect 17543 6953 17552 6987
rect 17500 6944 17552 6953
rect 13176 6604 13228 6656
rect 13268 6604 13320 6656
rect 16212 6876 16264 6928
rect 18052 6876 18104 6928
rect 14464 6808 14516 6860
rect 15200 6808 15252 6860
rect 16672 6808 16724 6860
rect 18604 6851 18656 6860
rect 18604 6817 18622 6851
rect 18622 6817 18656 6851
rect 18604 6808 18656 6817
rect 18972 6808 19024 6860
rect 13636 6783 13688 6792
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 15016 6647 15068 6656
rect 15016 6613 15025 6647
rect 15025 6613 15059 6647
rect 15059 6613 15068 6647
rect 15016 6604 15068 6613
rect 2755 6502 2807 6554
rect 2819 6502 2871 6554
rect 2883 6502 2935 6554
rect 2947 6502 2999 6554
rect 3011 6502 3063 6554
rect 7470 6502 7522 6554
rect 7534 6502 7586 6554
rect 7598 6502 7650 6554
rect 7662 6502 7714 6554
rect 7726 6502 7778 6554
rect 12185 6502 12237 6554
rect 12249 6502 12301 6554
rect 12313 6502 12365 6554
rect 12377 6502 12429 6554
rect 12441 6502 12493 6554
rect 16900 6502 16952 6554
rect 16964 6502 17016 6554
rect 17028 6502 17080 6554
rect 17092 6502 17144 6554
rect 17156 6502 17208 6554
rect 1032 6332 1084 6384
rect 1400 6400 1452 6452
rect 940 6196 992 6248
rect 1308 6239 1360 6248
rect 1308 6205 1317 6239
rect 1317 6205 1351 6239
rect 1351 6205 1360 6239
rect 1308 6196 1360 6205
rect 1584 6239 1636 6248
rect 1584 6205 1593 6239
rect 1593 6205 1627 6239
rect 1627 6205 1636 6239
rect 1584 6196 1636 6205
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 3240 6400 3292 6452
rect 3516 6400 3568 6452
rect 5540 6400 5592 6452
rect 5448 6332 5500 6384
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3148 6196 3200 6248
rect 3976 6239 4028 6248
rect 3976 6205 3977 6239
rect 3977 6205 4011 6239
rect 4011 6205 4028 6239
rect 3976 6196 4028 6205
rect 4896 6196 4948 6248
rect 5172 6196 5224 6248
rect 7104 6400 7156 6452
rect 9128 6400 9180 6452
rect 9588 6400 9640 6452
rect 10416 6400 10468 6452
rect 12164 6400 12216 6452
rect 12532 6400 12584 6452
rect 15752 6400 15804 6452
rect 16488 6400 16540 6452
rect 18144 6443 18196 6452
rect 18144 6409 18153 6443
rect 18153 6409 18187 6443
rect 18187 6409 18196 6443
rect 18144 6400 18196 6409
rect 9312 6332 9364 6384
rect 10968 6375 11020 6384
rect 4252 6171 4304 6180
rect 4252 6137 4261 6171
rect 4261 6137 4295 6171
rect 4295 6137 4304 6171
rect 4252 6128 4304 6137
rect 5724 6196 5776 6248
rect 10968 6341 10977 6375
rect 10977 6341 11011 6375
rect 11011 6341 11020 6375
rect 10968 6332 11020 6341
rect 13820 6332 13872 6384
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 6552 6196 6604 6248
rect 7380 6196 7432 6248
rect 9588 6264 9640 6316
rect 10784 6264 10836 6316
rect 5908 6171 5960 6180
rect 5908 6137 5917 6171
rect 5917 6137 5951 6171
rect 5951 6137 5960 6171
rect 5908 6128 5960 6137
rect 8392 6196 8444 6248
rect 7840 6128 7892 6180
rect 9680 6196 9732 6248
rect 11520 6264 11572 6316
rect 11980 6264 12032 6316
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 13452 6264 13504 6316
rect 1216 6060 1268 6112
rect 1308 6060 1360 6112
rect 2596 6060 2648 6112
rect 5448 6060 5500 6112
rect 7012 6060 7064 6112
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 8576 6060 8628 6112
rect 9404 6128 9456 6180
rect 11888 6239 11940 6248
rect 11888 6205 11897 6239
rect 11897 6205 11931 6239
rect 11931 6205 11940 6239
rect 11888 6196 11940 6205
rect 12992 6196 13044 6248
rect 13636 6196 13688 6248
rect 13912 6196 13964 6248
rect 9588 6060 9640 6112
rect 11612 6128 11664 6180
rect 11796 6128 11848 6180
rect 12624 6128 12676 6180
rect 12808 6128 12860 6180
rect 14464 6239 14516 6248
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 15476 6332 15528 6384
rect 15568 6264 15620 6316
rect 13268 6060 13320 6112
rect 14464 6060 14516 6112
rect 15200 6060 15252 6112
rect 15568 6171 15620 6180
rect 15568 6137 15577 6171
rect 15577 6137 15611 6171
rect 15611 6137 15620 6171
rect 15568 6128 15620 6137
rect 15752 6239 15804 6248
rect 15752 6205 15761 6239
rect 15761 6205 15795 6239
rect 15795 6205 15804 6239
rect 15752 6196 15804 6205
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 16120 6264 16172 6316
rect 16672 6239 16724 6248
rect 16672 6205 16681 6239
rect 16681 6205 16715 6239
rect 16715 6205 16724 6239
rect 16672 6196 16724 6205
rect 17224 6239 17276 6248
rect 17224 6205 17233 6239
rect 17233 6205 17267 6239
rect 17267 6205 17276 6239
rect 17224 6196 17276 6205
rect 17776 6239 17828 6248
rect 17776 6205 17785 6239
rect 17785 6205 17819 6239
rect 17819 6205 17828 6239
rect 17776 6196 17828 6205
rect 18604 6264 18656 6316
rect 18328 6239 18380 6248
rect 18328 6205 18337 6239
rect 18337 6205 18371 6239
rect 18371 6205 18380 6239
rect 18328 6196 18380 6205
rect 18420 6196 18472 6248
rect 5112 5958 5164 6010
rect 5176 5958 5228 6010
rect 5240 5958 5292 6010
rect 5304 5958 5356 6010
rect 5368 5958 5420 6010
rect 9827 5958 9879 6010
rect 9891 5958 9943 6010
rect 9955 5958 10007 6010
rect 10019 5958 10071 6010
rect 10083 5958 10135 6010
rect 14542 5958 14594 6010
rect 14606 5958 14658 6010
rect 14670 5958 14722 6010
rect 14734 5958 14786 6010
rect 14798 5958 14850 6010
rect 19257 5958 19309 6010
rect 19321 5958 19373 6010
rect 19385 5958 19437 6010
rect 19449 5958 19501 6010
rect 19513 5958 19565 6010
rect 1308 5856 1360 5908
rect 1860 5856 1912 5908
rect 1952 5856 2004 5908
rect 3332 5856 3384 5908
rect 6368 5899 6420 5908
rect 6368 5865 6377 5899
rect 6377 5865 6411 5899
rect 6411 5865 6420 5899
rect 6368 5856 6420 5865
rect 6828 5856 6880 5908
rect 8208 5856 8260 5908
rect 8852 5856 8904 5908
rect 8944 5856 8996 5908
rect 1216 5652 1268 5704
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 4896 5788 4948 5840
rect 1860 5720 1912 5729
rect 3424 5763 3476 5772
rect 3424 5729 3458 5763
rect 3458 5729 3476 5763
rect 3424 5720 3476 5729
rect 4160 5720 4212 5772
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 1952 5559 2004 5568
rect 1952 5525 1961 5559
rect 1961 5525 1995 5559
rect 1995 5525 2004 5559
rect 1952 5516 2004 5525
rect 4436 5652 4488 5704
rect 5724 5720 5776 5772
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 6736 5720 6788 5772
rect 6828 5720 6880 5772
rect 7104 5720 7156 5772
rect 8484 5763 8536 5772
rect 8484 5729 8493 5763
rect 8493 5729 8527 5763
rect 8527 5729 8536 5763
rect 8484 5720 8536 5729
rect 8576 5720 8628 5772
rect 9404 5856 9456 5908
rect 10784 5856 10836 5908
rect 6092 5652 6144 5704
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 9404 5763 9456 5772
rect 9404 5729 9413 5763
rect 9413 5729 9447 5763
rect 9447 5729 9456 5763
rect 9404 5720 9456 5729
rect 11704 5856 11756 5908
rect 12440 5856 12492 5908
rect 12532 5856 12584 5908
rect 13912 5856 13964 5908
rect 14280 5856 14332 5908
rect 12164 5788 12216 5840
rect 14188 5788 14240 5840
rect 11336 5763 11388 5772
rect 11336 5729 11345 5763
rect 11345 5729 11379 5763
rect 11379 5729 11388 5763
rect 11336 5720 11388 5729
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 11060 5652 11112 5704
rect 11980 5720 12032 5772
rect 14280 5720 14332 5772
rect 15016 5856 15068 5908
rect 15568 5856 15620 5908
rect 15660 5856 15712 5908
rect 15752 5856 15804 5908
rect 17500 5856 17552 5908
rect 17776 5856 17828 5908
rect 14740 5831 14792 5840
rect 14740 5797 14749 5831
rect 14749 5797 14783 5831
rect 14783 5797 14792 5831
rect 14740 5788 14792 5797
rect 15292 5788 15344 5840
rect 15108 5720 15160 5772
rect 9680 5627 9732 5636
rect 9680 5593 9689 5627
rect 9689 5593 9723 5627
rect 9723 5593 9732 5627
rect 9680 5584 9732 5593
rect 10600 5584 10652 5636
rect 10968 5584 11020 5636
rect 3516 5516 3568 5568
rect 4068 5516 4120 5568
rect 7932 5516 7984 5568
rect 9036 5559 9088 5568
rect 9036 5525 9045 5559
rect 9045 5525 9079 5559
rect 9079 5525 9088 5559
rect 9036 5516 9088 5525
rect 9312 5516 9364 5568
rect 9404 5516 9456 5568
rect 10508 5516 10560 5568
rect 10692 5516 10744 5568
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 15660 5720 15712 5772
rect 16304 5763 16356 5772
rect 16304 5729 16313 5763
rect 16313 5729 16347 5763
rect 16347 5729 16356 5763
rect 16304 5720 16356 5729
rect 16488 5763 16540 5772
rect 16488 5729 16497 5763
rect 16497 5729 16531 5763
rect 16531 5729 16540 5763
rect 16488 5720 16540 5729
rect 17224 5788 17276 5840
rect 18328 5856 18380 5908
rect 17408 5763 17460 5772
rect 17408 5729 17417 5763
rect 17417 5729 17451 5763
rect 17451 5729 17460 5763
rect 17408 5720 17460 5729
rect 18144 5720 18196 5772
rect 18328 5720 18380 5772
rect 18512 5763 18564 5772
rect 18512 5729 18521 5763
rect 18521 5729 18555 5763
rect 18555 5729 18564 5763
rect 18512 5720 18564 5729
rect 11796 5584 11848 5636
rect 15384 5516 15436 5568
rect 16120 5559 16172 5568
rect 16120 5525 16129 5559
rect 16129 5525 16163 5559
rect 16163 5525 16172 5559
rect 16120 5516 16172 5525
rect 2755 5414 2807 5466
rect 2819 5414 2871 5466
rect 2883 5414 2935 5466
rect 2947 5414 2999 5466
rect 3011 5414 3063 5466
rect 7470 5414 7522 5466
rect 7534 5414 7586 5466
rect 7598 5414 7650 5466
rect 7662 5414 7714 5466
rect 7726 5414 7778 5466
rect 12185 5414 12237 5466
rect 12249 5414 12301 5466
rect 12313 5414 12365 5466
rect 12377 5414 12429 5466
rect 12441 5414 12493 5466
rect 16900 5414 16952 5466
rect 16964 5414 17016 5466
rect 17028 5414 17080 5466
rect 17092 5414 17144 5466
rect 17156 5414 17208 5466
rect 1492 5312 1544 5364
rect 1860 5312 1912 5364
rect 7840 5312 7892 5364
rect 7932 5312 7984 5364
rect 9404 5312 9456 5364
rect 9496 5355 9548 5364
rect 9496 5321 9505 5355
rect 9505 5321 9539 5355
rect 9539 5321 9548 5355
rect 9496 5312 9548 5321
rect 6736 5244 6788 5296
rect 10784 5312 10836 5364
rect 10876 5312 10928 5364
rect 9864 5244 9916 5296
rect 10600 5244 10652 5296
rect 11336 5244 11388 5296
rect 11980 5244 12032 5296
rect 12072 5244 12124 5296
rect 13360 5312 13412 5364
rect 14096 5355 14148 5364
rect 14096 5321 14105 5355
rect 14105 5321 14139 5355
rect 14139 5321 14148 5355
rect 14096 5312 14148 5321
rect 14372 5312 14424 5364
rect 14464 5312 14516 5364
rect 1400 5176 1452 5228
rect 3056 5176 3108 5228
rect 8024 5176 8076 5228
rect 1216 5151 1268 5160
rect 1216 5117 1225 5151
rect 1225 5117 1259 5151
rect 1259 5117 1268 5151
rect 1216 5108 1268 5117
rect 1308 5151 1360 5160
rect 1308 5117 1317 5151
rect 1317 5117 1351 5151
rect 1351 5117 1360 5151
rect 1308 5108 1360 5117
rect 4252 5108 4304 5160
rect 4988 5108 5040 5160
rect 5448 5151 5500 5160
rect 5448 5117 5482 5151
rect 5482 5117 5500 5151
rect 5448 5108 5500 5117
rect 1952 5083 2004 5092
rect 1952 5049 1986 5083
rect 1986 5049 2004 5083
rect 1952 5040 2004 5049
rect 4068 5040 4120 5092
rect 1584 4972 1636 5024
rect 9036 5040 9088 5092
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 9864 5083 9916 5092
rect 9864 5049 9873 5083
rect 9873 5049 9907 5083
rect 9907 5049 9916 5083
rect 9864 5040 9916 5049
rect 9588 4972 9640 5024
rect 10232 5108 10284 5160
rect 10416 5151 10468 5160
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 10508 5108 10560 5160
rect 10600 5083 10652 5092
rect 10600 5049 10609 5083
rect 10609 5049 10643 5083
rect 10643 5049 10652 5083
rect 10600 5040 10652 5049
rect 10692 4972 10744 5024
rect 11060 5108 11112 5160
rect 11704 5108 11756 5160
rect 12072 5108 12124 5160
rect 13820 5244 13872 5296
rect 15200 5176 15252 5228
rect 16120 5176 16172 5228
rect 11244 5040 11296 5092
rect 11796 5040 11848 5092
rect 12440 5040 12492 5092
rect 12532 5083 12584 5092
rect 12532 5049 12541 5083
rect 12541 5049 12575 5083
rect 12575 5049 12584 5083
rect 12532 5040 12584 5049
rect 12900 5040 12952 5092
rect 13820 5108 13872 5160
rect 14372 5108 14424 5160
rect 14740 5108 14792 5160
rect 15292 5151 15344 5160
rect 15292 5117 15301 5151
rect 15301 5117 15335 5151
rect 15335 5117 15344 5151
rect 15292 5108 15344 5117
rect 15384 5108 15436 5160
rect 18052 5108 18104 5160
rect 16304 5040 16356 5092
rect 17408 5040 17460 5092
rect 13820 4972 13872 5024
rect 14464 5015 14516 5024
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14464 4972 14516 4981
rect 16764 5015 16816 5024
rect 16764 4981 16773 5015
rect 16773 4981 16807 5015
rect 16807 4981 16816 5015
rect 16764 4972 16816 4981
rect 18144 4972 18196 5024
rect 18788 5015 18840 5024
rect 18788 4981 18797 5015
rect 18797 4981 18831 5015
rect 18831 4981 18840 5015
rect 18788 4972 18840 4981
rect 5112 4870 5164 4922
rect 5176 4870 5228 4922
rect 5240 4870 5292 4922
rect 5304 4870 5356 4922
rect 5368 4870 5420 4922
rect 9827 4870 9879 4922
rect 9891 4870 9943 4922
rect 9955 4870 10007 4922
rect 10019 4870 10071 4922
rect 10083 4870 10135 4922
rect 14542 4870 14594 4922
rect 14606 4870 14658 4922
rect 14670 4870 14722 4922
rect 14734 4870 14786 4922
rect 14798 4870 14850 4922
rect 19257 4870 19309 4922
rect 19321 4870 19373 4922
rect 19385 4870 19437 4922
rect 19449 4870 19501 4922
rect 19513 4870 19565 4922
rect 1308 4768 1360 4820
rect 1676 4768 1728 4820
rect 5816 4768 5868 4820
rect 8484 4768 8536 4820
rect 10416 4768 10468 4820
rect 10968 4768 11020 4820
rect 12348 4768 12400 4820
rect 14372 4768 14424 4820
rect 16028 4768 16080 4820
rect 16764 4768 16816 4820
rect 1400 4632 1452 4684
rect 1492 4675 1544 4684
rect 1492 4641 1501 4675
rect 1501 4641 1535 4675
rect 1535 4641 1544 4675
rect 1492 4632 1544 4641
rect 4436 4632 4488 4684
rect 6368 4675 6420 4684
rect 6368 4641 6402 4675
rect 6402 4641 6420 4675
rect 6368 4632 6420 4641
rect 10692 4700 10744 4752
rect 11336 4700 11388 4752
rect 12072 4700 12124 4752
rect 12624 4700 12676 4752
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 1124 4471 1176 4480
rect 1124 4437 1133 4471
rect 1133 4437 1167 4471
rect 1167 4437 1176 4471
rect 1124 4428 1176 4437
rect 2596 4428 2648 4480
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 8392 4428 8444 4480
rect 9036 4428 9088 4480
rect 10508 4675 10560 4684
rect 10508 4641 10526 4675
rect 10526 4641 10560 4675
rect 10508 4632 10560 4641
rect 10968 4675 11020 4684
rect 10968 4641 10977 4675
rect 10977 4641 11011 4675
rect 11011 4641 11020 4675
rect 10968 4632 11020 4641
rect 11060 4675 11112 4684
rect 11060 4641 11069 4675
rect 11069 4641 11103 4675
rect 11103 4641 11112 4675
rect 11060 4632 11112 4641
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 11428 4632 11480 4641
rect 10784 4607 10836 4616
rect 10784 4573 10793 4607
rect 10793 4573 10827 4607
rect 10827 4573 10836 4607
rect 10784 4564 10836 4573
rect 11612 4632 11664 4684
rect 12348 4675 12400 4684
rect 12348 4641 12357 4675
rect 12357 4641 12391 4675
rect 12391 4641 12400 4675
rect 12348 4632 12400 4641
rect 15384 4632 15436 4684
rect 16488 4632 16540 4684
rect 17408 4743 17460 4752
rect 17408 4709 17417 4743
rect 17417 4709 17451 4743
rect 17451 4709 17460 4743
rect 17408 4700 17460 4709
rect 18512 4768 18564 4820
rect 18972 4700 19024 4752
rect 12992 4564 13044 4616
rect 13084 4496 13136 4548
rect 11612 4428 11664 4480
rect 16764 4428 16816 4480
rect 18052 4632 18104 4684
rect 18328 4632 18380 4684
rect 18788 4675 18840 4684
rect 18788 4641 18806 4675
rect 18806 4641 18840 4675
rect 18788 4632 18840 4641
rect 2755 4326 2807 4378
rect 2819 4326 2871 4378
rect 2883 4326 2935 4378
rect 2947 4326 2999 4378
rect 3011 4326 3063 4378
rect 7470 4326 7522 4378
rect 7534 4326 7586 4378
rect 7598 4326 7650 4378
rect 7662 4326 7714 4378
rect 7726 4326 7778 4378
rect 12185 4326 12237 4378
rect 12249 4326 12301 4378
rect 12313 4326 12365 4378
rect 12377 4326 12429 4378
rect 12441 4326 12493 4378
rect 16900 4326 16952 4378
rect 16964 4326 17016 4378
rect 17028 4326 17080 4378
rect 17092 4326 17144 4378
rect 17156 4326 17208 4378
rect 1400 4224 1452 4276
rect 1124 4020 1176 4072
rect 1400 4063 1452 4072
rect 1400 4029 1409 4063
rect 1409 4029 1443 4063
rect 1443 4029 1452 4063
rect 1400 4020 1452 4029
rect 10232 4224 10284 4276
rect 10508 4224 10560 4276
rect 11520 4224 11572 4276
rect 1952 4156 2004 4208
rect 1676 4063 1728 4072
rect 1676 4029 1685 4063
rect 1685 4029 1719 4063
rect 1719 4029 1728 4063
rect 1676 4020 1728 4029
rect 4988 4088 5040 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 1308 3952 1360 4004
rect 5448 3952 5500 4004
rect 7288 3952 7340 4004
rect 1124 3884 1176 3936
rect 2044 3927 2096 3936
rect 2044 3893 2053 3927
rect 2053 3893 2087 3927
rect 2087 3893 2096 3927
rect 2044 3884 2096 3893
rect 8668 3884 8720 3936
rect 8852 3952 8904 4004
rect 10784 4020 10836 4072
rect 12532 4224 12584 4276
rect 14004 4224 14056 4276
rect 15936 4224 15988 4276
rect 17224 4224 17276 4276
rect 18328 4267 18380 4276
rect 18328 4233 18337 4267
rect 18337 4233 18371 4267
rect 18371 4233 18380 4267
rect 18328 4224 18380 4233
rect 18512 4224 18564 4276
rect 16764 4156 16816 4208
rect 13820 4020 13872 4072
rect 15384 4088 15436 4140
rect 15568 4088 15620 4140
rect 12808 3952 12860 4004
rect 11060 3884 11112 3936
rect 14372 3952 14424 4004
rect 15200 4020 15252 4072
rect 16120 4063 16172 4072
rect 16120 4029 16129 4063
rect 16129 4029 16163 4063
rect 16163 4029 16172 4063
rect 16120 4020 16172 4029
rect 16948 4063 17000 4072
rect 16948 4029 16957 4063
rect 16957 4029 16991 4063
rect 16991 4029 17000 4063
rect 16948 4020 17000 4029
rect 17316 4020 17368 4072
rect 18144 3952 18196 4004
rect 17868 3884 17920 3936
rect 5112 3782 5164 3834
rect 5176 3782 5228 3834
rect 5240 3782 5292 3834
rect 5304 3782 5356 3834
rect 5368 3782 5420 3834
rect 9827 3782 9879 3834
rect 9891 3782 9943 3834
rect 9955 3782 10007 3834
rect 10019 3782 10071 3834
rect 10083 3782 10135 3834
rect 14542 3782 14594 3834
rect 14606 3782 14658 3834
rect 14670 3782 14722 3834
rect 14734 3782 14786 3834
rect 14798 3782 14850 3834
rect 19257 3782 19309 3834
rect 19321 3782 19373 3834
rect 19385 3782 19437 3834
rect 19449 3782 19501 3834
rect 19513 3782 19565 3834
rect 1124 3723 1176 3732
rect 1124 3689 1133 3723
rect 1133 3689 1167 3723
rect 1167 3689 1176 3723
rect 1124 3680 1176 3689
rect 1676 3680 1728 3732
rect 4896 3680 4948 3732
rect 5632 3680 5684 3732
rect 6368 3680 6420 3732
rect 9128 3680 9180 3732
rect 10324 3680 10376 3732
rect 10692 3680 10744 3732
rect 1308 3587 1360 3596
rect 1308 3553 1317 3587
rect 1317 3553 1351 3587
rect 1351 3553 1360 3587
rect 1308 3544 1360 3553
rect 1584 3476 1636 3528
rect 1676 3476 1728 3528
rect 2596 3612 2648 3664
rect 2228 3587 2280 3596
rect 2228 3553 2262 3587
rect 2262 3553 2280 3587
rect 2228 3544 2280 3553
rect 14464 3680 14516 3732
rect 15108 3680 15160 3732
rect 15384 3680 15436 3732
rect 3700 3544 3752 3596
rect 5448 3544 5500 3596
rect 6092 3544 6144 3596
rect 6368 3544 6420 3596
rect 8760 3544 8812 3596
rect 12992 3587 13044 3596
rect 12992 3553 13001 3587
rect 13001 3553 13035 3587
rect 13035 3553 13044 3587
rect 12992 3544 13044 3553
rect 13084 3544 13136 3596
rect 14372 3544 14424 3596
rect 6552 3476 6604 3528
rect 9036 3476 9088 3528
rect 15108 3544 15160 3596
rect 15292 3476 15344 3528
rect 1860 3408 1912 3460
rect 4620 3408 4672 3460
rect 1768 3340 1820 3392
rect 2228 3340 2280 3392
rect 6460 3408 6512 3460
rect 15384 3408 15436 3460
rect 16304 3680 16356 3732
rect 16764 3723 16816 3732
rect 16764 3689 16773 3723
rect 16773 3689 16807 3723
rect 16807 3689 16816 3723
rect 16764 3680 16816 3689
rect 16948 3680 17000 3732
rect 17500 3680 17552 3732
rect 17868 3612 17920 3664
rect 15936 3476 15988 3528
rect 16120 3408 16172 3460
rect 18972 3587 19024 3596
rect 18972 3553 18981 3587
rect 18981 3553 19015 3587
rect 19015 3553 19024 3587
rect 18972 3544 19024 3553
rect 6368 3383 6420 3392
rect 6368 3349 6377 3383
rect 6377 3349 6411 3383
rect 6411 3349 6420 3383
rect 6368 3340 6420 3349
rect 15752 3383 15804 3392
rect 15752 3349 15761 3383
rect 15761 3349 15795 3383
rect 15795 3349 15804 3383
rect 15752 3340 15804 3349
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 2755 3238 2807 3290
rect 2819 3238 2871 3290
rect 2883 3238 2935 3290
rect 2947 3238 2999 3290
rect 3011 3238 3063 3290
rect 7470 3238 7522 3290
rect 7534 3238 7586 3290
rect 7598 3238 7650 3290
rect 7662 3238 7714 3290
rect 7726 3238 7778 3290
rect 12185 3238 12237 3290
rect 12249 3238 12301 3290
rect 12313 3238 12365 3290
rect 12377 3238 12429 3290
rect 12441 3238 12493 3290
rect 16900 3238 16952 3290
rect 16964 3238 17016 3290
rect 17028 3238 17080 3290
rect 17092 3238 17144 3290
rect 17156 3238 17208 3290
rect 1308 2975 1360 2984
rect 1308 2941 1317 2975
rect 1317 2941 1351 2975
rect 1351 2941 1360 2975
rect 1308 2932 1360 2941
rect 1860 3136 1912 3188
rect 4804 3136 4856 3188
rect 7288 3179 7340 3188
rect 7288 3145 7297 3179
rect 7297 3145 7331 3179
rect 7331 3145 7340 3179
rect 7288 3136 7340 3145
rect 8392 3136 8444 3188
rect 8760 3179 8812 3188
rect 8760 3145 8769 3179
rect 8769 3145 8803 3179
rect 8803 3145 8812 3179
rect 8760 3136 8812 3145
rect 11336 3136 11388 3188
rect 12808 3136 12860 3188
rect 13084 3136 13136 3188
rect 15108 3179 15160 3188
rect 15108 3145 15117 3179
rect 15117 3145 15151 3179
rect 15151 3145 15160 3179
rect 15108 3136 15160 3145
rect 15292 3136 15344 3188
rect 15752 3179 15804 3188
rect 15752 3145 15761 3179
rect 15761 3145 15795 3179
rect 15795 3145 15804 3179
rect 15752 3136 15804 3145
rect 16120 3179 16172 3188
rect 16120 3145 16129 3179
rect 16129 3145 16163 3179
rect 16163 3145 16172 3179
rect 16120 3136 16172 3145
rect 17224 3136 17276 3188
rect 2228 2932 2280 2984
rect 5540 2932 5592 2984
rect 6368 2932 6420 2984
rect 7656 2975 7708 2984
rect 7656 2941 7665 2975
rect 7665 2941 7699 2975
rect 7699 2941 7708 2975
rect 7656 2932 7708 2941
rect 12532 3000 12584 3052
rect 15568 3068 15620 3120
rect 15844 3068 15896 3120
rect 12808 2975 12860 2984
rect 12808 2941 12817 2975
rect 12817 2941 12851 2975
rect 12851 2941 12860 2975
rect 12808 2932 12860 2941
rect 16304 3000 16356 3052
rect 1952 2907 2004 2916
rect 1952 2873 1986 2907
rect 1986 2873 2004 2907
rect 1952 2864 2004 2873
rect 2412 2864 2464 2916
rect 13268 2864 13320 2916
rect 16488 2975 16540 2984
rect 16488 2941 16497 2975
rect 16497 2941 16531 2975
rect 16531 2941 16540 2975
rect 16488 2932 16540 2941
rect 16028 2864 16080 2916
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 18972 3000 19024 3052
rect 16764 2932 16816 2984
rect 1216 2839 1268 2848
rect 1216 2805 1225 2839
rect 1225 2805 1259 2839
rect 1259 2805 1268 2839
rect 1216 2796 1268 2805
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 1676 2796 1728 2848
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 6920 2839 6972 2848
rect 6920 2805 6929 2839
rect 6929 2805 6963 2839
rect 6963 2805 6972 2839
rect 6920 2796 6972 2805
rect 15292 2796 15344 2848
rect 15936 2796 15988 2848
rect 16396 2839 16448 2848
rect 16396 2805 16405 2839
rect 16405 2805 16439 2839
rect 16439 2805 16448 2839
rect 16396 2796 16448 2805
rect 16580 2796 16632 2848
rect 17776 2864 17828 2916
rect 5112 2694 5164 2746
rect 5176 2694 5228 2746
rect 5240 2694 5292 2746
rect 5304 2694 5356 2746
rect 5368 2694 5420 2746
rect 9827 2694 9879 2746
rect 9891 2694 9943 2746
rect 9955 2694 10007 2746
rect 10019 2694 10071 2746
rect 10083 2694 10135 2746
rect 14542 2694 14594 2746
rect 14606 2694 14658 2746
rect 14670 2694 14722 2746
rect 14734 2694 14786 2746
rect 14798 2694 14850 2746
rect 19257 2694 19309 2746
rect 19321 2694 19373 2746
rect 19385 2694 19437 2746
rect 19449 2694 19501 2746
rect 19513 2694 19565 2746
rect 1492 2592 1544 2644
rect 1952 2635 2004 2644
rect 1952 2601 1961 2635
rect 1961 2601 1995 2635
rect 1995 2601 2004 2635
rect 1952 2592 2004 2601
rect 1768 2524 1820 2576
rect 1860 2524 1912 2576
rect 1216 2499 1268 2508
rect 1216 2465 1225 2499
rect 1225 2465 1259 2499
rect 1259 2465 1268 2499
rect 1216 2456 1268 2465
rect 1492 2499 1544 2508
rect 1492 2465 1501 2499
rect 1501 2465 1535 2499
rect 1535 2465 1544 2499
rect 1492 2456 1544 2465
rect 1308 2388 1360 2440
rect 2228 2456 2280 2508
rect 2504 2456 2556 2508
rect 3700 2592 3752 2644
rect 4160 2592 4212 2644
rect 4620 2592 4672 2644
rect 5632 2592 5684 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 7380 2592 7432 2644
rect 3240 2524 3292 2576
rect 1400 2295 1452 2304
rect 1400 2261 1409 2295
rect 1409 2261 1443 2295
rect 1443 2261 1452 2295
rect 1400 2252 1452 2261
rect 2596 2252 2648 2304
rect 3608 2499 3660 2508
rect 3608 2465 3617 2499
rect 3617 2465 3651 2499
rect 3651 2465 3660 2499
rect 3608 2456 3660 2465
rect 5540 2524 5592 2576
rect 4988 2499 5040 2508
rect 4988 2465 4997 2499
rect 4997 2465 5031 2499
rect 5031 2465 5040 2499
rect 4988 2456 5040 2465
rect 5816 2524 5868 2576
rect 8392 2524 8444 2576
rect 4988 2320 5040 2372
rect 6368 2456 6420 2508
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 8208 2388 8260 2440
rect 8668 2456 8720 2508
rect 9312 2524 9364 2576
rect 3516 2295 3568 2304
rect 3516 2261 3525 2295
rect 3525 2261 3559 2295
rect 3559 2261 3568 2295
rect 3516 2252 3568 2261
rect 3700 2252 3752 2304
rect 5540 2295 5592 2304
rect 5540 2261 5549 2295
rect 5549 2261 5583 2295
rect 5583 2261 5592 2295
rect 5540 2252 5592 2261
rect 6092 2295 6144 2304
rect 6092 2261 6101 2295
rect 6101 2261 6135 2295
rect 6135 2261 6144 2295
rect 6092 2252 6144 2261
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 8208 2252 8260 2261
rect 8484 2295 8536 2304
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 9680 2499 9732 2508
rect 9680 2465 9689 2499
rect 9689 2465 9723 2499
rect 9723 2465 9732 2499
rect 9680 2456 9732 2465
rect 10600 2635 10652 2644
rect 10600 2601 10609 2635
rect 10609 2601 10643 2635
rect 10643 2601 10652 2635
rect 10600 2592 10652 2601
rect 13452 2524 13504 2576
rect 15292 2592 15344 2644
rect 15660 2592 15712 2644
rect 16580 2592 16632 2644
rect 17316 2592 17368 2644
rect 17868 2592 17920 2644
rect 10232 2388 10284 2440
rect 10876 2456 10928 2508
rect 8484 2252 8536 2261
rect 8944 2252 8996 2304
rect 9128 2295 9180 2304
rect 9128 2261 9137 2295
rect 9137 2261 9171 2295
rect 9171 2261 9180 2295
rect 9128 2252 9180 2261
rect 9588 2252 9640 2304
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 10140 2252 10192 2304
rect 11060 2499 11112 2508
rect 11060 2465 11069 2499
rect 11069 2465 11103 2499
rect 11103 2465 11112 2499
rect 11060 2456 11112 2465
rect 12532 2456 12584 2508
rect 12716 2499 12768 2508
rect 12716 2465 12750 2499
rect 12750 2465 12768 2499
rect 12716 2456 12768 2465
rect 14004 2456 14056 2508
rect 15660 2499 15712 2508
rect 15660 2465 15669 2499
rect 15669 2465 15703 2499
rect 15703 2465 15712 2499
rect 15660 2456 15712 2465
rect 16120 2456 16172 2508
rect 17776 2524 17828 2576
rect 16396 2320 16448 2372
rect 11336 2295 11388 2304
rect 11336 2261 11345 2295
rect 11345 2261 11379 2295
rect 11379 2261 11388 2295
rect 11336 2252 11388 2261
rect 11980 2252 12032 2304
rect 14280 2252 14332 2304
rect 15752 2295 15804 2304
rect 15752 2261 15761 2295
rect 15761 2261 15795 2295
rect 15795 2261 15804 2295
rect 15752 2252 15804 2261
rect 15936 2252 15988 2304
rect 19064 2295 19116 2304
rect 19064 2261 19073 2295
rect 19073 2261 19107 2295
rect 19107 2261 19116 2295
rect 19064 2252 19116 2261
rect 2755 2150 2807 2202
rect 2819 2150 2871 2202
rect 2883 2150 2935 2202
rect 2947 2150 2999 2202
rect 3011 2150 3063 2202
rect 7470 2150 7522 2202
rect 7534 2150 7586 2202
rect 7598 2150 7650 2202
rect 7662 2150 7714 2202
rect 7726 2150 7778 2202
rect 12185 2150 12237 2202
rect 12249 2150 12301 2202
rect 12313 2150 12365 2202
rect 12377 2150 12429 2202
rect 12441 2150 12493 2202
rect 16900 2150 16952 2202
rect 16964 2150 17016 2202
rect 17028 2150 17080 2202
rect 17092 2150 17144 2202
rect 17156 2150 17208 2202
rect 1216 2048 1268 2100
rect 1400 2048 1452 2100
rect 2504 2048 2556 2100
rect 2780 2048 2832 2100
rect 3516 2048 3568 2100
rect 1216 1887 1268 1896
rect 1216 1853 1225 1887
rect 1225 1853 1259 1887
rect 1259 1853 1268 1887
rect 1216 1844 1268 1853
rect 4160 2048 4212 2100
rect 7012 2091 7064 2100
rect 7012 2057 7021 2091
rect 7021 2057 7055 2091
rect 7055 2057 7064 2091
rect 7012 2048 7064 2057
rect 7472 2048 7524 2100
rect 8208 2048 8260 2100
rect 8576 2091 8628 2100
rect 8576 2057 8585 2091
rect 8585 2057 8619 2091
rect 8619 2057 8628 2091
rect 8576 2048 8628 2057
rect 2228 1912 2280 1964
rect 2412 1912 2464 1964
rect 3240 1912 3292 1964
rect 2596 1887 2648 1896
rect 2596 1853 2605 1887
rect 2605 1853 2639 1887
rect 2639 1853 2648 1887
rect 2596 1844 2648 1853
rect 2780 1844 2832 1896
rect 3700 1912 3752 1964
rect 3516 1844 3568 1896
rect 6920 1912 6972 1964
rect 3884 1887 3936 1896
rect 3884 1853 3893 1887
rect 3893 1853 3927 1887
rect 3927 1853 3936 1887
rect 3884 1844 3936 1853
rect 5632 1887 5684 1896
rect 5632 1853 5666 1887
rect 5666 1853 5684 1887
rect 5632 1844 5684 1853
rect 5908 1844 5960 1896
rect 7196 1887 7248 1896
rect 7196 1853 7205 1887
rect 7205 1853 7239 1887
rect 7239 1853 7248 1887
rect 7196 1844 7248 1853
rect 7564 1912 7616 1964
rect 7840 1912 7892 1964
rect 8484 1980 8536 2032
rect 10232 2048 10284 2100
rect 11336 2048 11388 2100
rect 12072 2048 12124 2100
rect 12716 2048 12768 2100
rect 13268 2091 13320 2100
rect 13268 2057 13277 2091
rect 13277 2057 13311 2091
rect 13311 2057 13320 2091
rect 13268 2048 13320 2057
rect 10140 1980 10192 2032
rect 11980 1980 12032 2032
rect 9036 1955 9088 1964
rect 9036 1921 9045 1955
rect 9045 1921 9079 1955
rect 9079 1921 9088 1955
rect 9036 1912 9088 1921
rect 10784 1912 10836 1964
rect 8392 1844 8444 1896
rect 4436 1776 4488 1828
rect 1492 1708 1544 1760
rect 2688 1708 2740 1760
rect 4896 1708 4948 1760
rect 7380 1708 7432 1760
rect 9680 1844 9732 1896
rect 14004 1980 14056 2032
rect 8944 1776 8996 1828
rect 10324 1776 10376 1828
rect 11428 1776 11480 1828
rect 13084 1844 13136 1896
rect 14188 1844 14240 1896
rect 15660 2048 15712 2100
rect 16672 2091 16724 2100
rect 16672 2057 16681 2091
rect 16681 2057 16715 2091
rect 16715 2057 16724 2091
rect 16672 2048 16724 2057
rect 17960 2048 18012 2100
rect 18512 1912 18564 1964
rect 15016 1863 15025 1896
rect 15025 1863 15059 1896
rect 15059 1863 15068 1896
rect 15016 1844 15068 1863
rect 15292 1887 15344 1896
rect 15292 1853 15301 1887
rect 15301 1853 15335 1887
rect 15335 1853 15344 1887
rect 15292 1844 15344 1853
rect 16488 1844 16540 1896
rect 19064 1887 19116 1896
rect 19064 1853 19073 1887
rect 19073 1853 19107 1887
rect 19107 1853 19116 1887
rect 19064 1844 19116 1853
rect 10416 1708 10468 1760
rect 10600 1708 10652 1760
rect 12164 1708 12216 1760
rect 13176 1708 13228 1760
rect 13912 1751 13964 1760
rect 13912 1717 13921 1751
rect 13921 1717 13955 1751
rect 13955 1717 13964 1751
rect 13912 1708 13964 1717
rect 15200 1776 15252 1828
rect 15752 1776 15804 1828
rect 16304 1776 16356 1828
rect 16580 1776 16632 1828
rect 15660 1708 15712 1760
rect 16212 1708 16264 1760
rect 5112 1606 5164 1658
rect 5176 1606 5228 1658
rect 5240 1606 5292 1658
rect 5304 1606 5356 1658
rect 5368 1606 5420 1658
rect 9827 1606 9879 1658
rect 9891 1606 9943 1658
rect 9955 1606 10007 1658
rect 10019 1606 10071 1658
rect 10083 1606 10135 1658
rect 14542 1606 14594 1658
rect 14606 1606 14658 1658
rect 14670 1606 14722 1658
rect 14734 1606 14786 1658
rect 14798 1606 14850 1658
rect 19257 1606 19309 1658
rect 19321 1606 19373 1658
rect 19385 1606 19437 1658
rect 19449 1606 19501 1658
rect 19513 1606 19565 1658
rect 1400 1504 1452 1556
rect 1492 1547 1544 1556
rect 1492 1513 1501 1547
rect 1501 1513 1535 1547
rect 1535 1513 1544 1547
rect 1492 1504 1544 1513
rect 4436 1504 4488 1556
rect 4804 1547 4856 1556
rect 4804 1513 4813 1547
rect 4813 1513 4847 1547
rect 4847 1513 4856 1547
rect 4804 1504 4856 1513
rect 4988 1547 5040 1556
rect 4988 1513 4997 1547
rect 4997 1513 5031 1547
rect 5031 1513 5040 1547
rect 4988 1504 5040 1513
rect 5540 1504 5592 1556
rect 2044 1436 2096 1488
rect 3240 1436 3292 1488
rect 3884 1436 3936 1488
rect 1676 1343 1728 1352
rect 1676 1309 1685 1343
rect 1685 1309 1719 1343
rect 1719 1309 1728 1343
rect 1676 1300 1728 1309
rect 5172 1411 5224 1420
rect 5172 1377 5181 1411
rect 5181 1377 5215 1411
rect 5215 1377 5224 1411
rect 5172 1368 5224 1377
rect 5356 1368 5408 1420
rect 5816 1504 5868 1556
rect 6920 1436 6972 1488
rect 6368 1411 6420 1420
rect 6368 1377 6377 1411
rect 6377 1377 6411 1411
rect 6411 1377 6420 1411
rect 6368 1368 6420 1377
rect 7012 1368 7064 1420
rect 8300 1547 8352 1556
rect 8300 1513 8309 1547
rect 8309 1513 8343 1547
rect 8343 1513 8352 1547
rect 8300 1504 8352 1513
rect 8484 1504 8536 1556
rect 8760 1504 8812 1556
rect 9128 1504 9180 1556
rect 9588 1504 9640 1556
rect 10416 1547 10468 1556
rect 10416 1513 10425 1547
rect 10425 1513 10459 1547
rect 10459 1513 10468 1547
rect 10416 1504 10468 1513
rect 7196 1411 7248 1420
rect 7196 1377 7230 1411
rect 7230 1377 7248 1411
rect 7196 1368 7248 1377
rect 10324 1368 10376 1420
rect 2780 1232 2832 1284
rect 3332 1232 3384 1284
rect 6552 1300 6604 1352
rect 8392 1343 8444 1352
rect 6092 1232 6144 1284
rect 8392 1309 8401 1343
rect 8401 1309 8435 1343
rect 8435 1309 8444 1343
rect 8392 1300 8444 1309
rect 10600 1411 10652 1420
rect 10600 1377 10609 1411
rect 10609 1377 10643 1411
rect 10643 1377 10652 1411
rect 10600 1368 10652 1377
rect 11060 1547 11112 1556
rect 11060 1513 11069 1547
rect 11069 1513 11103 1547
rect 11103 1513 11112 1547
rect 11060 1504 11112 1513
rect 11336 1504 11388 1556
rect 11428 1504 11480 1556
rect 11244 1411 11296 1420
rect 11244 1377 11253 1411
rect 11253 1377 11287 1411
rect 11287 1377 11296 1411
rect 11244 1368 11296 1377
rect 11428 1368 11480 1420
rect 12164 1411 12216 1420
rect 12164 1377 12173 1411
rect 12173 1377 12207 1411
rect 12207 1377 12216 1411
rect 12164 1368 12216 1377
rect 12716 1504 12768 1556
rect 14188 1504 14240 1556
rect 14924 1504 14976 1556
rect 15200 1504 15252 1556
rect 13912 1436 13964 1488
rect 13176 1411 13228 1420
rect 13176 1377 13185 1411
rect 13185 1377 13219 1411
rect 13219 1377 13228 1411
rect 13176 1368 13228 1377
rect 13452 1411 13504 1420
rect 13452 1377 13461 1411
rect 13461 1377 13495 1411
rect 13495 1377 13504 1411
rect 13452 1368 13504 1377
rect 13544 1368 13596 1420
rect 15016 1436 15068 1488
rect 16120 1504 16172 1556
rect 16212 1547 16264 1556
rect 16212 1513 16221 1547
rect 16221 1513 16255 1547
rect 16255 1513 16264 1547
rect 16212 1504 16264 1513
rect 18236 1504 18288 1556
rect 13176 1232 13228 1284
rect 11244 1164 11296 1216
rect 14464 1164 14516 1216
rect 15660 1411 15712 1420
rect 15660 1377 15669 1411
rect 15669 1377 15703 1411
rect 15703 1377 15712 1411
rect 15660 1368 15712 1377
rect 16396 1368 16448 1420
rect 16488 1411 16540 1420
rect 16488 1377 16497 1411
rect 16497 1377 16531 1411
rect 16531 1377 16540 1411
rect 16488 1368 16540 1377
rect 16580 1368 16632 1420
rect 16120 1300 16172 1352
rect 2755 1062 2807 1114
rect 2819 1062 2871 1114
rect 2883 1062 2935 1114
rect 2947 1062 2999 1114
rect 3011 1062 3063 1114
rect 7470 1062 7522 1114
rect 7534 1062 7586 1114
rect 7598 1062 7650 1114
rect 7662 1062 7714 1114
rect 7726 1062 7778 1114
rect 12185 1062 12237 1114
rect 12249 1062 12301 1114
rect 12313 1062 12365 1114
rect 12377 1062 12429 1114
rect 12441 1062 12493 1114
rect 16900 1062 16952 1114
rect 16964 1062 17016 1114
rect 17028 1062 17080 1114
rect 17092 1062 17144 1114
rect 17156 1062 17208 1114
rect 2228 1003 2280 1012
rect 2228 969 2237 1003
rect 2237 969 2271 1003
rect 2271 969 2280 1003
rect 2228 960 2280 969
rect 4896 960 4948 1012
rect 7196 1003 7248 1012
rect 7196 969 7205 1003
rect 7205 969 7239 1003
rect 7239 969 7248 1003
rect 7196 960 7248 969
rect 11152 960 11204 1012
rect 11888 960 11940 1012
rect 13544 960 13596 1012
rect 1952 892 2004 944
rect 11796 892 11848 944
rect 12900 935 12952 944
rect 12900 901 12909 935
rect 12909 901 12943 935
rect 12943 901 12952 935
rect 12900 892 12952 901
rect 2044 824 2096 876
rect 13912 1003 13964 1012
rect 13912 969 13921 1003
rect 13921 969 13955 1003
rect 13955 969 13964 1003
rect 13912 960 13964 969
rect 14188 1003 14240 1012
rect 14188 969 14197 1003
rect 14197 969 14231 1003
rect 14231 969 14240 1003
rect 14188 960 14240 969
rect 14464 1003 14516 1012
rect 14464 969 14473 1003
rect 14473 969 14507 1003
rect 14507 969 14516 1003
rect 14464 960 14516 969
rect 15936 960 15988 1012
rect 16304 960 16356 1012
rect 848 799 900 808
rect 848 765 857 799
rect 857 765 891 799
rect 891 765 900 799
rect 848 756 900 765
rect 1308 756 1360 808
rect 3608 756 3660 808
rect 6920 756 6972 808
rect 10416 799 10468 808
rect 10416 765 10425 799
rect 10425 765 10459 799
rect 10459 765 10468 799
rect 10416 756 10468 765
rect 13176 756 13228 808
rect 11796 731 11848 740
rect 11796 697 11805 731
rect 11805 697 11839 731
rect 11839 697 11848 731
rect 11796 688 11848 697
rect 12256 688 12308 740
rect 13084 731 13136 740
rect 13084 697 13093 731
rect 13093 697 13127 731
rect 13127 697 13136 731
rect 13084 688 13136 697
rect 16120 799 16172 808
rect 16120 765 16129 799
rect 16129 765 16163 799
rect 16163 765 16172 799
rect 16120 756 16172 765
rect 16304 756 16356 808
rect 16580 799 16632 808
rect 16580 765 16589 799
rect 16589 765 16623 799
rect 16623 765 16632 799
rect 16580 756 16632 765
rect 18512 799 18564 808
rect 18512 765 18521 799
rect 18521 765 18555 799
rect 18555 765 18564 799
rect 18512 756 18564 765
rect 19064 799 19116 808
rect 19064 765 19073 799
rect 19073 765 19107 799
rect 19107 765 19116 799
rect 19064 756 19116 765
rect 5112 518 5164 570
rect 5176 518 5228 570
rect 5240 518 5292 570
rect 5304 518 5356 570
rect 5368 518 5420 570
rect 9827 518 9879 570
rect 9891 518 9943 570
rect 9955 518 10007 570
rect 10019 518 10071 570
rect 10083 518 10135 570
rect 14542 518 14594 570
rect 14606 518 14658 570
rect 14670 518 14722 570
rect 14734 518 14786 570
rect 14798 518 14850 570
rect 19257 518 19309 570
rect 19321 518 19373 570
rect 19385 518 19437 570
rect 19449 518 19501 570
rect 19513 518 19565 570
<< metal2 >>
rect 1122 19816 1178 19825
rect 1122 19751 1178 19760
rect 754 19136 810 19145
rect 754 19071 810 19080
rect 768 18834 796 19071
rect 756 18828 808 18834
rect 756 18770 808 18776
rect 1136 18766 1164 19751
rect 11610 19600 11666 20000
rect 5112 19068 5420 19077
rect 5112 19066 5118 19068
rect 5174 19066 5198 19068
rect 5254 19066 5278 19068
rect 5334 19066 5358 19068
rect 5414 19066 5420 19068
rect 5174 19014 5176 19066
rect 5356 19014 5358 19066
rect 5112 19012 5118 19014
rect 5174 19012 5198 19014
rect 5254 19012 5278 19014
rect 5334 19012 5358 19014
rect 5414 19012 5420 19014
rect 5112 19003 5420 19012
rect 9827 19068 10135 19077
rect 9827 19066 9833 19068
rect 9889 19066 9913 19068
rect 9969 19066 9993 19068
rect 10049 19066 10073 19068
rect 10129 19066 10135 19068
rect 9889 19014 9891 19066
rect 10071 19014 10073 19066
rect 9827 19012 9833 19014
rect 9889 19012 9913 19014
rect 9969 19012 9993 19014
rect 10049 19012 10073 19014
rect 10129 19012 10135 19014
rect 9827 19003 10135 19012
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 1124 18760 1176 18766
rect 1124 18702 1176 18708
rect 848 18624 900 18630
rect 848 18566 900 18572
rect 860 18465 888 18566
rect 2755 18524 3063 18533
rect 2755 18522 2761 18524
rect 2817 18522 2841 18524
rect 2897 18522 2921 18524
rect 2977 18522 3001 18524
rect 3057 18522 3063 18524
rect 2817 18470 2819 18522
rect 2999 18470 3001 18522
rect 2755 18468 2761 18470
rect 2817 18468 2841 18470
rect 2897 18468 2921 18470
rect 2977 18468 3001 18470
rect 3057 18468 3063 18470
rect 846 18456 902 18465
rect 2755 18459 3063 18468
rect 7470 18524 7778 18533
rect 7470 18522 7476 18524
rect 7532 18522 7556 18524
rect 7612 18522 7636 18524
rect 7692 18522 7716 18524
rect 7772 18522 7778 18524
rect 7532 18470 7534 18522
rect 7714 18470 7716 18522
rect 7470 18468 7476 18470
rect 7532 18468 7556 18470
rect 7612 18468 7636 18470
rect 7692 18468 7716 18470
rect 7772 18468 7778 18470
rect 7470 18459 7778 18468
rect 10428 18426 10456 18838
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11440 18426 11468 18566
rect 846 18391 902 18400
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 10520 18306 10548 18362
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 10336 18278 10548 18306
rect 848 18216 900 18222
rect 848 18158 900 18164
rect 860 17785 888 18158
rect 846 17776 902 17785
rect 846 17711 902 17720
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1504 17134 1532 17614
rect 1596 17202 1624 17614
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1872 17134 1900 17478
rect 2240 17338 2268 17478
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 848 17128 900 17134
rect 846 17096 848 17105
rect 1492 17128 1544 17134
rect 900 17096 902 17105
rect 1492 17070 1544 17076
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 846 17031 902 17040
rect 1872 16794 1900 17070
rect 2240 16794 2268 17274
rect 2332 16998 2360 17682
rect 2424 17678 2452 18226
rect 10336 18222 10364 18278
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 8392 18216 8444 18222
rect 10324 18216 10376 18222
rect 8392 18158 8444 18164
rect 10152 18176 10324 18204
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2608 17814 2636 18022
rect 2596 17808 2648 17814
rect 2596 17750 2648 17756
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 2700 17490 2728 18158
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 4160 18148 4212 18154
rect 4160 18090 4212 18096
rect 2608 17462 2728 17490
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2332 16794 2360 16934
rect 2608 16810 2636 17462
rect 2755 17436 3063 17445
rect 2755 17434 2761 17436
rect 2817 17434 2841 17436
rect 2897 17434 2921 17436
rect 2977 17434 3001 17436
rect 3057 17434 3063 17436
rect 2817 17382 2819 17434
rect 2999 17382 3001 17434
rect 2755 17380 2761 17382
rect 2817 17380 2841 17382
rect 2897 17380 2921 17382
rect 2977 17380 3001 17382
rect 3057 17380 3063 17382
rect 2755 17371 3063 17380
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 2608 16794 2820 16810
rect 3160 16794 3188 17002
rect 3804 16998 3832 18090
rect 4172 17746 4200 18090
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 5112 17980 5420 17989
rect 5112 17978 5118 17980
rect 5174 17978 5198 17980
rect 5254 17978 5278 17980
rect 5334 17978 5358 17980
rect 5414 17978 5420 17980
rect 5174 17926 5176 17978
rect 5356 17926 5358 17978
rect 5112 17924 5118 17926
rect 5174 17924 5198 17926
rect 5254 17924 5278 17926
rect 5334 17924 5358 17926
rect 5414 17924 5420 17926
rect 5112 17915 5420 17924
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 3884 17060 3936 17066
rect 3884 17002 3936 17008
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3712 16794 3740 16934
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2608 16788 2832 16794
rect 2608 16782 2780 16788
rect 1412 16046 1440 16730
rect 2608 16726 2636 16782
rect 2780 16730 2832 16736
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 16182 1624 16594
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 2412 16448 2464 16454
rect 2464 16408 2544 16436
rect 2412 16390 2464 16396
rect 1584 16176 1636 16182
rect 1584 16118 1636 16124
rect 1872 16046 1900 16390
rect 2516 16114 2544 16408
rect 2755 16348 3063 16357
rect 2755 16346 2761 16348
rect 2817 16346 2841 16348
rect 2897 16346 2921 16348
rect 2977 16346 3001 16348
rect 3057 16346 3063 16348
rect 2817 16294 2819 16346
rect 2999 16294 3001 16346
rect 2755 16292 2761 16294
rect 2817 16292 2841 16294
rect 2897 16292 2921 16294
rect 2977 16292 3001 16294
rect 3057 16292 3063 16294
rect 2755 16283 3063 16292
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 2228 15904 2280 15910
rect 2228 15846 2280 15852
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 1780 15706 1808 15846
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 2240 15638 2268 15846
rect 2228 15632 2280 15638
rect 2228 15574 2280 15580
rect 1492 15564 1544 15570
rect 1492 15506 1544 15512
rect 1504 14958 1532 15506
rect 2044 15428 2096 15434
rect 2044 15370 2096 15376
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1688 14634 1716 15302
rect 1596 14618 1716 14634
rect 1584 14612 1716 14618
rect 1636 14606 1716 14612
rect 1584 14554 1636 14560
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1412 14074 1440 14214
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1596 13870 1624 14554
rect 1688 14482 1716 14606
rect 2056 14550 2084 15370
rect 2240 15366 2268 15574
rect 2332 15502 2360 15846
rect 2424 15570 2452 15846
rect 2516 15638 2544 16050
rect 3252 16046 3280 16526
rect 3804 16454 3832 16934
rect 3896 16794 3924 17002
rect 4080 16998 4108 17478
rect 4172 17202 4200 17682
rect 4356 17338 4384 17818
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4448 17338 4476 17682
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 4080 16658 4108 16934
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3422 16144 3478 16153
rect 3422 16079 3478 16088
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 2504 15632 2556 15638
rect 2504 15574 2556 15580
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2044 14544 2096 14550
rect 2044 14486 2096 14492
rect 2240 14482 2268 15302
rect 2332 14958 2360 15438
rect 2755 15260 3063 15269
rect 2755 15258 2761 15260
rect 2817 15258 2841 15260
rect 2897 15258 2921 15260
rect 2977 15258 3001 15260
rect 3057 15258 3063 15260
rect 2817 15206 2819 15258
rect 2999 15206 3001 15258
rect 2755 15204 2761 15206
rect 2817 15204 2841 15206
rect 2897 15204 2921 15206
rect 2977 15204 3001 15206
rect 3057 15204 3063 15206
rect 2755 15195 3063 15204
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1964 14074 1992 14214
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1780 13870 1808 14010
rect 1964 13954 1992 14010
rect 1964 13938 2176 13954
rect 1964 13932 2188 13938
rect 1964 13926 2136 13932
rect 2136 13874 2188 13880
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1596 13462 1624 13806
rect 1584 13456 1636 13462
rect 1584 13398 1636 13404
rect 1216 13388 1268 13394
rect 1216 13330 1268 13336
rect 1228 12102 1256 13330
rect 1308 12368 1360 12374
rect 1308 12310 1360 12316
rect 1216 12096 1268 12102
rect 1216 12038 1268 12044
rect 1228 11558 1256 12038
rect 1216 11552 1268 11558
rect 1216 11494 1268 11500
rect 1228 11150 1256 11494
rect 1320 11354 1348 12310
rect 1780 11694 1808 13806
rect 2424 12374 2452 15030
rect 3344 14958 3372 15506
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 2872 14884 2924 14890
rect 2872 14826 2924 14832
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 14618 2636 14758
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2608 14074 2636 14554
rect 2884 14550 2912 14826
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2755 14172 3063 14181
rect 2755 14170 2761 14172
rect 2817 14170 2841 14172
rect 2897 14170 2921 14172
rect 2977 14170 3001 14172
rect 3057 14170 3063 14172
rect 2817 14118 2819 14170
rect 2999 14118 3001 14170
rect 2755 14116 2761 14118
rect 2817 14116 2841 14118
rect 2897 14116 2921 14118
rect 2977 14116 3001 14118
rect 3057 14116 3063 14118
rect 2755 14107 3063 14116
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 3344 13938 3372 14894
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 2516 13394 2544 13670
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2608 13190 2636 13670
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2608 12918 2636 13126
rect 2755 13084 3063 13093
rect 2755 13082 2761 13084
rect 2817 13082 2841 13084
rect 2897 13082 2921 13084
rect 2977 13082 3001 13084
rect 3057 13082 3063 13084
rect 2817 13030 2819 13082
rect 2999 13030 3001 13082
rect 2755 13028 2761 13030
rect 2817 13028 2841 13030
rect 2897 13028 2921 13030
rect 2977 13028 3001 13030
rect 3057 13028 3063 13030
rect 2755 13019 3063 13028
rect 2596 12912 2648 12918
rect 2596 12854 2648 12860
rect 3160 12714 3188 13670
rect 3252 13462 3280 13738
rect 3344 13462 3372 13874
rect 3240 13456 3292 13462
rect 3240 13398 3292 13404
rect 3332 13456 3384 13462
rect 3332 13398 3384 13404
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3252 12850 3280 13262
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2412 12368 2464 12374
rect 2412 12310 2464 12316
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1400 11620 1452 11626
rect 1400 11562 1452 11568
rect 1308 11348 1360 11354
rect 1308 11290 1360 11296
rect 1216 11144 1268 11150
rect 1216 11086 1268 11092
rect 1228 10130 1256 11086
rect 1216 10124 1268 10130
rect 1216 10066 1268 10072
rect 1032 9512 1084 9518
rect 1032 9454 1084 9460
rect 1044 9042 1072 9454
rect 1124 9444 1176 9450
rect 1124 9386 1176 9392
rect 1136 9042 1164 9386
rect 1032 9036 1084 9042
rect 1032 8978 1084 8984
rect 1124 9036 1176 9042
rect 1124 8978 1176 8984
rect 1032 8424 1084 8430
rect 1032 8366 1084 8372
rect 940 7812 992 7818
rect 940 7754 992 7760
rect 952 6730 980 7754
rect 1044 7546 1072 8366
rect 1136 8362 1164 8978
rect 1124 8356 1176 8362
rect 1124 8298 1176 8304
rect 1032 7540 1084 7546
rect 1032 7482 1084 7488
rect 940 6724 992 6730
rect 940 6666 992 6672
rect 952 6254 980 6666
rect 1044 6644 1072 7482
rect 1136 6866 1164 8298
rect 1216 8288 1268 8294
rect 1216 8230 1268 8236
rect 1228 8090 1256 8230
rect 1216 8084 1268 8090
rect 1216 8026 1268 8032
rect 1228 7528 1256 8026
rect 1320 7818 1348 11290
rect 1412 11286 1440 11562
rect 1400 11280 1452 11286
rect 1400 11222 1452 11228
rect 1412 8634 1440 11222
rect 1780 11218 1808 11630
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 2424 10606 2452 12038
rect 2516 11830 2544 12582
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2608 11898 2636 12242
rect 2755 11996 3063 12005
rect 2755 11994 2761 11996
rect 2817 11994 2841 11996
rect 2897 11994 2921 11996
rect 2977 11994 3001 11996
rect 3057 11994 3063 11996
rect 2817 11942 2819 11994
rect 2999 11942 3001 11994
rect 2755 11940 2761 11942
rect 2817 11940 2841 11942
rect 2897 11940 2921 11942
rect 2977 11940 3001 11942
rect 3057 11940 3063 11942
rect 2755 11931 3063 11940
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 2755 10908 3063 10917
rect 2755 10906 2761 10908
rect 2817 10906 2841 10908
rect 2897 10906 2921 10908
rect 2977 10906 3001 10908
rect 3057 10906 3063 10908
rect 2817 10854 2819 10906
rect 2999 10854 3001 10906
rect 2755 10852 2761 10854
rect 2817 10852 2841 10854
rect 2897 10852 2921 10854
rect 2977 10852 3001 10854
rect 3057 10852 3063 10854
rect 2755 10843 3063 10852
rect 3160 10606 3188 10950
rect 3252 10674 3280 11222
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3344 10606 3372 11494
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 1584 10192 1636 10198
rect 1584 10134 1636 10140
rect 1596 9178 1624 10134
rect 2516 9722 2544 10542
rect 3068 10452 3096 10542
rect 3068 10424 3188 10452
rect 2755 9820 3063 9829
rect 2755 9818 2761 9820
rect 2817 9818 2841 9820
rect 2897 9818 2921 9820
rect 2977 9818 3001 9820
rect 3057 9818 3063 9820
rect 2817 9766 2819 9818
rect 2999 9766 3001 9818
rect 2755 9764 2761 9766
rect 2817 9764 2841 9766
rect 2897 9764 2921 9766
rect 2977 9764 3001 9766
rect 3057 9764 3063 9766
rect 2755 9755 3063 9764
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 3160 9178 3188 10424
rect 3436 10198 3464 16079
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3528 14890 3556 15914
rect 3620 15570 3648 15982
rect 4172 15570 4200 17138
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4264 16522 4292 17070
rect 4356 16726 4384 17070
rect 4816 16794 4844 17070
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 5000 16794 5028 17002
rect 5112 16892 5420 16901
rect 5112 16890 5118 16892
rect 5174 16890 5198 16892
rect 5254 16890 5278 16892
rect 5334 16890 5358 16892
rect 5414 16890 5420 16892
rect 5174 16838 5176 16890
rect 5356 16838 5358 16890
rect 5112 16836 5118 16838
rect 5174 16836 5198 16838
rect 5254 16836 5278 16838
rect 5334 16836 5358 16838
rect 5414 16836 5420 16838
rect 5112 16827 5420 16836
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 4344 16720 4396 16726
rect 4344 16662 4396 16668
rect 5000 16658 5028 16730
rect 5736 16658 5764 18022
rect 6104 16794 6132 18022
rect 6288 17814 6316 18022
rect 6276 17808 6328 17814
rect 6276 17750 6328 17756
rect 8404 17746 8432 18158
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 6276 17604 6328 17610
rect 6276 17546 6328 17552
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6288 16658 6316 17546
rect 6564 16794 6592 17682
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 5000 16250 5028 16594
rect 5552 16250 5580 16594
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 5920 16250 5948 16526
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5112 15804 5420 15813
rect 5112 15802 5118 15804
rect 5174 15802 5198 15804
rect 5254 15802 5278 15804
rect 5334 15802 5358 15804
rect 5414 15802 5420 15804
rect 5174 15750 5176 15802
rect 5356 15750 5358 15802
rect 5112 15748 5118 15750
rect 5174 15748 5198 15750
rect 5254 15748 5278 15750
rect 5334 15748 5358 15750
rect 5414 15748 5420 15750
rect 5112 15739 5420 15748
rect 3608 15564 3660 15570
rect 3608 15506 3660 15512
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 5356 15360 5408 15366
rect 5460 15348 5488 15846
rect 5552 15706 5580 16186
rect 6012 16114 6040 16594
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 6288 15434 6316 15846
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 5408 15320 5488 15348
rect 5356 15302 5408 15308
rect 5368 14890 5396 15302
rect 3516 14884 3568 14890
rect 3516 14826 3568 14832
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3528 12374 3556 13194
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3528 10810 3556 12174
rect 3620 12102 3648 12378
rect 3896 12306 3924 12582
rect 3988 12306 4016 12922
rect 4172 12782 4200 13398
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4264 12850 4292 13262
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4264 12730 4292 12786
rect 4264 12702 4384 12730
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11801 3648 12038
rect 3896 11898 3924 12242
rect 4264 12170 4292 12582
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3606 11792 3662 11801
rect 3606 11727 3662 11736
rect 3988 11694 4016 12038
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3988 11218 4016 11630
rect 4356 11286 4384 12702
rect 4448 12434 4476 14214
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4540 13394 4568 13670
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4540 12782 4568 13330
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4448 12406 4568 12434
rect 4436 12164 4488 12170
rect 4436 12106 4488 12112
rect 4448 11762 4476 12106
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1412 7954 1440 8570
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1308 7812 1360 7818
rect 1308 7754 1360 7760
rect 1228 7500 1348 7528
rect 1124 6860 1176 6866
rect 1124 6802 1176 6808
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1124 6656 1176 6662
rect 1044 6616 1124 6644
rect 1044 6390 1072 6616
rect 1124 6598 1176 6604
rect 1032 6384 1084 6390
rect 1032 6326 1084 6332
rect 940 6248 992 6254
rect 940 6190 992 6196
rect 1228 6118 1256 6802
rect 1320 6254 1348 7500
rect 1504 6866 1532 8910
rect 1688 8430 1716 8978
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 8090 1716 8366
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1596 7546 1624 7890
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1400 6724 1452 6730
rect 1400 6666 1452 6672
rect 1412 6458 1440 6666
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1596 6254 1624 6598
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1216 6112 1268 6118
rect 1216 6054 1268 6060
rect 1308 6112 1360 6118
rect 1308 6054 1360 6060
rect 1228 5710 1256 6054
rect 1320 5914 1348 6054
rect 1872 5914 1900 6190
rect 1964 5914 1992 9114
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2962 8936 3018 8945
rect 2608 8498 2636 8910
rect 2962 8871 3018 8880
rect 2976 8838 3004 8871
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2755 8732 3063 8741
rect 2755 8730 2761 8732
rect 2817 8730 2841 8732
rect 2897 8730 2921 8732
rect 2977 8730 3001 8732
rect 3057 8730 3063 8732
rect 2817 8678 2819 8730
rect 2999 8678 3001 8730
rect 2755 8676 2761 8678
rect 2817 8676 2841 8678
rect 2897 8676 2921 8678
rect 2977 8676 3001 8678
rect 3057 8676 3063 8678
rect 2755 8667 3063 8676
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 2056 7886 2084 8230
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7206 2084 7822
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 2148 7546 2176 7754
rect 2608 7546 2636 8434
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 2755 7644 3063 7653
rect 2755 7642 2761 7644
rect 2817 7642 2841 7644
rect 2897 7642 2921 7644
rect 2977 7642 3001 7644
rect 3057 7642 3063 7644
rect 2817 7590 2819 7642
rect 2999 7590 3001 7642
rect 2755 7588 2761 7590
rect 2817 7588 2841 7590
rect 2897 7588 2921 7590
rect 2977 7588 3001 7590
rect 3057 7588 3063 7590
rect 2755 7579 3063 7588
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2608 6866 2636 7278
rect 2884 7206 2912 7482
rect 3160 7206 3188 7890
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3252 7274 3280 7822
rect 3344 7546 3372 8026
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2608 6118 2636 6802
rect 3160 6662 3188 7142
rect 3252 7002 3280 7210
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2755 6556 3063 6565
rect 2755 6554 2761 6556
rect 2817 6554 2841 6556
rect 2897 6554 2921 6556
rect 2977 6554 3001 6556
rect 3057 6554 3063 6556
rect 2817 6502 2819 6554
rect 2999 6502 3001 6554
rect 2755 6500 2761 6502
rect 2817 6500 2841 6502
rect 2897 6500 2921 6502
rect 2977 6500 3001 6502
rect 3057 6500 3063 6502
rect 2755 6491 3063 6500
rect 3160 6254 3188 6598
rect 3252 6458 3280 6938
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 3344 5914 3372 7482
rect 4080 7410 4108 7754
rect 4172 7410 4200 9046
rect 4540 9042 4568 12406
rect 4632 9518 4660 14758
rect 5112 14716 5420 14725
rect 5112 14714 5118 14716
rect 5174 14714 5198 14716
rect 5254 14714 5278 14716
rect 5334 14714 5358 14716
rect 5414 14714 5420 14716
rect 5174 14662 5176 14714
rect 5356 14662 5358 14714
rect 5112 14660 5118 14662
rect 5174 14660 5198 14662
rect 5254 14660 5278 14662
rect 5334 14660 5358 14662
rect 5414 14660 5420 14662
rect 5112 14651 5420 14660
rect 5920 14618 5948 14826
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5920 13870 5948 14418
rect 6288 14346 6316 14758
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5112 13628 5420 13637
rect 5112 13626 5118 13628
rect 5174 13626 5198 13628
rect 5254 13626 5278 13628
rect 5334 13626 5358 13628
rect 5414 13626 5420 13628
rect 5174 13574 5176 13626
rect 5356 13574 5358 13626
rect 5112 13572 5118 13574
rect 5174 13572 5198 13574
rect 5254 13572 5278 13574
rect 5334 13572 5358 13574
rect 5414 13572 5420 13574
rect 5112 13563 5420 13572
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4724 12374 4752 12786
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4908 12238 4936 13330
rect 5644 12986 5672 13806
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6104 13394 6132 13466
rect 6288 13394 6316 13738
rect 6380 13394 6408 14758
rect 6472 14618 6500 15506
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6564 15162 6592 15438
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6656 14498 6684 16390
rect 6748 15178 6776 17478
rect 6840 17338 6868 17478
rect 7470 17436 7778 17445
rect 7470 17434 7476 17436
rect 7532 17434 7556 17436
rect 7612 17434 7636 17436
rect 7692 17434 7716 17436
rect 7772 17434 7778 17436
rect 7532 17382 7534 17434
rect 7714 17382 7716 17434
rect 7470 17380 7476 17382
rect 7532 17380 7556 17382
rect 7612 17380 7636 17382
rect 7692 17380 7716 17382
rect 7772 17380 7778 17382
rect 7470 17371 7778 17380
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 8128 17134 8156 17682
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 7760 16658 7788 17002
rect 7944 16794 7972 17070
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6840 15978 6868 16390
rect 7470 16348 7778 16357
rect 7470 16346 7476 16348
rect 7532 16346 7556 16348
rect 7612 16346 7636 16348
rect 7692 16346 7716 16348
rect 7772 16346 7778 16348
rect 7532 16294 7534 16346
rect 7714 16294 7716 16346
rect 7470 16292 7476 16294
rect 7532 16292 7556 16294
rect 7612 16292 7636 16294
rect 7692 16292 7716 16294
rect 7772 16292 7778 16294
rect 7470 16283 7778 16292
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7576 15706 7604 15914
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7852 15706 7880 15846
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 6748 15150 6868 15178
rect 6472 14470 6684 14498
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5112 12540 5420 12549
rect 5112 12538 5118 12540
rect 5174 12538 5198 12540
rect 5254 12538 5278 12540
rect 5334 12538 5358 12540
rect 5414 12538 5420 12540
rect 5174 12486 5176 12538
rect 5356 12486 5358 12538
rect 5112 12484 5118 12486
rect 5174 12484 5198 12486
rect 5254 12484 5278 12486
rect 5334 12484 5358 12486
rect 5414 12484 5420 12486
rect 5112 12475 5420 12484
rect 5460 12442 5488 12650
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5644 12306 5672 12922
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4724 11830 4752 12038
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 4724 11626 4752 11766
rect 4816 11694 4844 12038
rect 5092 11694 5120 12242
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5736 11762 5764 12038
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 4724 11218 4752 11562
rect 5000 11218 5028 11562
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 5112 11452 5420 11461
rect 5112 11450 5118 11452
rect 5174 11450 5198 11452
rect 5254 11450 5278 11452
rect 5334 11450 5358 11452
rect 5414 11450 5420 11452
rect 5174 11398 5176 11450
rect 5356 11398 5358 11450
rect 5112 11396 5118 11398
rect 5174 11396 5198 11398
rect 5254 11396 5278 11398
rect 5334 11396 5358 11398
rect 5414 11396 5420 11398
rect 5112 11387 5420 11396
rect 5828 11218 5856 11494
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5000 10674 5028 11154
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5112 10364 5420 10373
rect 5112 10362 5118 10364
rect 5174 10362 5198 10364
rect 5254 10362 5278 10364
rect 5334 10362 5358 10364
rect 5414 10362 5420 10364
rect 5174 10310 5176 10362
rect 5356 10310 5358 10362
rect 5112 10308 5118 10310
rect 5174 10308 5198 10310
rect 5254 10308 5278 10310
rect 5334 10308 5358 10310
rect 5414 10308 5420 10310
rect 5112 10299 5420 10308
rect 5460 10130 5488 10950
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5644 10470 5672 10542
rect 6012 10470 6040 10950
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5644 10266 5672 10406
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4804 9512 4856 9518
rect 5540 9512 5592 9518
rect 4804 9454 4856 9460
rect 5262 9480 5318 9489
rect 4816 9178 4844 9454
rect 5540 9454 5592 9460
rect 5262 9415 5264 9424
rect 5316 9415 5318 9424
rect 5264 9386 5316 9392
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4908 9058 4936 9318
rect 5112 9276 5420 9285
rect 5112 9274 5118 9276
rect 5174 9274 5198 9276
rect 5254 9274 5278 9276
rect 5334 9274 5358 9276
rect 5414 9274 5420 9276
rect 5174 9222 5176 9274
rect 5356 9222 5358 9274
rect 5112 9220 5118 9222
rect 5174 9220 5198 9222
rect 5254 9220 5278 9222
rect 5334 9220 5358 9222
rect 5414 9220 5420 9222
rect 5112 9211 5420 9220
rect 5354 9072 5410 9081
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4804 9036 4856 9042
rect 4908 9030 5354 9058
rect 5354 9007 5356 9016
rect 4804 8978 4856 8984
rect 5408 9007 5410 9016
rect 5460 9024 5488 9318
rect 5552 9178 5580 9454
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5644 9042 5672 10202
rect 6012 10130 6040 10406
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5722 10024 5778 10033
rect 5722 9959 5778 9968
rect 5736 9518 5764 9959
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5632 9036 5684 9042
rect 5460 8996 5580 9024
rect 5356 8978 5408 8984
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4724 8634 4752 8910
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4632 8090 4660 8366
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4528 8016 4580 8022
rect 4724 7970 4752 8230
rect 4580 7964 4752 7970
rect 4528 7958 4752 7964
rect 4540 7942 4752 7958
rect 4724 7886 4752 7942
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4540 7750 4568 7822
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4080 7002 4108 7346
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4172 6866 4200 7346
rect 4356 6882 4384 7686
rect 4540 7478 4568 7686
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4160 6860 4212 6866
rect 4356 6854 4476 6882
rect 4160 6802 4212 6808
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3528 6458 3556 6666
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 1308 5908 1360 5914
rect 1308 5850 1360 5856
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 1216 5704 1268 5710
rect 1216 5646 1268 5652
rect 1228 5166 1256 5646
rect 1320 5166 1348 5850
rect 3344 5794 3372 5850
rect 3344 5778 3464 5794
rect 1860 5772 1912 5778
rect 3344 5772 3476 5778
rect 3344 5766 3424 5772
rect 1860 5714 1912 5720
rect 3424 5714 3476 5720
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1216 5160 1268 5166
rect 1216 5102 1268 5108
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4826 1348 5102
rect 1308 4820 1360 4826
rect 1308 4762 1360 4768
rect 1412 4690 1440 5170
rect 1504 4690 1532 5306
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1124 4480 1176 4486
rect 1124 4422 1176 4428
rect 1136 4078 1164 4422
rect 1412 4282 1440 4626
rect 1596 4622 1624 4966
rect 1688 4826 1716 5510
rect 1872 5370 1900 5714
rect 3528 5574 3556 6258
rect 3988 6254 4016 6598
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 4172 5778 4200 6802
rect 4448 6662 4476 6854
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1964 5098 1992 5510
rect 2755 5468 3063 5477
rect 2755 5466 2761 5468
rect 2817 5466 2841 5468
rect 2897 5466 2921 5468
rect 2977 5466 3001 5468
rect 3057 5466 3063 5468
rect 2817 5414 2819 5466
rect 2999 5414 3001 5466
rect 2755 5412 2761 5414
rect 2817 5412 2841 5414
rect 2897 5412 2921 5414
rect 2977 5412 3001 5414
rect 3057 5412 3063 5414
rect 2755 5403 3063 5412
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3068 5137 3096 5170
rect 3054 5128 3110 5137
rect 1952 5092 2004 5098
rect 4080 5098 4108 5510
rect 4264 5166 4292 6122
rect 4448 5710 4476 6598
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 3054 5063 3110 5072
rect 4068 5092 4120 5098
rect 1952 5034 2004 5040
rect 4068 5034 4120 5040
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 1688 4162 1716 4762
rect 1964 4214 1992 5034
rect 4448 4690 4476 5646
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 1596 4134 1716 4162
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 1124 4072 1176 4078
rect 1124 4014 1176 4020
rect 1400 4072 1452 4078
rect 1596 4026 1624 4134
rect 1452 4020 1624 4026
rect 1400 4014 1624 4020
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1308 4004 1360 4010
rect 1412 3998 1624 4014
rect 1308 3946 1360 3952
rect 1124 3936 1176 3942
rect 1124 3878 1176 3884
rect 1136 3738 1164 3878
rect 1124 3732 1176 3738
rect 1124 3674 1176 3680
rect 1136 1986 1164 3674
rect 1320 3602 1348 3946
rect 1308 3596 1360 3602
rect 1308 3538 1360 3544
rect 1320 2990 1348 3538
rect 1596 3534 1624 3998
rect 1688 3738 1716 4014
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1676 3528 1728 3534
rect 1964 3482 1992 4150
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1676 3470 1728 3476
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 1688 2854 1716 3470
rect 1872 3466 1992 3482
rect 1860 3460 1992 3466
rect 1912 3454 1992 3460
rect 1860 3402 1912 3408
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1216 2848 1268 2854
rect 1492 2848 1544 2854
rect 1268 2796 1348 2802
rect 1216 2790 1348 2796
rect 1492 2790 1544 2796
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1228 2774 1348 2790
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 1228 2106 1256 2450
rect 1320 2446 1348 2774
rect 1504 2650 1532 2790
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 1504 2514 1532 2586
rect 1492 2508 1544 2514
rect 1492 2450 1544 2456
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 1400 2304 1452 2310
rect 1400 2246 1452 2252
rect 1412 2106 1440 2246
rect 1216 2100 1268 2106
rect 1216 2042 1268 2048
rect 1400 2100 1452 2106
rect 1400 2042 1452 2048
rect 1136 1958 1256 1986
rect 1228 1902 1256 1958
rect 1216 1896 1268 1902
rect 1216 1838 1268 1844
rect 1412 1562 1440 2042
rect 1492 1760 1544 1766
rect 1492 1702 1544 1708
rect 1504 1562 1532 1702
rect 1400 1556 1452 1562
rect 1400 1498 1452 1504
rect 1492 1556 1544 1562
rect 1492 1498 1544 1504
rect 1688 1358 1716 2790
rect 1780 2582 1808 3334
rect 1872 3194 1900 3402
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 2056 3074 2084 3878
rect 2608 3670 2636 4422
rect 2755 4380 3063 4389
rect 2755 4378 2761 4380
rect 2817 4378 2841 4380
rect 2897 4378 2921 4380
rect 2977 4378 3001 4380
rect 3057 4378 3063 4380
rect 2817 4326 2819 4378
rect 2999 4326 3001 4378
rect 2755 4324 2761 4326
rect 2817 4324 2841 4326
rect 2897 4324 2921 4326
rect 2977 4324 3001 4326
rect 3057 4324 3063 4326
rect 2755 4315 3063 4324
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 2240 3398 2268 3538
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2755 3292 3063 3301
rect 2755 3290 2761 3292
rect 2817 3290 2841 3292
rect 2897 3290 2921 3292
rect 2977 3290 3001 3292
rect 3057 3290 3063 3292
rect 2817 3238 2819 3290
rect 2999 3238 3001 3290
rect 2755 3236 2761 3238
rect 2817 3236 2841 3238
rect 2897 3236 2921 3238
rect 2977 3236 3001 3238
rect 3057 3236 3063 3238
rect 2755 3227 3063 3236
rect 1872 3046 2084 3074
rect 1872 2582 1900 3046
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 1952 2916 2004 2922
rect 1952 2858 2004 2864
rect 1964 2650 1992 2858
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 1768 2576 1820 2582
rect 1768 2518 1820 2524
rect 1860 2576 1912 2582
rect 1860 2518 1912 2524
rect 2240 2514 2268 2926
rect 2412 2916 2464 2922
rect 2412 2858 2464 2864
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2424 1970 2452 2858
rect 3712 2650 3740 3538
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4632 2650 4660 3402
rect 4816 3194 4844 8978
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5184 8430 5212 8842
rect 5172 8424 5224 8430
rect 5460 8412 5488 8842
rect 5552 8838 5580 8996
rect 5632 8978 5684 8984
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5540 8424 5592 8430
rect 5460 8384 5540 8412
rect 5172 8366 5224 8372
rect 5540 8366 5592 8372
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5112 8188 5420 8197
rect 5112 8186 5118 8188
rect 5174 8186 5198 8188
rect 5254 8186 5278 8188
rect 5334 8186 5358 8188
rect 5414 8186 5420 8188
rect 5174 8134 5176 8186
rect 5356 8134 5358 8186
rect 5112 8132 5118 8134
rect 5174 8132 5198 8134
rect 5254 8132 5278 8134
rect 5334 8132 5358 8134
rect 5414 8132 5420 8134
rect 5112 8123 5420 8132
rect 5460 7954 5488 8230
rect 5552 8090 5580 8366
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4908 7342 4936 7754
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4908 7206 4936 7278
rect 5460 7274 5488 7890
rect 5644 7342 5672 8570
rect 5736 8090 5764 9318
rect 5920 9178 5948 9862
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 6012 8838 6040 9590
rect 6104 9330 6132 11494
rect 6380 11014 6408 13126
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6472 10810 6500 14470
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6564 13394 6592 14010
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6196 9926 6224 9998
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6196 9518 6224 9862
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6184 9376 6236 9382
rect 6104 9324 6184 9330
rect 6104 9318 6236 9324
rect 6104 9302 6224 9318
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 6012 8634 6040 8774
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5920 7546 5948 8366
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 6934 4936 7142
rect 5000 6984 5028 7210
rect 5112 7100 5420 7109
rect 5112 7098 5118 7100
rect 5174 7098 5198 7100
rect 5254 7098 5278 7100
rect 5334 7098 5358 7100
rect 5414 7098 5420 7100
rect 5174 7046 5176 7098
rect 5356 7046 5358 7098
rect 5112 7044 5118 7046
rect 5174 7044 5198 7046
rect 5254 7044 5278 7046
rect 5334 7044 5358 7046
rect 5414 7044 5420 7046
rect 5112 7035 5420 7044
rect 5172 6996 5224 7002
rect 5000 6956 5172 6984
rect 5172 6938 5224 6944
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4908 6254 4936 6870
rect 5184 6254 5212 6938
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5460 6390 5488 6598
rect 5552 6458 5580 6598
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 6012 6254 6040 7278
rect 6196 6866 6224 9302
rect 6274 9072 6330 9081
rect 6274 9007 6276 9016
rect 6328 9007 6330 9016
rect 6276 8978 6328 8984
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6288 8430 6316 8774
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6288 7818 6316 8366
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 6000 6248 6052 6254
rect 6052 6196 6132 6202
rect 6000 6190 6132 6196
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5112 6012 5420 6021
rect 5112 6010 5118 6012
rect 5174 6010 5198 6012
rect 5254 6010 5278 6012
rect 5334 6010 5358 6012
rect 5414 6010 5420 6012
rect 5174 5958 5176 6010
rect 5356 5958 5358 6010
rect 5112 5956 5118 5958
rect 5174 5956 5198 5958
rect 5254 5956 5278 5958
rect 5334 5956 5358 5958
rect 5414 5956 5420 5958
rect 5112 5947 5420 5956
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4908 3738 4936 5782
rect 5460 5166 5488 6054
rect 5736 5778 5764 6190
rect 5908 6180 5960 6186
rect 6012 6174 6132 6190
rect 5908 6122 5960 6128
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5000 4146 5028 5102
rect 5112 4924 5420 4933
rect 5112 4922 5118 4924
rect 5174 4922 5198 4924
rect 5254 4922 5278 4924
rect 5334 4922 5358 4924
rect 5414 4922 5420 4924
rect 5174 4870 5176 4922
rect 5356 4870 5358 4922
rect 5112 4868 5118 4870
rect 5174 4868 5198 4870
rect 5254 4868 5278 4870
rect 5334 4868 5358 4870
rect 5414 4868 5420 4870
rect 5112 4859 5420 4868
rect 5828 4826 5856 5714
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5112 3836 5420 3845
rect 5112 3834 5118 3836
rect 5174 3834 5198 3836
rect 5254 3834 5278 3836
rect 5334 3834 5358 3836
rect 5414 3834 5420 3836
rect 5174 3782 5176 3834
rect 5356 3782 5358 3834
rect 5112 3780 5118 3782
rect 5174 3780 5198 3782
rect 5254 3780 5278 3782
rect 5334 3780 5358 3782
rect 5414 3780 5420 3782
rect 5112 3771 5420 3780
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5460 3602 5488 3946
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5112 2748 5420 2757
rect 5112 2746 5118 2748
rect 5174 2746 5198 2748
rect 5254 2746 5278 2748
rect 5334 2746 5358 2748
rect 5414 2746 5420 2748
rect 5174 2694 5176 2746
rect 5356 2694 5358 2746
rect 5112 2692 5118 2694
rect 5174 2692 5198 2694
rect 5254 2692 5278 2694
rect 5334 2692 5358 2694
rect 5414 2692 5420 2694
rect 5112 2683 5420 2692
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2516 2106 2544 2450
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2504 2100 2556 2106
rect 2504 2042 2556 2048
rect 2228 1964 2280 1970
rect 2228 1906 2280 1912
rect 2412 1964 2464 1970
rect 2412 1906 2464 1912
rect 2044 1488 2096 1494
rect 2044 1430 2096 1436
rect 1676 1352 1728 1358
rect 1676 1294 1728 1300
rect 1952 944 2004 950
rect 1952 886 2004 892
rect 848 808 900 814
rect 676 768 848 796
rect 676 400 704 768
rect 848 750 900 756
rect 1308 808 1360 814
rect 1308 750 1360 756
rect 1320 400 1348 750
rect 1964 400 1992 886
rect 2056 882 2084 1430
rect 2240 1018 2268 1906
rect 2608 1902 2636 2246
rect 2755 2204 3063 2213
rect 2755 2202 2761 2204
rect 2817 2202 2841 2204
rect 2897 2202 2921 2204
rect 2977 2202 3001 2204
rect 3057 2202 3063 2204
rect 2817 2150 2819 2202
rect 2999 2150 3001 2202
rect 2755 2148 2761 2150
rect 2817 2148 2841 2150
rect 2897 2148 2921 2150
rect 2977 2148 3001 2150
rect 3057 2148 3063 2150
rect 2755 2139 3063 2148
rect 2780 2100 2832 2106
rect 2780 2042 2832 2048
rect 2792 1902 2820 2042
rect 3252 1970 3280 2518
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3528 2106 3556 2246
rect 3516 2100 3568 2106
rect 3516 2042 3568 2048
rect 3240 1964 3292 1970
rect 3240 1906 3292 1912
rect 2596 1896 2648 1902
rect 2596 1838 2648 1844
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 2688 1760 2740 1766
rect 2740 1708 2820 1714
rect 2688 1702 2820 1708
rect 2700 1686 2820 1702
rect 2792 1290 2820 1686
rect 3252 1494 3280 1906
rect 3528 1902 3556 2042
rect 3516 1896 3568 1902
rect 3516 1838 3568 1844
rect 3240 1488 3292 1494
rect 3240 1430 3292 1436
rect 3620 1306 3648 2450
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 3712 1970 3740 2246
rect 4172 2106 4200 2586
rect 5552 2582 5580 2926
rect 5644 2650 5672 3674
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5828 2582 5856 2790
rect 5540 2576 5592 2582
rect 4908 2514 5028 2530
rect 5540 2518 5592 2524
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 4908 2508 5040 2514
rect 4908 2502 4988 2508
rect 4160 2100 4212 2106
rect 4160 2042 4212 2048
rect 3700 1964 3752 1970
rect 3700 1906 3752 1912
rect 3884 1896 3936 1902
rect 3884 1838 3936 1844
rect 4802 1864 4858 1873
rect 3896 1494 3924 1838
rect 4436 1828 4488 1834
rect 4802 1799 4858 1808
rect 4436 1770 4488 1776
rect 4448 1562 4476 1770
rect 4816 1562 4844 1799
rect 4908 1766 4936 2502
rect 4988 2450 5040 2456
rect 5552 2394 5580 2518
rect 4988 2372 5040 2378
rect 5552 2366 5672 2394
rect 4988 2314 5040 2320
rect 4896 1760 4948 1766
rect 4896 1702 4948 1708
rect 4436 1556 4488 1562
rect 4436 1498 4488 1504
rect 4804 1556 4856 1562
rect 4804 1498 4856 1504
rect 3884 1488 3936 1494
rect 3884 1430 3936 1436
rect 3344 1290 3648 1306
rect 2780 1284 2832 1290
rect 2780 1226 2832 1232
rect 3332 1284 3648 1290
rect 3384 1278 3648 1284
rect 3332 1226 3384 1232
rect 2755 1116 3063 1125
rect 2755 1114 2761 1116
rect 2817 1114 2841 1116
rect 2897 1114 2921 1116
rect 2977 1114 3001 1116
rect 3057 1114 3063 1116
rect 2817 1062 2819 1114
rect 2999 1062 3001 1114
rect 2755 1060 2761 1062
rect 2817 1060 2841 1062
rect 2897 1060 2921 1062
rect 2977 1060 3001 1062
rect 3057 1060 3063 1062
rect 2755 1051 3063 1060
rect 2228 1012 2280 1018
rect 2228 954 2280 960
rect 2044 876 2096 882
rect 2044 818 2096 824
rect 3620 814 3648 1278
rect 4908 1408 4936 1702
rect 5000 1562 5028 2314
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5112 1660 5420 1669
rect 5112 1658 5118 1660
rect 5174 1658 5198 1660
rect 5254 1658 5278 1660
rect 5334 1658 5358 1660
rect 5414 1658 5420 1660
rect 5174 1606 5176 1658
rect 5356 1606 5358 1658
rect 5112 1604 5118 1606
rect 5174 1604 5198 1606
rect 5254 1604 5278 1606
rect 5334 1604 5358 1606
rect 5414 1604 5420 1606
rect 5112 1595 5420 1604
rect 5552 1562 5580 2246
rect 5644 1902 5672 2366
rect 5632 1896 5684 1902
rect 5632 1838 5684 1844
rect 4988 1556 5040 1562
rect 4988 1498 5040 1504
rect 5540 1556 5592 1562
rect 5540 1498 5592 1504
rect 5172 1420 5224 1426
rect 4908 1380 5172 1408
rect 4908 1018 4936 1380
rect 5172 1362 5224 1368
rect 5356 1420 5408 1426
rect 5644 1408 5672 1838
rect 5828 1562 5856 2518
rect 5920 1902 5948 6122
rect 6104 5710 6132 6174
rect 6380 5914 6408 10542
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6564 7342 6592 9522
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6104 3602 6132 4558
rect 6380 3738 6408 4626
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6380 3398 6408 3538
rect 6472 3466 6500 7142
rect 6564 6254 6592 7278
rect 6656 6746 6684 14214
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6748 12374 6776 13262
rect 6840 12986 6868 15150
rect 7300 14804 7328 15506
rect 7392 15162 7420 15506
rect 7470 15260 7778 15269
rect 7470 15258 7476 15260
rect 7532 15258 7556 15260
rect 7612 15258 7636 15260
rect 7692 15258 7716 15260
rect 7772 15258 7778 15260
rect 7532 15206 7534 15258
rect 7714 15206 7716 15258
rect 7470 15204 7476 15206
rect 7532 15204 7556 15206
rect 7612 15204 7636 15206
rect 7692 15204 7716 15206
rect 7772 15204 7778 15206
rect 7470 15195 7778 15204
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7380 14816 7432 14822
rect 7300 14776 7380 14804
rect 7380 14758 7432 14764
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 13938 7328 14214
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7392 13870 7420 14758
rect 7576 14618 7604 14894
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7852 14346 7880 14894
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7470 14172 7778 14181
rect 7470 14170 7476 14172
rect 7532 14170 7556 14172
rect 7612 14170 7636 14172
rect 7692 14170 7716 14172
rect 7772 14170 7778 14172
rect 7532 14118 7534 14170
rect 7714 14118 7716 14170
rect 7470 14116 7476 14118
rect 7532 14116 7556 14118
rect 7612 14116 7636 14118
rect 7692 14116 7716 14118
rect 7772 14116 7778 14118
rect 7470 14107 7778 14116
rect 7852 14074 7880 14282
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7748 14000 7800 14006
rect 7800 13948 7880 13954
rect 7748 13942 7880 13948
rect 7760 13926 7880 13942
rect 7380 13864 7432 13870
rect 7300 13812 7380 13818
rect 7300 13806 7432 13812
rect 7300 13790 7420 13806
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 7024 13394 7052 13670
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7116 12434 7144 12718
rect 7024 12406 7144 12434
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6748 10130 6776 12310
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6748 9518 6776 10066
rect 6840 9722 6868 10066
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6920 6792 6972 6798
rect 6656 6740 6920 6746
rect 6656 6734 6972 6740
rect 6656 6718 6960 6734
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6840 5914 6868 6718
rect 7024 6118 7052 12406
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7208 10810 7236 12174
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7208 9178 7236 10746
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7116 7954 7144 8978
rect 7300 8022 7328 13790
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7392 12850 7420 13466
rect 7668 13394 7696 13670
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7470 13084 7778 13093
rect 7470 13082 7476 13084
rect 7532 13082 7556 13084
rect 7612 13082 7636 13084
rect 7692 13082 7716 13084
rect 7772 13082 7778 13084
rect 7532 13030 7534 13082
rect 7714 13030 7716 13082
rect 7470 13028 7476 13030
rect 7532 13028 7556 13030
rect 7612 13028 7636 13030
rect 7692 13028 7716 13030
rect 7772 13028 7778 13030
rect 7470 13019 7778 13028
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7852 12434 7880 13926
rect 7944 13462 7972 14486
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 8036 13274 8064 13806
rect 7392 12406 7880 12434
rect 7944 13246 8064 13274
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7116 7410 7144 7890
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7116 6730 7144 7346
rect 7392 6866 7420 12406
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7470 11996 7778 12005
rect 7470 11994 7476 11996
rect 7532 11994 7556 11996
rect 7612 11994 7636 11996
rect 7692 11994 7716 11996
rect 7772 11994 7778 11996
rect 7532 11942 7534 11994
rect 7714 11942 7716 11994
rect 7470 11940 7476 11942
rect 7532 11940 7556 11942
rect 7612 11940 7636 11942
rect 7692 11940 7716 11942
rect 7772 11940 7778 11942
rect 7470 11931 7778 11940
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7576 11354 7604 11630
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7852 11234 7880 12242
rect 7760 11218 7880 11234
rect 7748 11212 7880 11218
rect 7800 11206 7880 11212
rect 7748 11154 7800 11160
rect 7470 10908 7778 10917
rect 7470 10906 7476 10908
rect 7532 10906 7556 10908
rect 7612 10906 7636 10908
rect 7692 10906 7716 10908
rect 7772 10906 7778 10908
rect 7532 10854 7534 10906
rect 7714 10854 7716 10906
rect 7470 10852 7476 10854
rect 7532 10852 7556 10854
rect 7612 10852 7636 10854
rect 7692 10852 7716 10854
rect 7772 10852 7778 10854
rect 7470 10843 7778 10852
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 10033 7604 10066
rect 7760 10062 7788 10406
rect 7748 10056 7800 10062
rect 7562 10024 7618 10033
rect 7748 9998 7800 10004
rect 7562 9959 7618 9968
rect 7470 9820 7778 9829
rect 7470 9818 7476 9820
rect 7532 9818 7556 9820
rect 7612 9818 7636 9820
rect 7692 9818 7716 9820
rect 7772 9818 7778 9820
rect 7532 9766 7534 9818
rect 7714 9766 7716 9818
rect 7470 9764 7476 9766
rect 7532 9764 7556 9766
rect 7612 9764 7636 9766
rect 7692 9764 7716 9766
rect 7772 9764 7778 9766
rect 7470 9755 7778 9764
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7838 9480 7894 9489
rect 7668 9042 7696 9454
rect 7838 9415 7894 9424
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7470 8732 7778 8741
rect 7470 8730 7476 8732
rect 7532 8730 7556 8732
rect 7612 8730 7636 8732
rect 7692 8730 7716 8732
rect 7772 8730 7778 8732
rect 7532 8678 7534 8730
rect 7714 8678 7716 8730
rect 7470 8676 7476 8678
rect 7532 8676 7556 8678
rect 7612 8676 7636 8678
rect 7692 8676 7716 8678
rect 7772 8676 7778 8678
rect 7470 8667 7778 8676
rect 7852 8430 7880 9415
rect 7944 9110 7972 13246
rect 8128 12986 8156 16934
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8220 16250 8248 16594
rect 8404 16454 8432 17682
rect 8496 17338 8524 18090
rect 10152 18086 10180 18176
rect 10324 18158 10376 18164
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9416 17338 9444 17750
rect 9600 17338 9628 18022
rect 9827 17980 10135 17989
rect 9827 17978 9833 17980
rect 9889 17978 9913 17980
rect 9969 17978 9993 17980
rect 10049 17978 10073 17980
rect 10129 17978 10135 17980
rect 9889 17926 9891 17978
rect 10071 17926 10073 17978
rect 9827 17924 9833 17926
rect 9889 17924 9913 17926
rect 9969 17924 9993 17926
rect 10049 17924 10073 17926
rect 10129 17924 10135 17926
rect 9827 17915 10135 17924
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9692 17218 9720 17682
rect 9876 17542 9904 17818
rect 10244 17814 10272 18022
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9600 17190 9720 17218
rect 9324 16998 9352 17138
rect 9600 17134 9628 17190
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9588 17128 9640 17134
rect 9784 17082 9812 17478
rect 10152 17338 10180 17682
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 9588 17070 9640 17076
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8404 16046 8432 16390
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8220 14006 8248 14894
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 8036 12434 8064 12718
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8036 12406 8156 12434
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 10674 8064 11494
rect 8128 11370 8156 12406
rect 8220 12102 8248 12582
rect 8312 12434 8340 15302
rect 8404 14414 8432 15982
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8588 14278 8616 14894
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8956 14498 8984 14758
rect 8864 14482 8984 14498
rect 9048 14482 9076 14894
rect 8852 14476 8984 14482
rect 8904 14470 8984 14476
rect 8852 14418 8904 14424
rect 8668 14340 8720 14346
rect 8668 14282 8720 14288
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8588 13870 8616 14214
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8588 13462 8616 13806
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8680 13394 8708 14282
rect 8956 13938 8984 14470
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9140 14362 9168 15914
rect 9048 14334 9168 14362
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 9048 13734 9076 14334
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 13870 9168 14214
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8312 12406 8432 12434
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8128 11342 8248 11370
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8128 10674 8156 11222
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7470 7644 7778 7653
rect 7470 7642 7476 7644
rect 7532 7642 7556 7644
rect 7612 7642 7636 7644
rect 7692 7642 7716 7644
rect 7772 7642 7778 7644
rect 7532 7590 7534 7642
rect 7714 7590 7716 7642
rect 7470 7588 7476 7590
rect 7532 7588 7556 7590
rect 7612 7588 7636 7590
rect 7692 7588 7716 7590
rect 7772 7588 7778 7590
rect 7470 7579 7778 7588
rect 8220 7546 8248 11342
rect 8404 8430 8432 12406
rect 8588 8634 8616 13126
rect 8760 12776 8812 12782
rect 8666 12744 8722 12753
rect 8760 12718 8812 12724
rect 8666 12679 8668 12688
rect 8720 12679 8722 12688
rect 8668 12650 8720 12656
rect 8666 12336 8722 12345
rect 8666 12271 8722 12280
rect 8680 11694 8708 12271
rect 8772 11694 8800 12718
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 9048 9178 9076 13670
rect 9140 9518 9168 13806
rect 9324 12850 9352 16186
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9416 14958 9444 15098
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9508 14498 9536 17070
rect 9692 17054 9812 17082
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9600 14958 9628 15030
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9600 14618 9628 14758
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9508 14470 9628 14498
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9232 12442 9260 12718
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9508 12306 9536 12582
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9232 9722 9260 11630
rect 9508 11626 9536 12242
rect 9600 12238 9628 14470
rect 9584 12232 9636 12238
rect 9584 12174 9636 12180
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 8036 6934 8064 7142
rect 8404 7002 8432 7686
rect 8496 7410 8524 8230
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7116 6458 7144 6666
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 7116 5778 7144 6394
rect 7300 6361 7328 6598
rect 7286 6352 7342 6361
rect 7286 6287 7342 6296
rect 7392 6254 7420 6802
rect 7470 6556 7778 6565
rect 7470 6554 7476 6556
rect 7532 6554 7556 6556
rect 7612 6554 7636 6556
rect 7692 6554 7716 6556
rect 7772 6554 7778 6556
rect 7532 6502 7534 6554
rect 7714 6502 7716 6554
rect 7470 6500 7476 6502
rect 7532 6500 7556 6502
rect 7612 6500 7636 6502
rect 7692 6500 7716 6502
rect 7772 6500 7778 6502
rect 7470 6491 7778 6500
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 6748 5302 6776 5714
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6840 4146 6868 5714
rect 7470 5468 7778 5477
rect 7470 5466 7476 5468
rect 7532 5466 7556 5468
rect 7612 5466 7636 5468
rect 7692 5466 7716 5468
rect 7772 5466 7778 5468
rect 7532 5414 7534 5466
rect 7714 5414 7716 5466
rect 7470 5412 7476 5414
rect 7532 5412 7556 5414
rect 7612 5412 7636 5414
rect 7692 5412 7716 5414
rect 7772 5412 7778 5414
rect 7470 5403 7778 5412
rect 7852 5370 7880 6122
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7944 5370 7972 5510
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 8036 5234 8064 6870
rect 8496 6866 8524 7346
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8392 6860 8444 6866
rect 8312 6820 8392 6848
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5914 8248 6054
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7470 4380 7778 4389
rect 7470 4378 7476 4380
rect 7532 4378 7556 4380
rect 7612 4378 7636 4380
rect 7692 4378 7716 4380
rect 7772 4378 7778 4380
rect 7532 4326 7534 4378
rect 7714 4326 7716 4378
rect 7470 4324 7476 4326
rect 7532 4324 7556 4326
rect 7612 4324 7636 4326
rect 7692 4324 7716 4326
rect 7772 4324 7778 4326
rect 7470 4315 7778 4324
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6380 2990 6408 3334
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6380 2650 6408 2926
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6564 2514 6592 3470
rect 7300 3194 7328 3946
rect 7470 3292 7778 3301
rect 7470 3290 7476 3292
rect 7532 3290 7556 3292
rect 7612 3290 7636 3292
rect 7692 3290 7716 3292
rect 7772 3290 7778 3292
rect 7532 3238 7534 3290
rect 7714 3238 7716 3290
rect 7470 3236 7476 3238
rect 7532 3236 7556 3238
rect 7612 3236 7636 3238
rect 7692 3236 7716 3238
rect 7772 3236 7778 3238
rect 7470 3227 7778 3236
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 5816 1556 5868 1562
rect 5816 1498 5868 1504
rect 5408 1380 5672 1408
rect 5356 1362 5408 1368
rect 6104 1290 6132 2246
rect 6380 1426 6408 2450
rect 6368 1420 6420 1426
rect 6368 1362 6420 1368
rect 6564 1358 6592 2450
rect 6932 1970 6960 2790
rect 7668 2774 7696 2926
rect 7668 2746 7880 2774
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7012 2100 7064 2106
rect 7012 2042 7064 2048
rect 6920 1964 6972 1970
rect 6920 1906 6972 1912
rect 6932 1494 6960 1906
rect 6920 1488 6972 1494
rect 6920 1430 6972 1436
rect 6552 1352 6604 1358
rect 6552 1294 6604 1300
rect 6092 1284 6144 1290
rect 6092 1226 6144 1232
rect 4896 1012 4948 1018
rect 4896 954 4948 960
rect 6932 814 6960 1430
rect 7024 1426 7052 2042
rect 7196 1896 7248 1902
rect 7196 1838 7248 1844
rect 7208 1426 7236 1838
rect 7392 1766 7420 2586
rect 7470 2204 7778 2213
rect 7470 2202 7476 2204
rect 7532 2202 7556 2204
rect 7612 2202 7636 2204
rect 7692 2202 7716 2204
rect 7772 2202 7778 2204
rect 7532 2150 7534 2202
rect 7714 2150 7716 2202
rect 7470 2148 7476 2150
rect 7532 2148 7556 2150
rect 7612 2148 7636 2150
rect 7692 2148 7716 2150
rect 7772 2148 7778 2150
rect 7470 2139 7778 2148
rect 7472 2100 7524 2106
rect 7524 2060 7604 2088
rect 7472 2042 7524 2048
rect 7576 1970 7604 2060
rect 7852 1970 7880 2746
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8220 2310 8248 2382
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8220 2106 8248 2246
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 7840 1964 7892 1970
rect 7840 1906 7892 1912
rect 7380 1760 7432 1766
rect 7380 1702 7432 1708
rect 8312 1562 8340 6820
rect 8392 6802 8444 6808
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8404 4486 8432 6190
rect 8496 5930 8524 6802
rect 8588 6118 8616 7142
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8496 5902 8616 5930
rect 8588 5778 8616 5902
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8496 4826 8524 5714
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8680 3942 8708 8298
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8772 3754 8800 8978
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 8430 8892 8774
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 9048 8090 9076 9114
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9232 8838 9260 8978
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9324 8566 9352 11494
rect 9416 11014 9444 11494
rect 9600 11354 9628 11630
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9692 11234 9720 17054
rect 9827 16892 10135 16901
rect 9827 16890 9833 16892
rect 9889 16890 9913 16892
rect 9969 16890 9993 16892
rect 10049 16890 10073 16892
rect 10129 16890 10135 16892
rect 9889 16838 9891 16890
rect 10071 16838 10073 16890
rect 9827 16836 9833 16838
rect 9889 16836 9913 16838
rect 9969 16836 9993 16838
rect 10049 16836 10073 16838
rect 10129 16836 10135 16838
rect 9827 16827 10135 16836
rect 9827 15804 10135 15813
rect 9827 15802 9833 15804
rect 9889 15802 9913 15804
rect 9969 15802 9993 15804
rect 10049 15802 10073 15804
rect 10129 15802 10135 15804
rect 9889 15750 9891 15802
rect 10071 15750 10073 15802
rect 9827 15748 9833 15750
rect 9889 15748 9913 15750
rect 9969 15748 9993 15750
rect 10049 15748 10073 15750
rect 10129 15748 10135 15750
rect 9827 15739 10135 15748
rect 9827 14716 10135 14725
rect 9827 14714 9833 14716
rect 9889 14714 9913 14716
rect 9969 14714 9993 14716
rect 10049 14714 10073 14716
rect 10129 14714 10135 14716
rect 9889 14662 9891 14714
rect 10071 14662 10073 14714
rect 9827 14660 9833 14662
rect 9889 14660 9913 14662
rect 9969 14660 9993 14662
rect 10049 14660 10073 14662
rect 10129 14660 10135 14662
rect 9827 14651 10135 14660
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 9827 13628 10135 13637
rect 9827 13626 9833 13628
rect 9889 13626 9913 13628
rect 9969 13626 9993 13628
rect 10049 13626 10073 13628
rect 10129 13626 10135 13628
rect 9889 13574 9891 13626
rect 10071 13574 10073 13626
rect 9827 13572 9833 13574
rect 9889 13572 9913 13574
rect 9969 13572 9993 13574
rect 10049 13572 10073 13574
rect 10129 13572 10135 13574
rect 9827 13563 10135 13572
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 12918 10088 13126
rect 10048 12912 10100 12918
rect 10140 12912 10192 12918
rect 10048 12854 10100 12860
rect 10138 12880 10140 12889
rect 10192 12880 10194 12889
rect 10138 12815 10194 12824
rect 9827 12540 10135 12549
rect 9827 12538 9833 12540
rect 9889 12538 9913 12540
rect 9969 12538 9993 12540
rect 10049 12538 10073 12540
rect 10129 12538 10135 12540
rect 9889 12486 9891 12538
rect 10071 12486 10073 12538
rect 9827 12484 9833 12486
rect 9889 12484 9913 12486
rect 9969 12484 9993 12486
rect 10049 12484 10073 12486
rect 10129 12484 10135 12486
rect 9827 12475 10135 12484
rect 10244 12434 10272 14214
rect 9876 12406 10272 12434
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9784 11665 9812 12242
rect 9876 11694 9904 12406
rect 10336 12374 10364 17546
rect 10704 17542 10732 18022
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11256 17746 11284 17818
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 17134 10732 17478
rect 11164 17338 11192 17682
rect 11348 17592 11376 18022
rect 11428 17604 11480 17610
rect 11348 17564 11428 17592
rect 11428 17546 11480 17552
rect 11440 17338 11468 17546
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10888 16794 10916 17070
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 11072 16794 11100 17002
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10796 16046 10824 16730
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 11072 15706 11100 16458
rect 11164 16454 11192 17274
rect 11532 17218 11560 17478
rect 11624 17354 11652 19600
rect 14542 19068 14850 19077
rect 14542 19066 14548 19068
rect 14604 19066 14628 19068
rect 14684 19066 14708 19068
rect 14764 19066 14788 19068
rect 14844 19066 14850 19068
rect 14604 19014 14606 19066
rect 14786 19014 14788 19066
rect 14542 19012 14548 19014
rect 14604 19012 14628 19014
rect 14684 19012 14708 19014
rect 14764 19012 14788 19014
rect 14844 19012 14850 19014
rect 14542 19003 14850 19012
rect 19257 19068 19565 19077
rect 19257 19066 19263 19068
rect 19319 19066 19343 19068
rect 19399 19066 19423 19068
rect 19479 19066 19503 19068
rect 19559 19066 19565 19068
rect 19319 19014 19321 19066
rect 19501 19014 19503 19066
rect 19257 19012 19263 19014
rect 19319 19012 19343 19014
rect 19399 19012 19423 19014
rect 19479 19012 19503 19014
rect 19559 19012 19565 19014
rect 19257 19003 19565 19012
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11624 17326 11744 17354
rect 11808 17338 11836 18158
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 11256 17190 11560 17218
rect 11612 17196 11664 17202
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11164 16046 11192 16186
rect 11152 16040 11204 16046
rect 11150 16008 11152 16017
rect 11204 16008 11206 16017
rect 11150 15943 11206 15952
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10428 12850 10456 15098
rect 10704 14958 10732 15370
rect 11072 14958 11100 15642
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 13546 10640 14758
rect 10704 14482 10732 14894
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10520 13518 10640 13546
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10060 11762 10088 12174
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9864 11688 9916 11694
rect 9770 11656 9826 11665
rect 9864 11630 9916 11636
rect 9770 11591 9826 11600
rect 10152 11608 10180 12038
rect 10336 11801 10364 12174
rect 10322 11792 10378 11801
rect 10322 11727 10378 11736
rect 10152 11580 10272 11608
rect 9827 11452 10135 11461
rect 9827 11450 9833 11452
rect 9889 11450 9913 11452
rect 9969 11450 9993 11452
rect 10049 11450 10073 11452
rect 10129 11450 10135 11452
rect 9889 11398 9891 11450
rect 10071 11398 10073 11450
rect 9827 11396 9833 11398
rect 9889 11396 9913 11398
rect 9969 11396 9993 11398
rect 10049 11396 10073 11398
rect 10129 11396 10135 11398
rect 9827 11387 10135 11396
rect 9692 11218 9812 11234
rect 9496 11212 9548 11218
rect 9692 11212 9824 11218
rect 9692 11206 9772 11212
rect 9496 11154 9548 11160
rect 9772 11154 9824 11160
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9416 8634 9444 8842
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8864 7274 8892 7822
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8956 6866 8984 7890
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9034 7304 9090 7313
rect 9034 7239 9036 7248
rect 9088 7239 9090 7248
rect 9036 7210 9088 7216
rect 9140 7041 9168 7754
rect 9126 7032 9182 7041
rect 9126 6967 9182 6976
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 8956 5914 8984 6802
rect 9140 6458 9168 6802
rect 9232 6730 9260 8366
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9324 6390 9352 8366
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9416 6866 9444 8026
rect 9508 7818 9536 11154
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10810 9720 11086
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9876 10606 9904 11018
rect 10060 10810 10088 11154
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 9680 10600 9732 10606
rect 9864 10600 9916 10606
rect 9680 10542 9732 10548
rect 9770 10568 9826 10577
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9600 9178 9628 9998
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9586 9072 9642 9081
rect 9586 9007 9642 9016
rect 9600 8634 9628 9007
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9588 8084 9640 8090
rect 9692 8072 9720 10542
rect 9864 10542 9916 10548
rect 9770 10503 9772 10512
rect 9824 10503 9826 10512
rect 9772 10474 9824 10480
rect 9827 10364 10135 10373
rect 9827 10362 9833 10364
rect 9889 10362 9913 10364
rect 9969 10362 9993 10364
rect 10049 10362 10073 10364
rect 10129 10362 10135 10364
rect 9889 10310 9891 10362
rect 10071 10310 10073 10362
rect 9827 10308 9833 10310
rect 9889 10308 9913 10310
rect 9969 10308 9993 10310
rect 10049 10308 10073 10310
rect 10129 10308 10135 10310
rect 9827 10299 10135 10308
rect 10244 9926 10272 11580
rect 10336 10606 10364 11727
rect 10428 11694 10456 12786
rect 10520 12374 10548 13518
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10612 12434 10640 13330
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10704 12617 10732 12650
rect 10690 12608 10746 12617
rect 10690 12543 10746 12552
rect 10888 12442 10916 12718
rect 10876 12436 10928 12442
rect 10612 12406 10732 12434
rect 10508 12368 10560 12374
rect 10508 12310 10560 12316
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10428 9518 10456 11630
rect 10520 11354 10548 11630
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10704 11234 10732 12406
rect 10876 12378 10928 12384
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10520 11206 10732 11234
rect 10520 10742 10548 11206
rect 10508 10736 10560 10742
rect 10508 10678 10560 10684
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 9827 9276 10135 9285
rect 9827 9274 9833 9276
rect 9889 9274 9913 9276
rect 9969 9274 9993 9276
rect 10049 9274 10073 9276
rect 10129 9274 10135 9276
rect 9889 9222 9891 9274
rect 10071 9222 10073 9274
rect 9827 9220 9833 9222
rect 9889 9220 9913 9222
rect 9969 9220 9993 9222
rect 10049 9220 10073 9222
rect 10129 9220 10135 9222
rect 9827 9211 10135 9220
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 9772 8560 9824 8566
rect 9770 8528 9772 8537
rect 9824 8528 9826 8537
rect 9770 8463 9826 8472
rect 10140 8288 10192 8294
rect 10192 8248 10272 8276
rect 10140 8230 10192 8236
rect 9827 8188 10135 8197
rect 9827 8186 9833 8188
rect 9889 8186 9913 8188
rect 9969 8186 9993 8188
rect 10049 8186 10073 8188
rect 10129 8186 10135 8188
rect 9889 8134 9891 8186
rect 10071 8134 10073 8186
rect 9827 8132 9833 8134
rect 9889 8132 9913 8134
rect 9969 8132 9993 8134
rect 10049 8132 10073 8134
rect 10129 8132 10135 8134
rect 9827 8123 10135 8132
rect 10048 8084 10100 8090
rect 9692 8044 9904 8072
rect 9588 8026 9640 8032
rect 9600 7818 9628 8026
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9586 7304 9642 7313
rect 9586 7239 9642 7248
rect 9600 7206 9628 7239
rect 9876 7206 9904 8044
rect 10048 8026 10100 8032
rect 10060 7954 10088 8026
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9968 7274 9996 7822
rect 10060 7342 10088 7890
rect 10244 7342 10272 8248
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9494 7032 9550 7041
rect 9600 7018 9628 7142
rect 9827 7100 10135 7109
rect 9827 7098 9833 7100
rect 9889 7098 9913 7100
rect 9969 7098 9993 7100
rect 10049 7098 10073 7100
rect 10129 7098 10135 7100
rect 9889 7046 9891 7098
rect 10071 7046 10073 7098
rect 9827 7044 9833 7046
rect 9889 7044 9913 7046
rect 9969 7044 9993 7046
rect 10049 7044 10073 7046
rect 10129 7044 10135 7046
rect 9827 7035 10135 7044
rect 9600 6990 9720 7018
rect 9494 6967 9550 6976
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9416 6186 9444 6598
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8944 5908 8996 5914
rect 9404 5908 9456 5914
rect 8944 5850 8996 5856
rect 9324 5868 9404 5896
rect 8864 5817 8892 5850
rect 8850 5808 8906 5817
rect 8850 5743 8906 5752
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9034 5672 9090 5681
rect 9034 5607 9090 5616
rect 9048 5574 9076 5607
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9048 4486 9076 5034
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 8852 4004 8904 4010
rect 9048 3992 9076 4422
rect 8904 3964 9076 3992
rect 8852 3946 8904 3952
rect 8772 3726 8892 3754
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 3194 8800 3538
rect 8392 3188 8444 3194
rect 8760 3188 8812 3194
rect 8392 3130 8444 3136
rect 8588 3148 8760 3176
rect 8404 2582 8432 3130
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8496 2038 8524 2246
rect 8588 2106 8616 3148
rect 8760 3130 8812 3136
rect 8864 2774 8892 3726
rect 9048 3534 9076 3964
rect 9140 3738 9168 5714
rect 9324 5681 9352 5868
rect 9404 5850 9456 5856
rect 9402 5808 9458 5817
rect 9402 5743 9404 5752
rect 9456 5743 9458 5752
rect 9404 5714 9456 5720
rect 9310 5672 9366 5681
rect 9310 5607 9366 5616
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8772 2746 8892 2774
rect 8668 2508 8720 2514
rect 8772 2496 8800 2746
rect 8720 2468 8800 2496
rect 8668 2450 8720 2456
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8576 2100 8628 2106
rect 8628 2060 8800 2088
rect 8576 2042 8628 2048
rect 8484 2032 8536 2038
rect 8484 1974 8536 1980
rect 8392 1896 8444 1902
rect 8392 1838 8444 1844
rect 8300 1556 8352 1562
rect 8300 1498 8352 1504
rect 7012 1420 7064 1426
rect 7012 1362 7064 1368
rect 7196 1420 7248 1426
rect 7196 1362 7248 1368
rect 7208 1018 7236 1362
rect 8404 1358 8432 1838
rect 8496 1562 8524 1974
rect 8772 1562 8800 2060
rect 8956 1834 8984 2246
rect 9048 1970 9076 3470
rect 9324 2582 9352 5510
rect 9416 5370 9444 5510
rect 9508 5370 9536 6967
rect 9692 6934 9720 6990
rect 9680 6928 9732 6934
rect 9586 6896 9642 6905
rect 9680 6870 9732 6876
rect 10244 6866 10272 7278
rect 9586 6831 9642 6840
rect 10232 6860 10284 6866
rect 9600 6798 9628 6831
rect 10232 6802 10284 6808
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9600 6322 9628 6394
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9600 5030 9628 6054
rect 9692 5760 9720 6190
rect 9827 6012 10135 6021
rect 9827 6010 9833 6012
rect 9889 6010 9913 6012
rect 9969 6010 9993 6012
rect 10049 6010 10073 6012
rect 10129 6010 10135 6012
rect 9889 5958 9891 6010
rect 10071 5958 10073 6010
rect 9827 5956 9833 5958
rect 9889 5956 9913 5958
rect 9969 5956 9993 5958
rect 10049 5956 10073 5958
rect 10129 5956 10135 5958
rect 9827 5947 10135 5956
rect 9692 5732 9812 5760
rect 9678 5672 9734 5681
rect 9678 5607 9680 5616
rect 9732 5607 9734 5616
rect 9680 5578 9732 5584
rect 9680 5160 9732 5166
rect 9784 5148 9812 5732
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9732 5120 9812 5148
rect 9680 5102 9732 5108
rect 9876 5098 9904 5238
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9827 4924 10135 4933
rect 9827 4922 9833 4924
rect 9889 4922 9913 4924
rect 9969 4922 9993 4924
rect 10049 4922 10073 4924
rect 10129 4922 10135 4924
rect 9889 4870 9891 4922
rect 10071 4870 10073 4922
rect 9827 4868 9833 4870
rect 9889 4868 9913 4870
rect 9969 4868 9993 4870
rect 10049 4868 10073 4870
rect 10129 4868 10135 4870
rect 9827 4859 10135 4868
rect 10244 4282 10272 5102
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 9827 3836 10135 3845
rect 9827 3834 9833 3836
rect 9889 3834 9913 3836
rect 9969 3834 9993 3836
rect 10049 3834 10073 3836
rect 10129 3834 10135 3836
rect 9889 3782 9891 3834
rect 10071 3782 10073 3834
rect 9827 3780 9833 3782
rect 9889 3780 9913 3782
rect 9969 3780 9993 3782
rect 10049 3780 10073 3782
rect 10129 3780 10135 3782
rect 9827 3771 10135 3780
rect 10336 3738 10364 8978
rect 10428 8906 10456 9318
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 7954 10456 8230
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10428 7478 10456 7890
rect 10520 7546 10548 10678
rect 10796 10606 10824 12174
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10600 10056 10652 10062
rect 10704 10033 10732 10202
rect 10600 9998 10652 10004
rect 10690 10024 10746 10033
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10428 6458 10456 7142
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10612 5642 10640 9998
rect 10690 9959 10746 9968
rect 10692 9512 10744 9518
rect 10690 9480 10692 9489
rect 10744 9480 10746 9489
rect 10796 9450 10824 10542
rect 10690 9415 10746 9424
rect 10784 9444 10836 9450
rect 10704 9042 10732 9415
rect 10784 9386 10836 9392
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10704 8090 10732 8298
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 6322 10824 7686
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10796 5817 10824 5850
rect 10782 5808 10838 5817
rect 10782 5743 10838 5752
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10520 5166 10548 5510
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10428 4826 10456 5102
rect 10612 5098 10640 5238
rect 10600 5092 10652 5098
rect 10600 5034 10652 5040
rect 10704 5030 10732 5510
rect 10888 5370 10916 11562
rect 10980 10674 11008 13126
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10980 8514 11008 10474
rect 11072 10266 11100 14486
rect 11164 12850 11192 15846
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9518 11100 9930
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11164 9178 11192 12038
rect 11256 11898 11284 17190
rect 11612 17138 11664 17144
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11440 16658 11468 17070
rect 11624 16794 11652 17138
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11348 15552 11376 16118
rect 11440 15910 11468 16594
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11520 16176 11572 16182
rect 11520 16118 11572 16124
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11532 15638 11560 16118
rect 11624 16046 11652 16526
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11520 15632 11572 15638
rect 11520 15574 11572 15580
rect 11612 15564 11664 15570
rect 11348 15524 11468 15552
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11256 10470 11284 10746
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11256 9761 11284 10406
rect 11242 9752 11298 9761
rect 11242 9687 11298 9696
rect 11348 9518 11376 14214
rect 11440 10606 11468 15524
rect 11612 15506 11664 15512
rect 11624 15162 11652 15506
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11624 14482 11652 14758
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11624 11694 11652 12582
rect 11716 11898 11744 17326
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11900 16998 11928 17682
rect 11992 17338 12020 18770
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12185 18524 12493 18533
rect 12185 18522 12191 18524
rect 12247 18522 12271 18524
rect 12327 18522 12351 18524
rect 12407 18522 12431 18524
rect 12487 18522 12493 18524
rect 12247 18470 12249 18522
rect 12429 18470 12431 18522
rect 12185 18468 12191 18470
rect 12247 18468 12271 18470
rect 12327 18468 12351 18470
rect 12407 18468 12431 18470
rect 12487 18468 12493 18470
rect 12185 18459 12493 18468
rect 12544 18426 12572 18566
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12544 17746 12572 18362
rect 13004 18086 13032 18770
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13372 17746 13400 18022
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12185 17436 12493 17445
rect 12185 17434 12191 17436
rect 12247 17434 12271 17436
rect 12327 17434 12351 17436
rect 12407 17434 12431 17436
rect 12487 17434 12493 17436
rect 12247 17382 12249 17434
rect 12429 17382 12431 17434
rect 12185 17380 12191 17382
rect 12247 17380 12271 17382
rect 12327 17380 12351 17382
rect 12407 17380 12431 17382
rect 12487 17380 12493 17382
rect 12185 17371 12493 17380
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 15570 11928 16390
rect 11992 15706 12020 16594
rect 12185 16348 12493 16357
rect 12185 16346 12191 16348
rect 12247 16346 12271 16348
rect 12327 16346 12351 16348
rect 12407 16346 12431 16348
rect 12487 16346 12493 16348
rect 12247 16294 12249 16346
rect 12429 16294 12431 16346
rect 12185 16292 12191 16294
rect 12247 16292 12271 16294
rect 12327 16292 12351 16294
rect 12407 16292 12431 16294
rect 12487 16292 12493 16294
rect 12185 16283 12493 16292
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12084 15706 12112 15846
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11808 12646 11836 15302
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11702 11792 11758 11801
rect 11702 11727 11758 11736
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11716 11506 11744 11727
rect 11900 11540 11928 15506
rect 12084 15473 12112 15506
rect 12070 15464 12126 15473
rect 12070 15399 12126 15408
rect 12176 15348 12204 15846
rect 12360 15706 12388 15982
rect 12348 15700 12400 15706
rect 12400 15660 12664 15688
rect 12348 15642 12400 15648
rect 12084 15320 12204 15348
rect 12532 15360 12584 15366
rect 12084 15094 12112 15320
rect 12532 15302 12584 15308
rect 12185 15260 12493 15269
rect 12185 15258 12191 15260
rect 12247 15258 12271 15260
rect 12327 15258 12351 15260
rect 12407 15258 12431 15260
rect 12487 15258 12493 15260
rect 12247 15206 12249 15258
rect 12429 15206 12431 15258
rect 12185 15204 12191 15206
rect 12247 15204 12271 15206
rect 12327 15204 12351 15206
rect 12407 15204 12431 15206
rect 12487 15204 12493 15206
rect 12185 15195 12493 15204
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 12084 14618 12112 14758
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12268 14482 12296 15098
rect 12544 14958 12572 15302
rect 12636 15162 12664 15660
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12728 15162 12756 15506
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12820 15162 12848 15438
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12544 14414 12572 14758
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12185 14172 12493 14181
rect 12185 14170 12191 14172
rect 12247 14170 12271 14172
rect 12327 14170 12351 14172
rect 12407 14170 12431 14172
rect 12487 14170 12493 14172
rect 12247 14118 12249 14170
rect 12429 14118 12431 14170
rect 12185 14116 12191 14118
rect 12247 14116 12271 14118
rect 12327 14116 12351 14118
rect 12407 14116 12431 14118
rect 12487 14116 12493 14118
rect 12185 14107 12493 14116
rect 12544 13326 12572 14350
rect 12728 14074 12756 15098
rect 12820 15026 12848 15098
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12728 13462 12756 14010
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12185 13084 12493 13093
rect 12185 13082 12191 13084
rect 12247 13082 12271 13084
rect 12327 13082 12351 13084
rect 12407 13082 12431 13084
rect 12487 13082 12493 13084
rect 12247 13030 12249 13082
rect 12429 13030 12431 13082
rect 12185 13028 12191 13030
rect 12247 13028 12271 13030
rect 12327 13028 12351 13030
rect 12407 13028 12431 13030
rect 12487 13028 12493 13030
rect 12185 13019 12493 13028
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 11624 11478 11744 11506
rect 11808 11512 11928 11540
rect 11624 11218 11652 11478
rect 11808 11370 11836 11512
rect 11716 11342 11836 11370
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11624 9518 11652 11154
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11428 9512 11480 9518
rect 11612 9512 11664 9518
rect 11428 9454 11480 9460
rect 11532 9472 11612 9500
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8634 11100 8910
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10980 8498 11100 8514
rect 10980 8492 11112 8498
rect 10980 8486 11060 8492
rect 11060 8434 11112 8440
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 8129 11008 8230
rect 10966 8120 11022 8129
rect 11072 8106 11100 8434
rect 11164 8265 11192 8978
rect 11242 8936 11298 8945
rect 11242 8871 11298 8880
rect 11256 8430 11284 8871
rect 11348 8566 11376 9114
rect 11440 9110 11468 9454
rect 11428 9104 11480 9110
rect 11428 9046 11480 9052
rect 11532 9042 11560 9472
rect 11612 9454 11664 9460
rect 11716 9178 11744 11342
rect 12084 11268 12112 12582
rect 12544 12374 12572 13262
rect 12912 12918 12940 17478
rect 13556 17202 13584 18906
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18154 13952 18566
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13740 17882 13768 18022
rect 13924 17882 13952 18090
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13740 17338 13768 17682
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13924 17202 13952 17818
rect 14016 17746 14044 18702
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 14200 17610 14228 18770
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14384 17746 14412 18566
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14188 17604 14240 17610
rect 14188 17546 14240 17552
rect 14200 17270 14228 17546
rect 14292 17338 14320 17682
rect 14476 17678 14504 18158
rect 14832 18148 14884 18154
rect 14884 18108 14964 18136
rect 14832 18090 14884 18096
rect 14542 17980 14850 17989
rect 14542 17978 14548 17980
rect 14604 17978 14628 17980
rect 14684 17978 14708 17980
rect 14764 17978 14788 17980
rect 14844 17978 14850 17980
rect 14604 17926 14606 17978
rect 14786 17926 14788 17978
rect 14542 17924 14548 17926
rect 14604 17924 14628 17926
rect 14684 17924 14708 17926
rect 14764 17924 14788 17926
rect 14844 17924 14850 17926
rect 14542 17915 14850 17924
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 13188 16046 13216 16458
rect 13924 16046 13952 16662
rect 14108 16658 14136 16934
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14016 16250 14044 16390
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13188 15706 13216 15846
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13556 15570 13584 15846
rect 14016 15706 14044 16186
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14108 15570 14136 15846
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 13004 14074 13032 15506
rect 13266 15464 13322 15473
rect 13266 15399 13322 15408
rect 13280 14822 13308 15399
rect 13556 15366 13584 15506
rect 14292 15366 14320 16390
rect 14476 15570 14504 17614
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14568 17338 14596 17478
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14936 17134 14964 18108
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15120 17338 15148 17682
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14542 16892 14850 16901
rect 14542 16890 14548 16892
rect 14604 16890 14628 16892
rect 14684 16890 14708 16892
rect 14764 16890 14788 16892
rect 14844 16890 14850 16892
rect 14604 16838 14606 16890
rect 14786 16838 14788 16890
rect 14542 16836 14548 16838
rect 14604 16836 14628 16838
rect 14684 16836 14708 16838
rect 14764 16836 14788 16838
rect 14844 16836 14850 16838
rect 14542 16827 14850 16836
rect 14924 16788 14976 16794
rect 14924 16730 14976 16736
rect 14648 16720 14700 16726
rect 14832 16720 14884 16726
rect 14700 16680 14832 16708
rect 14648 16662 14700 16668
rect 14832 16662 14884 16668
rect 14844 16454 14872 16662
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14542 15804 14850 15813
rect 14542 15802 14548 15804
rect 14604 15802 14628 15804
rect 14684 15802 14708 15804
rect 14764 15802 14788 15804
rect 14844 15802 14850 15804
rect 14604 15750 14606 15802
rect 14786 15750 14788 15802
rect 14542 15748 14548 15750
rect 14604 15748 14628 15750
rect 14684 15748 14708 15750
rect 14764 15748 14788 15750
rect 14844 15748 14850 15750
rect 14542 15739 14850 15748
rect 14936 15638 14964 16730
rect 15120 16658 15148 17138
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15028 16538 15056 16594
rect 15212 16538 15240 16934
rect 15028 16510 15240 16538
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 14924 15632 14976 15638
rect 14924 15574 14976 15580
rect 15120 15570 15148 16390
rect 15212 15978 15240 16510
rect 15304 16250 15332 18158
rect 15396 18154 15424 18906
rect 18510 18864 18566 18873
rect 18510 18799 18512 18808
rect 18564 18799 18566 18808
rect 18512 18770 18564 18776
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 16900 18524 17208 18533
rect 16900 18522 16906 18524
rect 16962 18522 16986 18524
rect 17042 18522 17066 18524
rect 17122 18522 17146 18524
rect 17202 18522 17208 18524
rect 16962 18470 16964 18522
rect 17144 18470 17146 18522
rect 16900 18468 16906 18470
rect 16962 18468 16986 18470
rect 17042 18468 17066 18470
rect 17122 18468 17146 18470
rect 17202 18468 17208 18470
rect 16900 18459 17208 18468
rect 19076 18465 19104 18566
rect 19062 18456 19118 18465
rect 19062 18391 19118 18400
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15396 17134 15424 18090
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16592 17746 16620 18022
rect 16304 17740 16356 17746
rect 16224 17700 16304 17728
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 15580 16726 15608 17274
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14292 15162 14320 15302
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14292 14958 14320 15098
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14476 14890 14504 15506
rect 15120 14958 15148 15506
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13280 14074 13308 14758
rect 13924 14482 13952 14826
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13004 13258 13032 14010
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13096 13274 13124 13330
rect 12992 13252 13044 13258
rect 13096 13246 13308 13274
rect 12992 13194 13044 13200
rect 13280 13172 13308 13246
rect 13360 13184 13412 13190
rect 13280 13144 13360 13172
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12808 12300 12860 12306
rect 12912 12288 12940 12718
rect 12992 12640 13044 12646
rect 12990 12608 12992 12617
rect 13044 12608 13046 12617
rect 12990 12543 13046 12552
rect 12860 12260 12940 12288
rect 12808 12242 12860 12248
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12185 11996 12493 12005
rect 12185 11994 12191 11996
rect 12247 11994 12271 11996
rect 12327 11994 12351 11996
rect 12407 11994 12431 11996
rect 12487 11994 12493 11996
rect 12247 11942 12249 11994
rect 12429 11942 12431 11994
rect 12185 11940 12191 11942
rect 12247 11940 12271 11942
rect 12327 11940 12351 11942
rect 12407 11940 12431 11942
rect 12487 11940 12493 11942
rect 12185 11931 12493 11940
rect 12544 11898 12572 12038
rect 12912 11898 12940 12260
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12530 11792 12586 11801
rect 12530 11727 12586 11736
rect 12544 11694 12572 11727
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 11900 11240 12112 11268
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11808 10810 11836 11154
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11808 9722 11836 10610
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11624 8634 11652 8978
rect 11612 8628 11664 8634
rect 11808 8616 11836 9386
rect 11900 9042 11928 11240
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10674 12112 10950
rect 12185 10908 12493 10917
rect 12185 10906 12191 10908
rect 12247 10906 12271 10908
rect 12327 10906 12351 10908
rect 12407 10906 12431 10908
rect 12487 10906 12493 10908
rect 12247 10854 12249 10906
rect 12429 10854 12431 10906
rect 12185 10852 12191 10854
rect 12247 10852 12271 10854
rect 12327 10852 12351 10854
rect 12407 10852 12431 10854
rect 12487 10852 12493 10854
rect 12185 10843 12493 10852
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11992 10062 12020 10474
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11992 9450 12020 9862
rect 11980 9444 12032 9450
rect 11980 9386 12032 9392
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11992 8634 12020 8978
rect 11612 8570 11664 8576
rect 11716 8588 11836 8616
rect 11980 8628 12032 8634
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11610 8528 11666 8537
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11150 8256 11206 8265
rect 11150 8191 11206 8200
rect 11072 8078 11192 8106
rect 10966 8055 11022 8064
rect 10980 7886 11008 8055
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10968 7880 11020 7886
rect 11072 7857 11100 7958
rect 10968 7822 11020 7828
rect 11058 7848 11114 7857
rect 10980 7342 11008 7822
rect 11058 7783 11114 7792
rect 11164 7750 11192 8078
rect 11348 8022 11376 8502
rect 11610 8463 11666 8472
rect 11624 8430 11652 8463
rect 11612 8424 11664 8430
rect 11426 8392 11482 8401
rect 11612 8366 11664 8372
rect 11426 8327 11482 8336
rect 11440 8294 11468 8327
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11716 8072 11744 8588
rect 11980 8570 12032 8576
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11440 8044 11744 8072
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11348 7546 11376 7754
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11256 7342 11284 7482
rect 10968 7336 11020 7342
rect 11244 7336 11296 7342
rect 10968 7278 11020 7284
rect 11150 7304 11206 7313
rect 10980 6866 11008 7278
rect 11244 7278 11296 7284
rect 11150 7239 11152 7248
rect 11204 7239 11206 7248
rect 11152 7210 11204 7216
rect 11164 7018 11192 7210
rect 11164 6990 11376 7018
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 6662 11284 6734
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 10966 6488 11022 6497
rect 10966 6423 11022 6432
rect 10980 6390 11008 6423
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10796 5250 10824 5306
rect 10796 5222 10916 5250
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10888 4706 10916 5222
rect 10980 4826 11008 5578
rect 11072 5166 11100 5646
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10966 4720 11022 4729
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10520 4282 10548 4626
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10704 3738 10732 4694
rect 10888 4678 10966 4706
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10796 4078 10824 4558
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 9827 2748 10135 2757
rect 9827 2746 9833 2748
rect 9889 2746 9913 2748
rect 9969 2746 9993 2748
rect 10049 2746 10073 2748
rect 10129 2746 10135 2748
rect 9889 2694 9891 2746
rect 10071 2694 10073 2746
rect 9827 2692 9833 2694
rect 9889 2692 9913 2694
rect 9969 2692 9993 2694
rect 10049 2692 10073 2694
rect 10129 2692 10135 2694
rect 9827 2683 10135 2692
rect 10598 2680 10654 2689
rect 10598 2615 10600 2624
rect 10652 2615 10654 2624
rect 10600 2586 10652 2592
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 9954 2544 10010 2553
rect 9680 2508 9732 2514
rect 9954 2479 10010 2488
rect 9680 2450 9732 2456
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9036 1964 9088 1970
rect 9036 1906 9088 1912
rect 8944 1828 8996 1834
rect 8944 1770 8996 1776
rect 9140 1562 9168 2246
rect 9600 1562 9628 2246
rect 9692 1902 9720 2450
rect 9968 2310 9996 2479
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10152 2038 10180 2246
rect 10244 2106 10272 2382
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 10140 2032 10192 2038
rect 10140 1974 10192 1980
rect 10796 1970 10824 4014
rect 10888 2514 10916 4678
rect 10966 4655 10968 4664
rect 11020 4655 11022 4664
rect 11060 4684 11112 4690
rect 10968 4626 11020 4632
rect 11060 4626 11112 4632
rect 11072 3942 11100 4626
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 10784 1964 10836 1970
rect 10784 1906 10836 1912
rect 9680 1896 9732 1902
rect 9680 1838 9732 1844
rect 10324 1828 10376 1834
rect 10324 1770 10376 1776
rect 9827 1660 10135 1669
rect 9827 1658 9833 1660
rect 9889 1658 9913 1660
rect 9969 1658 9993 1660
rect 10049 1658 10073 1660
rect 10129 1658 10135 1660
rect 9889 1606 9891 1658
rect 10071 1606 10073 1658
rect 9827 1604 9833 1606
rect 9889 1604 9913 1606
rect 9969 1604 9993 1606
rect 10049 1604 10073 1606
rect 10129 1604 10135 1606
rect 9827 1595 10135 1604
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 8760 1556 8812 1562
rect 8760 1498 8812 1504
rect 9128 1556 9180 1562
rect 9128 1498 9180 1504
rect 9588 1556 9640 1562
rect 9588 1498 9640 1504
rect 10336 1426 10364 1770
rect 10416 1760 10468 1766
rect 10416 1702 10468 1708
rect 10600 1760 10652 1766
rect 10600 1702 10652 1708
rect 10428 1562 10456 1702
rect 10416 1556 10468 1562
rect 10416 1498 10468 1504
rect 10612 1426 10640 1702
rect 11072 1562 11100 2450
rect 11060 1556 11112 1562
rect 11060 1498 11112 1504
rect 10324 1420 10376 1426
rect 10324 1362 10376 1368
rect 10600 1420 10652 1426
rect 10600 1362 10652 1368
rect 8392 1352 8444 1358
rect 8392 1294 8444 1300
rect 7470 1116 7778 1125
rect 7470 1114 7476 1116
rect 7532 1114 7556 1116
rect 7612 1114 7636 1116
rect 7692 1114 7716 1116
rect 7772 1114 7778 1116
rect 7532 1062 7534 1114
rect 7714 1062 7716 1114
rect 7470 1060 7476 1062
rect 7532 1060 7556 1062
rect 7612 1060 7636 1062
rect 7692 1060 7716 1062
rect 7772 1060 7778 1062
rect 7470 1051 7778 1060
rect 11164 1018 11192 6598
rect 11256 5098 11284 6598
rect 11348 5778 11376 6990
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11348 4978 11376 5238
rect 11256 4950 11376 4978
rect 11256 4690 11284 4950
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11348 3194 11376 4694
rect 11440 4690 11468 8044
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11716 7750 11744 7890
rect 11808 7886 11836 8366
rect 11900 7954 11928 8366
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11532 7342 11560 7686
rect 11716 7342 11744 7686
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11532 6798 11560 7278
rect 11716 6934 11744 7278
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11532 5778 11560 6258
rect 11808 6186 11836 7346
rect 11900 7342 11928 7890
rect 11992 7410 12020 8230
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11900 6798 11928 7278
rect 11992 6798 12020 7346
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11900 6254 11928 6734
rect 11992 6322 12020 6734
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11624 5658 11652 6122
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11532 5630 11652 5658
rect 11428 4684 11480 4690
rect 11532 4672 11560 5630
rect 11716 5166 11744 5850
rect 11808 5642 11836 6122
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11808 5098 11836 5578
rect 11796 5092 11848 5098
rect 11796 5034 11848 5040
rect 11612 4684 11664 4690
rect 11532 4644 11612 4672
rect 11428 4626 11480 4632
rect 11612 4626 11664 4632
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11520 4276 11572 4282
rect 11624 4264 11652 4422
rect 11572 4236 11652 4264
rect 11520 4218 11572 4224
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11348 2106 11376 2246
rect 11336 2100 11388 2106
rect 11336 2042 11388 2048
rect 11348 1562 11376 2042
rect 11428 1828 11480 1834
rect 11428 1770 11480 1776
rect 11440 1562 11468 1770
rect 11336 1556 11388 1562
rect 11336 1498 11388 1504
rect 11428 1556 11480 1562
rect 11428 1498 11480 1504
rect 11440 1426 11468 1498
rect 11244 1420 11296 1426
rect 11244 1362 11296 1368
rect 11428 1420 11480 1426
rect 11428 1362 11480 1368
rect 11256 1222 11284 1362
rect 11244 1216 11296 1222
rect 11244 1158 11296 1164
rect 7196 1012 7248 1018
rect 7196 954 7248 960
rect 11152 1012 11204 1018
rect 11152 954 11204 960
rect 11808 950 11836 5034
rect 11900 1018 11928 6190
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11992 5302 12020 5714
rect 12084 5302 12112 10202
rect 12176 9926 12204 10542
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12185 9820 12493 9829
rect 12185 9818 12191 9820
rect 12247 9818 12271 9820
rect 12327 9818 12351 9820
rect 12407 9818 12431 9820
rect 12487 9818 12493 9820
rect 12247 9766 12249 9818
rect 12429 9766 12431 9818
rect 12185 9764 12191 9766
rect 12247 9764 12271 9766
rect 12327 9764 12351 9766
rect 12407 9764 12431 9766
rect 12487 9764 12493 9766
rect 12185 9755 12493 9764
rect 12544 9704 12572 9862
rect 12452 9676 12572 9704
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12268 9024 12296 9454
rect 12452 9110 12480 9676
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12544 9178 12572 9522
rect 12636 9178 12664 10406
rect 12714 10024 12770 10033
rect 12714 9959 12770 9968
rect 12728 9518 12756 9959
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12348 9036 12400 9042
rect 12268 8996 12348 9024
rect 12348 8978 12400 8984
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12185 8732 12493 8741
rect 12185 8730 12191 8732
rect 12247 8730 12271 8732
rect 12327 8730 12351 8732
rect 12407 8730 12431 8732
rect 12487 8730 12493 8732
rect 12247 8678 12249 8730
rect 12429 8678 12431 8730
rect 12185 8676 12191 8678
rect 12247 8676 12271 8678
rect 12327 8676 12351 8678
rect 12407 8676 12431 8678
rect 12487 8676 12493 8678
rect 12185 8667 12493 8676
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12176 8294 12204 8434
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12162 8120 12218 8129
rect 12268 8106 12296 8366
rect 12218 8078 12296 8106
rect 12346 8120 12402 8129
rect 12162 8055 12218 8064
rect 12346 8055 12348 8064
rect 12400 8055 12402 8064
rect 12348 8026 12400 8032
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12176 7750 12204 7958
rect 12254 7848 12310 7857
rect 12254 7783 12256 7792
rect 12308 7783 12310 7792
rect 12256 7754 12308 7760
rect 12164 7744 12216 7750
rect 12452 7732 12480 7958
rect 12544 7800 12572 8366
rect 12636 8090 12664 8774
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12728 7818 12756 8978
rect 12820 8242 12848 11562
rect 13280 11234 13308 13144
rect 13360 13126 13412 13132
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13372 12434 13400 12854
rect 13556 12782 13584 13330
rect 13740 13172 13768 13670
rect 13832 13530 13860 13670
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13820 13388 13872 13394
rect 13872 13348 13952 13376
rect 13820 13330 13872 13336
rect 13820 13184 13872 13190
rect 13740 13144 13820 13172
rect 13820 13126 13872 13132
rect 13924 12986 13952 13348
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13832 12782 13860 12922
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13372 12406 13492 12434
rect 13280 11206 13400 11234
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13096 10713 13124 11086
rect 13372 11014 13400 11206
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13082 10704 13138 10713
rect 13082 10639 13138 10648
rect 12990 9480 13046 9489
rect 12990 9415 13046 9424
rect 12820 8214 12940 8242
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12716 7812 12768 7818
rect 12544 7772 12664 7800
rect 12452 7704 12572 7732
rect 12164 7686 12216 7692
rect 12185 7644 12493 7653
rect 12185 7642 12191 7644
rect 12247 7642 12271 7644
rect 12327 7642 12351 7644
rect 12407 7642 12431 7644
rect 12487 7642 12493 7644
rect 12247 7590 12249 7642
rect 12429 7590 12431 7642
rect 12185 7588 12191 7590
rect 12247 7588 12271 7590
rect 12327 7588 12351 7590
rect 12407 7588 12431 7590
rect 12487 7588 12493 7590
rect 12185 7579 12493 7588
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12452 6746 12480 7482
rect 12544 7410 12572 7704
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 6866 12572 7142
rect 12636 7002 12664 7772
rect 12716 7754 12768 7760
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12452 6718 12572 6746
rect 12185 6556 12493 6565
rect 12185 6554 12191 6556
rect 12247 6554 12271 6556
rect 12327 6554 12351 6556
rect 12407 6554 12431 6556
rect 12487 6554 12493 6556
rect 12247 6502 12249 6554
rect 12429 6502 12431 6554
rect 12185 6500 12191 6502
rect 12247 6500 12271 6502
rect 12327 6500 12351 6502
rect 12407 6500 12431 6502
rect 12487 6500 12493 6502
rect 12185 6491 12493 6500
rect 12544 6458 12572 6718
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12176 5846 12204 6394
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12452 5914 12480 6258
rect 12544 6066 12572 6394
rect 12636 6186 12664 6802
rect 12728 6798 12756 7482
rect 12820 7206 12848 7890
rect 12912 7478 12940 8214
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 13004 7410 13032 9415
rect 13464 9058 13492 12406
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11762 13676 12038
rect 13924 11898 13952 12582
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 9722 13768 11494
rect 13832 11218 13860 11562
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13832 9450 13860 9590
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13544 9104 13596 9110
rect 13464 9052 13544 9058
rect 13464 9046 13596 9052
rect 13268 9036 13320 9042
rect 13464 9030 13584 9046
rect 13268 8978 13320 8984
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13188 8548 13216 8842
rect 13280 8786 13308 8978
rect 13280 8758 13584 8786
rect 13188 8520 13400 8548
rect 13084 8492 13136 8498
rect 13136 8452 13216 8480
rect 13084 8434 13136 8440
rect 13082 8392 13138 8401
rect 13082 8327 13138 8336
rect 13096 8090 13124 8327
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 6866 12848 7142
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12544 6038 12664 6066
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12185 5468 12493 5477
rect 12185 5466 12191 5468
rect 12247 5466 12271 5468
rect 12327 5466 12351 5468
rect 12407 5466 12431 5468
rect 12487 5466 12493 5468
rect 12247 5414 12249 5466
rect 12429 5414 12431 5466
rect 12185 5412 12191 5414
rect 12247 5412 12271 5414
rect 12327 5412 12351 5414
rect 12407 5412 12431 5414
rect 12487 5412 12493 5414
rect 12185 5403 12493 5412
rect 12544 5352 12572 5850
rect 12452 5324 12572 5352
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 11992 5148 12020 5238
rect 12072 5160 12124 5166
rect 11992 5120 12072 5148
rect 12072 5102 12124 5108
rect 12452 5098 12480 5324
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11992 2038 12020 2246
rect 12084 2106 12112 4694
rect 12360 4690 12388 4762
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12185 4380 12493 4389
rect 12185 4378 12191 4380
rect 12247 4378 12271 4380
rect 12327 4378 12351 4380
rect 12407 4378 12431 4380
rect 12487 4378 12493 4380
rect 12247 4326 12249 4378
rect 12429 4326 12431 4378
rect 12185 4324 12191 4326
rect 12247 4324 12271 4326
rect 12327 4324 12351 4326
rect 12407 4324 12431 4326
rect 12487 4324 12493 4326
rect 12185 4315 12493 4324
rect 12544 4282 12572 5034
rect 12636 4758 12664 6038
rect 12624 4752 12676 4758
rect 12728 4729 12756 6734
rect 12806 6352 12862 6361
rect 12806 6287 12862 6296
rect 12820 6186 12848 6287
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12912 5098 12940 6802
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13004 5710 13032 6190
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12624 4694 12676 4700
rect 12714 4720 12770 4729
rect 12714 4655 12770 4664
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12185 3292 12493 3301
rect 12185 3290 12191 3292
rect 12247 3290 12271 3292
rect 12327 3290 12351 3292
rect 12407 3290 12431 3292
rect 12487 3290 12493 3292
rect 12247 3238 12249 3290
rect 12429 3238 12431 3290
rect 12185 3236 12191 3238
rect 12247 3236 12271 3238
rect 12327 3236 12351 3238
rect 12407 3236 12431 3238
rect 12487 3236 12493 3238
rect 12185 3227 12493 3236
rect 12544 3058 12572 4218
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12820 3194 12848 3946
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12544 2514 12572 2994
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12820 2774 12848 2926
rect 12728 2746 12848 2774
rect 12728 2514 12756 2746
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12185 2204 12493 2213
rect 12185 2202 12191 2204
rect 12247 2202 12271 2204
rect 12327 2202 12351 2204
rect 12407 2202 12431 2204
rect 12487 2202 12493 2204
rect 12247 2150 12249 2202
rect 12429 2150 12431 2202
rect 12185 2148 12191 2150
rect 12247 2148 12271 2150
rect 12327 2148 12351 2150
rect 12407 2148 12431 2150
rect 12487 2148 12493 2150
rect 12185 2139 12493 2148
rect 12728 2106 12756 2450
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 12716 2100 12768 2106
rect 12716 2042 12768 2048
rect 11980 2032 12032 2038
rect 11980 1974 12032 1980
rect 12164 1760 12216 1766
rect 12164 1702 12216 1708
rect 12176 1426 12204 1702
rect 12728 1562 12756 2042
rect 12716 1556 12768 1562
rect 12716 1498 12768 1504
rect 12164 1420 12216 1426
rect 12164 1362 12216 1368
rect 12185 1116 12493 1125
rect 12185 1114 12191 1116
rect 12247 1114 12271 1116
rect 12327 1114 12351 1116
rect 12407 1114 12431 1116
rect 12487 1114 12493 1116
rect 12247 1062 12249 1114
rect 12429 1062 12431 1114
rect 12185 1060 12191 1062
rect 12247 1060 12271 1062
rect 12327 1060 12351 1062
rect 12407 1060 12431 1062
rect 12487 1060 12493 1062
rect 12185 1051 12493 1060
rect 11888 1012 11940 1018
rect 11888 954 11940 960
rect 12912 950 12940 5034
rect 13004 4622 13032 5646
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13004 3602 13032 4558
rect 13096 4554 13124 7890
rect 13188 6662 13216 8452
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 7818 13308 8366
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13280 7313 13308 7346
rect 13266 7304 13322 7313
rect 13266 7239 13322 7248
rect 13280 6866 13308 7239
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13280 6118 13308 6598
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13372 5370 13400 8520
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13464 6322 13492 7822
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13096 3194 13124 3538
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13096 1902 13124 3130
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 13280 2106 13308 2858
rect 13556 2774 13584 8758
rect 13648 8537 13676 9318
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13634 8528 13690 8537
rect 13634 8463 13690 8472
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13648 6798 13676 8366
rect 13740 7546 13768 8910
rect 13832 8294 13860 8978
rect 13924 8294 13952 10746
rect 14016 9518 14044 14758
rect 14476 14482 14504 14826
rect 14542 14716 14850 14725
rect 14542 14714 14548 14716
rect 14604 14714 14628 14716
rect 14684 14714 14708 14716
rect 14764 14714 14788 14716
rect 14844 14714 14850 14716
rect 14604 14662 14606 14714
rect 14786 14662 14788 14714
rect 14542 14660 14548 14662
rect 14604 14660 14628 14662
rect 14684 14660 14708 14662
rect 14764 14660 14788 14662
rect 14844 14660 14850 14662
rect 14542 14651 14850 14660
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14292 13938 14320 14418
rect 14476 13938 14504 14418
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15028 14074 15056 14214
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14292 13530 14320 13874
rect 15212 13870 15240 14554
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 14542 13628 14850 13637
rect 14542 13626 14548 13628
rect 14604 13626 14628 13628
rect 14684 13626 14708 13628
rect 14764 13626 14788 13628
rect 14844 13626 14850 13628
rect 14604 13574 14606 13626
rect 14786 13574 14788 13626
rect 14542 13572 14548 13574
rect 14604 13572 14628 13574
rect 14684 13572 14708 13574
rect 14764 13572 14788 13574
rect 14844 13572 14850 13574
rect 14542 13563 14850 13572
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14200 12617 14228 13126
rect 14568 12918 14596 13126
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14830 12880 14886 12889
rect 14372 12844 14424 12850
rect 14830 12815 14886 12824
rect 14924 12844 14976 12850
rect 14372 12786 14424 12792
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14186 12608 14242 12617
rect 14186 12543 14242 12552
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14108 11762 14136 12242
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14108 11354 14136 11698
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14108 10266 14136 11086
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14094 9616 14150 9625
rect 14094 9551 14150 9560
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 8974 14044 9318
rect 14108 9178 14136 9551
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13832 7274 13860 8230
rect 14016 7954 14044 8298
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13924 7002 13952 7822
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7546 14044 7686
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6254 13676 6734
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 14002 6352 14058 6361
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13832 5302 13860 6326
rect 14002 6287 14058 6296
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13924 5914 13952 6190
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13832 5166 13860 5238
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13832 4078 13860 4966
rect 14016 4282 14044 6287
rect 14108 5370 14136 8978
rect 14200 8430 14228 12543
rect 14292 12374 14320 12718
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14292 11898 14320 12310
rect 14384 12170 14412 12786
rect 14844 12782 14872 12815
rect 14924 12786 14976 12792
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14372 12164 14424 12170
rect 14372 12106 14424 12112
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14384 11642 14412 12106
rect 14476 11801 14504 12718
rect 14542 12540 14850 12549
rect 14542 12538 14548 12540
rect 14604 12538 14628 12540
rect 14684 12538 14708 12540
rect 14764 12538 14788 12540
rect 14844 12538 14850 12540
rect 14604 12486 14606 12538
rect 14786 12486 14788 12538
rect 14542 12484 14548 12486
rect 14604 12484 14628 12486
rect 14684 12484 14708 12486
rect 14764 12484 14788 12486
rect 14844 12484 14850 12486
rect 14542 12475 14850 12484
rect 14462 11792 14518 11801
rect 14462 11727 14518 11736
rect 14292 11614 14412 11642
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14292 10810 14320 11614
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14280 9512 14332 9518
rect 14278 9480 14280 9489
rect 14332 9480 14334 9489
rect 14278 9415 14334 9424
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 9178 14320 9318
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14200 7546 14228 7890
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14200 5846 14228 7346
rect 14292 5914 14320 8910
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13556 2746 13676 2774
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 13084 1896 13136 1902
rect 13084 1838 13136 1844
rect 13176 1760 13228 1766
rect 13176 1702 13228 1708
rect 13188 1426 13216 1702
rect 13464 1426 13492 2518
rect 13648 1873 13676 2746
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 14016 2038 14044 2450
rect 14292 2310 14320 5714
rect 14384 5370 14412 11494
rect 14476 11286 14504 11630
rect 14936 11558 14964 12786
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14542 11452 14850 11461
rect 14542 11450 14548 11452
rect 14604 11450 14628 11452
rect 14684 11450 14708 11452
rect 14764 11450 14788 11452
rect 14844 11450 14850 11452
rect 14604 11398 14606 11450
rect 14786 11398 14788 11450
rect 14542 11396 14548 11398
rect 14604 11396 14628 11398
rect 14684 11396 14708 11398
rect 14764 11396 14788 11398
rect 14844 11396 14850 11398
rect 14542 11387 14850 11396
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14568 10810 14596 11154
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14556 10804 14608 10810
rect 14476 10764 14556 10792
rect 14476 10130 14504 10764
rect 14556 10746 14608 10752
rect 14542 10364 14850 10373
rect 14542 10362 14548 10364
rect 14604 10362 14628 10364
rect 14684 10362 14708 10364
rect 14764 10362 14788 10364
rect 14844 10362 14850 10364
rect 14604 10310 14606 10362
rect 14786 10310 14788 10362
rect 14542 10308 14548 10310
rect 14604 10308 14628 10310
rect 14684 10308 14708 10310
rect 14764 10308 14788 10310
rect 14844 10308 14850 10310
rect 14542 10299 14850 10308
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14476 9178 14504 9318
rect 14542 9276 14850 9285
rect 14542 9274 14548 9276
rect 14604 9274 14628 9276
rect 14684 9274 14708 9276
rect 14764 9274 14788 9276
rect 14844 9274 14850 9276
rect 14604 9222 14606 9274
rect 14786 9222 14788 9274
rect 14542 9220 14548 9222
rect 14604 9220 14628 9222
rect 14684 9220 14708 9222
rect 14764 9220 14788 9222
rect 14844 9220 14850 9222
rect 14542 9211 14850 9220
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14936 8430 14964 10950
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14476 7274 14504 8230
rect 14542 8188 14850 8197
rect 14542 8186 14548 8188
rect 14604 8186 14628 8188
rect 14684 8186 14708 8188
rect 14764 8186 14788 8188
rect 14844 8186 14850 8188
rect 14604 8134 14606 8186
rect 14786 8134 14788 8186
rect 14542 8132 14548 8134
rect 14604 8132 14628 8134
rect 14684 8132 14708 8134
rect 14764 8132 14788 8134
rect 14844 8132 14850 8134
rect 14542 8123 14850 8132
rect 14936 8090 14964 8230
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14922 7984 14978 7993
rect 14556 7948 14608 7954
rect 14922 7919 14924 7928
rect 14556 7890 14608 7896
rect 14976 7919 14978 7928
rect 14924 7890 14976 7896
rect 14568 7478 14596 7890
rect 15028 7886 15056 13806
rect 15212 13462 15240 13806
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 15120 11642 15148 12038
rect 15120 11614 15240 11642
rect 15212 11354 15240 11614
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15304 11098 15332 13670
rect 15488 11778 15516 14350
rect 15672 13870 15700 14418
rect 16132 14414 16160 17478
rect 16224 16017 16252 17700
rect 16304 17682 16356 17688
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16684 17610 16712 18022
rect 18064 17814 18092 18158
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 18248 17882 18276 18090
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16210 16008 16266 16017
rect 16210 15943 16266 15952
rect 16224 14482 16252 15943
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15764 12306 15792 12582
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15212 11070 15332 11098
rect 15396 11750 15516 11778
rect 15672 11762 15700 12038
rect 15764 11762 15792 12038
rect 15660 11756 15712 11762
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15120 10130 15148 10542
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15120 8090 15148 9862
rect 15212 9110 15240 11070
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15304 10742 15332 10950
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15304 9450 15332 10678
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15290 9072 15346 9081
rect 15290 9007 15292 9016
rect 15344 9007 15346 9016
rect 15292 8978 15344 8984
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15016 7880 15068 7886
rect 15068 7840 15148 7868
rect 15016 7822 15068 7828
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14924 7472 14976 7478
rect 14924 7414 14976 7420
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 14476 6866 14504 7210
rect 14542 7100 14850 7109
rect 14542 7098 14548 7100
rect 14604 7098 14628 7100
rect 14684 7098 14708 7100
rect 14764 7098 14788 7100
rect 14844 7098 14850 7100
rect 14604 7046 14606 7098
rect 14786 7046 14788 7098
rect 14542 7044 14548 7046
rect 14604 7044 14628 7046
rect 14684 7044 14708 7046
rect 14764 7044 14788 7046
rect 14844 7044 14850 7046
rect 14542 7035 14850 7044
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14462 6352 14518 6361
rect 14462 6287 14518 6296
rect 14476 6254 14504 6287
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5370 14504 6054
rect 14542 6012 14850 6021
rect 14542 6010 14548 6012
rect 14604 6010 14628 6012
rect 14684 6010 14708 6012
rect 14764 6010 14788 6012
rect 14844 6010 14850 6012
rect 14604 5958 14606 6010
rect 14786 5958 14788 6010
rect 14542 5956 14548 5958
rect 14604 5956 14628 5958
rect 14684 5956 14708 5958
rect 14764 5956 14788 5958
rect 14844 5956 14850 5958
rect 14542 5947 14850 5956
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14752 5166 14780 5782
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14384 4826 14412 5102
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14384 3602 14412 3946
rect 14476 3738 14504 4966
rect 14542 4924 14850 4933
rect 14542 4922 14548 4924
rect 14604 4922 14628 4924
rect 14684 4922 14708 4924
rect 14764 4922 14788 4924
rect 14844 4922 14850 4924
rect 14604 4870 14606 4922
rect 14786 4870 14788 4922
rect 14542 4868 14548 4870
rect 14604 4868 14628 4870
rect 14684 4868 14708 4870
rect 14764 4868 14788 4870
rect 14844 4868 14850 4870
rect 14542 4859 14850 4868
rect 14542 3836 14850 3845
rect 14542 3834 14548 3836
rect 14604 3834 14628 3836
rect 14684 3834 14708 3836
rect 14764 3834 14788 3836
rect 14844 3834 14850 3836
rect 14604 3782 14606 3834
rect 14786 3782 14788 3834
rect 14542 3780 14548 3782
rect 14604 3780 14628 3782
rect 14684 3780 14708 3782
rect 14764 3780 14788 3782
rect 14844 3780 14850 3782
rect 14542 3771 14850 3780
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14542 2748 14850 2757
rect 14542 2746 14548 2748
rect 14604 2746 14628 2748
rect 14684 2746 14708 2748
rect 14764 2746 14788 2748
rect 14844 2746 14850 2748
rect 14604 2694 14606 2746
rect 14786 2694 14788 2746
rect 14542 2692 14548 2694
rect 14604 2692 14628 2694
rect 14684 2692 14708 2694
rect 14764 2692 14788 2694
rect 14844 2692 14850 2694
rect 14542 2683 14850 2692
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14004 2032 14056 2038
rect 14004 1974 14056 1980
rect 14188 1896 14240 1902
rect 13634 1864 13690 1873
rect 14188 1838 14240 1844
rect 13634 1799 13690 1808
rect 13912 1760 13964 1766
rect 13912 1702 13964 1708
rect 13924 1494 13952 1702
rect 14200 1562 14228 1838
rect 14542 1660 14850 1669
rect 14542 1658 14548 1660
rect 14604 1658 14628 1660
rect 14684 1658 14708 1660
rect 14764 1658 14788 1660
rect 14844 1658 14850 1660
rect 14604 1606 14606 1658
rect 14786 1606 14788 1658
rect 14542 1604 14548 1606
rect 14604 1604 14628 1606
rect 14684 1604 14708 1606
rect 14764 1604 14788 1606
rect 14844 1604 14850 1606
rect 14542 1595 14850 1604
rect 14936 1562 14964 7414
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15028 5914 15056 6598
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 15120 5778 15148 7840
rect 15212 7546 15240 8366
rect 15290 7984 15346 7993
rect 15290 7919 15346 7928
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15212 6118 15240 6802
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15212 5234 15240 6054
rect 15304 5846 15332 7919
rect 15396 7750 15424 11750
rect 15660 11698 15712 11704
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15488 11218 15516 11630
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15580 10538 15608 11222
rect 15672 11014 15700 11698
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15856 10130 15884 12038
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15856 8974 15884 10066
rect 15948 9382 15976 14282
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 13394 16068 13670
rect 16132 13530 16160 14214
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16224 13530 16252 13738
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16040 12374 16068 13330
rect 16224 12714 16252 13466
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16028 12368 16080 12374
rect 16028 12310 16080 12316
rect 16040 11898 16068 12310
rect 16224 12238 16252 12650
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16316 11778 16344 17546
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 16776 17338 16804 17478
rect 16900 17436 17208 17445
rect 16900 17434 16906 17436
rect 16962 17434 16986 17436
rect 17042 17434 17066 17436
rect 17122 17434 17146 17436
rect 17202 17434 17208 17436
rect 16962 17382 16964 17434
rect 17144 17382 17146 17434
rect 16900 17380 16906 17382
rect 16962 17380 16986 17382
rect 17042 17380 17066 17382
rect 17122 17380 17146 17382
rect 17202 17380 17208 17382
rect 16900 17371 17208 17380
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16776 17134 16804 17274
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16684 16794 16712 16934
rect 16960 16794 16988 16934
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 17236 16590 17264 17478
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17328 16522 17356 17002
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 16900 16348 17208 16357
rect 16900 16346 16906 16348
rect 16962 16346 16986 16348
rect 17042 16346 17066 16348
rect 17122 16346 17146 16348
rect 17202 16346 17208 16348
rect 16962 16294 16964 16346
rect 17144 16294 17146 16346
rect 16900 16292 16906 16294
rect 16962 16292 16986 16294
rect 17042 16292 17066 16294
rect 17122 16292 17146 16294
rect 17202 16292 17208 16294
rect 16900 16283 17208 16292
rect 17236 16046 17264 16390
rect 17512 16250 17540 16594
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17328 15706 17356 15846
rect 17512 15706 17540 16186
rect 17788 16182 17816 17070
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17880 16658 17908 16934
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17880 16250 17908 16594
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17776 16176 17828 16182
rect 17776 16118 17828 16124
rect 17788 16046 17816 16118
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16132 11750 16344 11778
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15948 9058 15976 9318
rect 15948 9030 16068 9058
rect 15844 8968 15896 8974
rect 15936 8968 15988 8974
rect 15844 8910 15896 8916
rect 15934 8936 15936 8945
rect 15988 8936 15990 8945
rect 15934 8871 15990 8880
rect 16040 8566 16068 9030
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15488 6390 15516 8434
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15580 7954 15608 8298
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15660 7948 15712 7954
rect 15712 7908 15976 7936
rect 15660 7890 15712 7896
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15580 6322 15608 7890
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15856 7410 15884 7754
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15856 6474 15884 7346
rect 15764 6458 15884 6474
rect 15752 6452 15884 6458
rect 15804 6446 15884 6452
rect 15752 6394 15804 6400
rect 15764 6338 15792 6394
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15672 6310 15792 6338
rect 15568 6180 15620 6186
rect 15568 6122 15620 6128
rect 15580 5914 15608 6122
rect 15672 5914 15700 6310
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15764 5914 15792 6190
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15292 5840 15344 5846
rect 15856 5817 15884 6190
rect 15292 5782 15344 5788
rect 15842 5808 15898 5817
rect 15660 5772 15712 5778
rect 15842 5743 15898 5752
rect 15660 5714 15712 5720
rect 15290 5672 15346 5681
rect 15290 5607 15346 5616
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15304 5166 15332 5607
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15396 5166 15424 5510
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15396 4146 15424 4626
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15106 3768 15162 3777
rect 15106 3703 15108 3712
rect 15160 3703 15162 3712
rect 15108 3674 15160 3680
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15120 3194 15148 3538
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15212 2122 15240 4014
rect 15396 3738 15424 4082
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15304 3194 15332 3470
rect 15396 3466 15424 3674
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15304 2854 15332 3130
rect 15580 3126 15608 4082
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15304 2650 15332 2790
rect 15672 2650 15700 5714
rect 15948 4282 15976 7908
rect 16040 4826 16068 8366
rect 16132 6322 16160 11750
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11218 16252 11494
rect 16316 11354 16344 11630
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16408 11234 16436 14758
rect 16500 13870 16528 14758
rect 16592 14482 16620 15302
rect 16900 15260 17208 15269
rect 16900 15258 16906 15260
rect 16962 15258 16986 15260
rect 17042 15258 17066 15260
rect 17122 15258 17146 15260
rect 17202 15258 17208 15260
rect 16962 15206 16964 15258
rect 17144 15206 17146 15258
rect 16900 15204 16906 15206
rect 16962 15204 16986 15206
rect 17042 15204 17066 15206
rect 17122 15204 17146 15206
rect 17202 15204 17208 15206
rect 16900 15195 17208 15204
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16900 14172 17208 14181
rect 16900 14170 16906 14172
rect 16962 14170 16986 14172
rect 17042 14170 17066 14172
rect 17122 14170 17146 14172
rect 17202 14170 17208 14172
rect 16962 14118 16964 14170
rect 17144 14118 17146 14170
rect 16900 14116 16906 14118
rect 16962 14116 16986 14118
rect 17042 14116 17066 14118
rect 17122 14116 17146 14118
rect 17202 14116 17208 14118
rect 16900 14107 17208 14116
rect 17420 14074 17448 15302
rect 17512 15194 17540 15642
rect 17880 15366 17908 15982
rect 17972 15910 18000 17070
rect 18064 16726 18092 17750
rect 18248 16998 18276 17818
rect 19076 17785 19104 18158
rect 19257 17980 19565 17989
rect 19257 17978 19263 17980
rect 19319 17978 19343 17980
rect 19399 17978 19423 17980
rect 19479 17978 19503 17980
rect 19559 17978 19565 17980
rect 19319 17926 19321 17978
rect 19501 17926 19503 17978
rect 19257 17924 19263 17926
rect 19319 17924 19343 17926
rect 19399 17924 19423 17926
rect 19479 17924 19503 17926
rect 19559 17924 19565 17926
rect 19257 17915 19565 17924
rect 19062 17776 19118 17785
rect 18788 17740 18840 17746
rect 19062 17711 19118 17720
rect 18788 17682 18840 17688
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18708 17338 18736 17478
rect 18800 17338 18828 17682
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 19062 17096 19118 17105
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18248 16794 18276 16934
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 18064 15194 18092 16662
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18420 16176 18472 16182
rect 18420 16118 18472 16124
rect 18432 15706 18460 16118
rect 18616 15910 18644 16594
rect 18708 16454 18736 17070
rect 19062 17031 19118 17040
rect 19076 16658 19104 17031
rect 19257 16892 19565 16901
rect 19257 16890 19263 16892
rect 19319 16890 19343 16892
rect 19399 16890 19423 16892
rect 19479 16890 19503 16892
rect 19559 16890 19565 16892
rect 19319 16838 19321 16890
rect 19501 16838 19503 16890
rect 19257 16836 19263 16838
rect 19319 16836 19343 16838
rect 19399 16836 19423 16838
rect 19479 16836 19503 16838
rect 19559 16836 19565 16838
rect 19257 16827 19565 16836
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 19257 15804 19565 15813
rect 19257 15802 19263 15804
rect 19319 15802 19343 15804
rect 19399 15802 19423 15804
rect 19479 15802 19503 15804
rect 19559 15802 19565 15804
rect 19319 15750 19321 15802
rect 19501 15750 19503 15802
rect 19257 15748 19263 15750
rect 19319 15748 19343 15750
rect 19399 15748 19423 15750
rect 19479 15748 19503 15750
rect 19559 15748 19565 15750
rect 19257 15739 19565 15748
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18236 15632 18288 15638
rect 18236 15574 18288 15580
rect 17512 15166 17632 15194
rect 17604 14958 17632 15166
rect 17788 15166 18092 15194
rect 17788 14958 17816 15166
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17788 13870 17816 14894
rect 18248 14822 18276 15574
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16500 11694 16528 13126
rect 16592 12345 16620 13670
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 16900 13084 17208 13093
rect 16900 13082 16906 13084
rect 16962 13082 16986 13084
rect 17042 13082 17066 13084
rect 17122 13082 17146 13084
rect 17202 13082 17208 13084
rect 16962 13030 16964 13082
rect 17144 13030 17146 13082
rect 16900 13028 16906 13030
rect 16962 13028 16986 13030
rect 17042 13028 17066 13030
rect 17122 13028 17146 13030
rect 17202 13028 17208 13030
rect 16900 13019 17208 13028
rect 17236 12782 17264 13398
rect 17788 13326 17816 13806
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17590 13016 17646 13025
rect 17590 12951 17592 12960
rect 17644 12951 17646 12960
rect 17592 12922 17644 12928
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17590 12744 17646 12753
rect 17590 12679 17646 12688
rect 17604 12442 17632 12679
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 16578 12336 16634 12345
rect 16578 12271 16634 12280
rect 17314 12336 17370 12345
rect 17314 12271 17316 12280
rect 17368 12271 17370 12280
rect 17316 12242 17368 12248
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16316 11206 16436 11234
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 9178 16252 10406
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16316 8430 16344 11206
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10062 16436 10406
rect 16592 10146 16620 12174
rect 16900 11996 17208 12005
rect 16900 11994 16906 11996
rect 16962 11994 16986 11996
rect 17042 11994 17066 11996
rect 17122 11994 17146 11996
rect 17202 11994 17208 11996
rect 16962 11942 16964 11994
rect 17144 11942 17146 11994
rect 16900 11940 16906 11942
rect 16962 11940 16986 11942
rect 17042 11940 17066 11942
rect 17122 11940 17146 11942
rect 17202 11940 17208 11942
rect 16900 11931 17208 11940
rect 18156 11642 18184 13670
rect 18340 12986 18368 15302
rect 18708 15162 18736 15506
rect 18892 15162 18920 15506
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18432 12782 18460 14486
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18524 13870 18552 14214
rect 18616 13870 18644 14826
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18708 14482 18736 14758
rect 18892 14634 18920 15098
rect 18972 14952 19024 14958
rect 18972 14894 19024 14900
rect 18800 14606 18920 14634
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18432 11898 18460 12718
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18616 11694 18644 13330
rect 18708 12986 18736 14418
rect 18800 13802 18828 14606
rect 18984 14550 19012 14894
rect 19257 14716 19565 14725
rect 19257 14714 19263 14716
rect 19319 14714 19343 14716
rect 19399 14714 19423 14716
rect 19479 14714 19503 14716
rect 19559 14714 19565 14716
rect 19319 14662 19321 14714
rect 19501 14662 19503 14714
rect 19257 14660 19263 14662
rect 19319 14660 19343 14662
rect 19399 14660 19423 14662
rect 19479 14660 19503 14662
rect 19559 14660 19565 14662
rect 19257 14651 19565 14660
rect 18972 14544 19024 14550
rect 18972 14486 19024 14492
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 18892 14074 18920 14418
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18892 12782 18920 14010
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18880 12776 18932 12782
rect 18800 12736 18880 12764
rect 18800 12322 18828 12736
rect 18880 12718 18932 12724
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18708 12306 18828 12322
rect 18892 12306 18920 12582
rect 18696 12300 18828 12306
rect 18748 12294 18828 12300
rect 18696 12242 18748 12248
rect 18800 11898 18828 12294
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18420 11688 18472 11694
rect 18156 11614 18276 11642
rect 18604 11688 18656 11694
rect 18472 11636 18552 11642
rect 18420 11630 18552 11636
rect 18604 11630 18656 11636
rect 18432 11614 18552 11630
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 17696 11218 17724 11494
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 16900 10908 17208 10917
rect 16900 10906 16906 10908
rect 16962 10906 16986 10908
rect 17042 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17208 10908
rect 16962 10854 16964 10906
rect 17144 10854 17146 10906
rect 16900 10852 16906 10854
rect 16962 10852 16986 10854
rect 17042 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17208 10854
rect 16900 10843 17208 10852
rect 16670 10568 16726 10577
rect 17696 10538 17724 11154
rect 16670 10503 16726 10512
rect 17684 10532 17736 10538
rect 16500 10118 16620 10146
rect 16684 10130 16712 10503
rect 17684 10474 17736 10480
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16672 10124 16724 10130
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16224 6934 16252 7890
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16316 7546 16344 7822
rect 16408 7750 16436 8230
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16316 5778 16344 7278
rect 16500 6458 16528 10118
rect 16672 10066 16724 10072
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 8090 16620 9998
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16684 9042 16712 9522
rect 16776 9450 16804 10406
rect 17316 10056 17368 10062
rect 17314 10024 17316 10033
rect 17368 10024 17370 10033
rect 17314 9959 17370 9968
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 16900 9820 17208 9829
rect 16900 9818 16906 9820
rect 16962 9818 16986 9820
rect 17042 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17208 9820
rect 16962 9766 16964 9818
rect 17144 9766 17146 9818
rect 16900 9764 16906 9766
rect 16962 9764 16986 9766
rect 17042 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17208 9766
rect 16900 9755 17208 9764
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16764 9444 16816 9450
rect 16764 9386 16816 9392
rect 17052 9110 17080 9454
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16684 8498 16712 8978
rect 16900 8732 17208 8741
rect 16900 8730 16906 8732
rect 16962 8730 16986 8732
rect 17042 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17208 8732
rect 16962 8678 16964 8730
rect 17144 8678 17146 8730
rect 16900 8676 16906 8678
rect 16962 8676 16986 8678
rect 17042 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17208 8678
rect 16900 8667 17208 8676
rect 17328 8566 17356 9046
rect 17512 8634 17540 9862
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17788 8634 17816 9658
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16684 6866 16712 8298
rect 17328 8022 17356 8502
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17696 7954 17724 8434
rect 17880 8430 17908 8978
rect 17972 8498 18000 11154
rect 18156 11014 18184 11494
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18248 10810 18276 11614
rect 18524 11558 18552 11614
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18248 10198 18276 10746
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17880 7993 17908 8366
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 17866 7984 17922 7993
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17684 7948 17736 7954
rect 17866 7919 17922 7928
rect 17684 7890 17736 7896
rect 16900 7644 17208 7653
rect 16900 7642 16906 7644
rect 16962 7642 16986 7644
rect 17042 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17208 7644
rect 16962 7590 16964 7642
rect 17144 7590 17146 7642
rect 16900 7588 16906 7590
rect 16962 7588 16986 7590
rect 17042 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17208 7590
rect 16900 7579 17208 7588
rect 17236 7342 17264 7890
rect 17696 7342 17724 7890
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16900 6556 17208 6565
rect 16900 6554 16906 6556
rect 16962 6554 16986 6556
rect 17042 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17208 6556
rect 16962 6502 16964 6554
rect 17144 6502 17146 6554
rect 16900 6500 16906 6502
rect 16962 6500 16986 6502
rect 17042 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17208 6502
rect 16900 6491 17208 6500
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 17236 6254 17264 7278
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17512 6905 17540 6938
rect 17498 6896 17554 6905
rect 17880 6882 17908 7278
rect 17498 6831 17554 6840
rect 17788 6854 17908 6882
rect 17788 6254 17816 6854
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 16132 5234 16160 5510
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16316 5098 16344 5714
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16500 4690 16528 5714
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15764 3194 15792 3334
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15844 3120 15896 3126
rect 15844 3062 15896 3068
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 15212 2094 15332 2122
rect 15672 2106 15700 2450
rect 15752 2304 15804 2310
rect 15856 2292 15884 3062
rect 15948 2854 15976 3470
rect 16132 3466 16160 4014
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16132 3194 16160 3402
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16316 3058 16344 3674
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 16040 2774 16068 2858
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16040 2746 16160 2774
rect 16132 2514 16160 2746
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 15936 2304 15988 2310
rect 15856 2264 15936 2292
rect 15752 2246 15804 2252
rect 15936 2246 15988 2252
rect 15304 1902 15332 2094
rect 15660 2100 15712 2106
rect 15660 2042 15712 2048
rect 15016 1896 15068 1902
rect 15016 1838 15068 1844
rect 15292 1896 15344 1902
rect 15292 1838 15344 1844
rect 14188 1556 14240 1562
rect 14188 1498 14240 1504
rect 14924 1556 14976 1562
rect 14924 1498 14976 1504
rect 13912 1488 13964 1494
rect 13912 1430 13964 1436
rect 13176 1420 13228 1426
rect 13176 1362 13228 1368
rect 13452 1420 13504 1426
rect 13452 1362 13504 1368
rect 13544 1420 13596 1426
rect 13544 1362 13596 1368
rect 13176 1284 13228 1290
rect 13176 1226 13228 1232
rect 11796 944 11848 950
rect 11796 886 11848 892
rect 12900 944 12952 950
rect 12900 886 12952 892
rect 13188 814 13216 1226
rect 13556 1018 13584 1362
rect 13924 1018 13952 1430
rect 14200 1018 14228 1498
rect 15028 1494 15056 1838
rect 15764 1834 15792 2246
rect 15200 1828 15252 1834
rect 15200 1770 15252 1776
rect 15752 1828 15804 1834
rect 15752 1770 15804 1776
rect 15212 1562 15240 1770
rect 15660 1760 15712 1766
rect 15660 1702 15712 1708
rect 15200 1556 15252 1562
rect 15200 1498 15252 1504
rect 15016 1488 15068 1494
rect 15016 1430 15068 1436
rect 15672 1426 15700 1702
rect 15660 1420 15712 1426
rect 15660 1362 15712 1368
rect 14464 1216 14516 1222
rect 14464 1158 14516 1164
rect 14476 1018 14504 1158
rect 15948 1018 15976 2246
rect 16132 1562 16160 2450
rect 16408 2378 16436 2790
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 16304 1828 16356 1834
rect 16304 1770 16356 1776
rect 16212 1760 16264 1766
rect 16212 1702 16264 1708
rect 16224 1562 16252 1702
rect 16120 1556 16172 1562
rect 16120 1498 16172 1504
rect 16212 1556 16264 1562
rect 16212 1498 16264 1504
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 13544 1012 13596 1018
rect 13544 954 13596 960
rect 13912 1012 13964 1018
rect 13912 954 13964 960
rect 14188 1012 14240 1018
rect 14188 954 14240 960
rect 14464 1012 14516 1018
rect 14464 954 14516 960
rect 15936 1012 15988 1018
rect 15936 954 15988 960
rect 16132 814 16160 1294
rect 16316 1018 16344 1770
rect 16408 1426 16436 2314
rect 16500 1986 16528 2926
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16592 2650 16620 2790
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16684 2106 16712 6190
rect 17236 5846 17264 6190
rect 17788 5914 17816 6190
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 16900 5468 17208 5477
rect 16900 5466 16906 5468
rect 16962 5466 16986 5468
rect 17042 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17208 5468
rect 16962 5414 16964 5466
rect 17144 5414 17146 5466
rect 16900 5412 16906 5414
rect 16962 5412 16986 5414
rect 17042 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17208 5414
rect 16900 5403 17208 5412
rect 17420 5098 17448 5714
rect 17408 5092 17460 5098
rect 17408 5034 17460 5040
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16776 4826 16804 4966
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 17420 4758 17448 5034
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16776 4214 16804 4422
rect 16900 4380 17208 4389
rect 16900 4378 16906 4380
rect 16962 4378 16986 4380
rect 17042 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17208 4380
rect 16962 4326 16964 4378
rect 17144 4326 17146 4378
rect 16900 4324 16906 4326
rect 16962 4324 16986 4326
rect 17042 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17208 4326
rect 16900 4315 17208 4324
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16762 3768 16818 3777
rect 16960 3738 16988 4014
rect 16762 3703 16764 3712
rect 16816 3703 16818 3712
rect 16948 3732 17000 3738
rect 16764 3674 16816 3680
rect 16948 3674 17000 3680
rect 16960 3380 16988 3674
rect 16776 3352 16988 3380
rect 16776 2990 16804 3352
rect 16900 3292 17208 3301
rect 16900 3290 16906 3292
rect 16962 3290 16986 3292
rect 17042 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17208 3292
rect 16962 3238 16964 3290
rect 17144 3238 17146 3290
rect 16900 3236 16906 3238
rect 16962 3236 16986 3238
rect 17042 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17208 3238
rect 16900 3227 17208 3236
rect 17236 3194 17264 4218
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17328 3398 17356 4014
rect 17512 3738 17540 5850
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17880 3670 17908 3878
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 17328 2650 17356 3334
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17788 2582 17816 2858
rect 17880 2650 17908 3606
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 16900 2204 17208 2213
rect 16900 2202 16906 2204
rect 16962 2202 16986 2204
rect 17042 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17208 2204
rect 16962 2150 16964 2202
rect 17144 2150 17146 2202
rect 16900 2148 16906 2150
rect 16962 2148 16986 2150
rect 17042 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17208 2150
rect 16900 2139 17208 2148
rect 17972 2106 18000 8298
rect 18064 7818 18092 8298
rect 18052 7812 18104 7818
rect 18052 7754 18104 7760
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 18064 5166 18092 6870
rect 18156 6458 18184 8434
rect 18248 8430 18276 9318
rect 18524 9194 18552 11494
rect 18616 11150 18644 11630
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18708 10606 18736 10950
rect 18892 10606 18920 12242
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18800 9586 18828 10474
rect 18892 10130 18920 10542
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18984 9722 19012 13670
rect 19257 13628 19565 13637
rect 19257 13626 19263 13628
rect 19319 13626 19343 13628
rect 19399 13626 19423 13628
rect 19479 13626 19503 13628
rect 19559 13626 19565 13628
rect 19319 13574 19321 13626
rect 19501 13574 19503 13626
rect 19257 13572 19263 13574
rect 19319 13572 19343 13574
rect 19399 13572 19423 13574
rect 19479 13572 19503 13574
rect 19559 13572 19565 13574
rect 19257 13563 19565 13572
rect 19257 12540 19565 12549
rect 19257 12538 19263 12540
rect 19319 12538 19343 12540
rect 19399 12538 19423 12540
rect 19479 12538 19503 12540
rect 19559 12538 19565 12540
rect 19319 12486 19321 12538
rect 19501 12486 19503 12538
rect 19257 12484 19263 12486
rect 19319 12484 19343 12486
rect 19399 12484 19423 12486
rect 19479 12484 19503 12486
rect 19559 12484 19565 12486
rect 19257 12475 19565 12484
rect 19062 11656 19118 11665
rect 19062 11591 19118 11600
rect 19076 11218 19104 11591
rect 19257 11452 19565 11461
rect 19257 11450 19263 11452
rect 19319 11450 19343 11452
rect 19399 11450 19423 11452
rect 19479 11450 19503 11452
rect 19559 11450 19565 11452
rect 19319 11398 19321 11450
rect 19501 11398 19503 11450
rect 19257 11396 19263 11398
rect 19319 11396 19343 11398
rect 19399 11396 19423 11398
rect 19479 11396 19503 11398
rect 19559 11396 19565 11398
rect 19257 11387 19565 11396
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 19257 10364 19565 10373
rect 19257 10362 19263 10364
rect 19319 10362 19343 10364
rect 19399 10362 19423 10364
rect 19479 10362 19503 10364
rect 19559 10362 19565 10364
rect 19319 10310 19321 10362
rect 19501 10310 19503 10362
rect 19257 10308 19263 10310
rect 19319 10308 19343 10310
rect 19399 10308 19423 10310
rect 19479 10308 19503 10310
rect 19559 10308 19565 10310
rect 19257 10299 19565 10308
rect 18972 9716 19024 9722
rect 18892 9676 18972 9704
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18524 9178 18644 9194
rect 18512 9172 18644 9178
rect 18564 9166 18644 9172
rect 18512 9114 18564 9120
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18432 6338 18460 8978
rect 18524 8362 18552 8978
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18616 7970 18644 9166
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8294 18736 8774
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18524 7954 18644 7970
rect 18512 7948 18644 7954
rect 18564 7942 18644 7948
rect 18512 7890 18564 7896
rect 18524 7546 18552 7890
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18708 7410 18736 8230
rect 18892 7546 18920 9676
rect 18972 9658 19024 9664
rect 19257 9276 19565 9285
rect 19257 9274 19263 9276
rect 19319 9274 19343 9276
rect 19399 9274 19423 9276
rect 19479 9274 19503 9276
rect 19559 9274 19565 9276
rect 19319 9222 19321 9274
rect 19501 9222 19503 9274
rect 19257 9220 19263 9222
rect 19319 9220 19343 9222
rect 19399 9220 19423 9222
rect 19479 9220 19503 9222
rect 19559 9220 19565 9222
rect 19257 9211 19565 9220
rect 19257 8188 19565 8197
rect 19257 8186 19263 8188
rect 19319 8186 19343 8188
rect 19399 8186 19423 8188
rect 19479 8186 19503 8188
rect 19559 8186 19565 8188
rect 19319 8134 19321 8186
rect 19501 8134 19503 8186
rect 19257 8132 19263 8134
rect 19319 8132 19343 8134
rect 19399 8132 19423 8134
rect 19479 8132 19503 8134
rect 19559 8132 19565 8134
rect 19257 8123 19565 8132
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18616 6866 18644 7142
rect 18984 6866 19012 7958
rect 19257 7100 19565 7109
rect 19257 7098 19263 7100
rect 19319 7098 19343 7100
rect 19399 7098 19423 7100
rect 19479 7098 19503 7100
rect 19559 7098 19565 7100
rect 19319 7046 19321 7098
rect 19501 7046 19503 7098
rect 19257 7044 19263 7046
rect 19319 7044 19343 7046
rect 19399 7044 19423 7046
rect 19479 7044 19503 7046
rect 19559 7044 19565 7046
rect 19257 7035 19565 7044
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 18248 6310 18460 6338
rect 18616 6322 18644 6802
rect 18604 6316 18656 6322
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18064 4690 18092 5102
rect 18156 5030 18184 5714
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18156 4010 18184 4966
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 16672 2100 16724 2106
rect 16672 2042 16724 2048
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 16500 1958 16620 1986
rect 16488 1896 16540 1902
rect 16488 1838 16540 1844
rect 16500 1426 16528 1838
rect 16592 1834 16620 1958
rect 16580 1828 16632 1834
rect 16580 1770 16632 1776
rect 18248 1562 18276 6310
rect 18604 6258 18656 6264
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18340 5914 18368 6190
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18432 5794 18460 6190
rect 19257 6012 19565 6021
rect 19257 6010 19263 6012
rect 19319 6010 19343 6012
rect 19399 6010 19423 6012
rect 19479 6010 19503 6012
rect 19559 6010 19565 6012
rect 19319 5958 19321 6010
rect 19501 5958 19503 6010
rect 19257 5956 19263 5958
rect 19319 5956 19343 5958
rect 19399 5956 19423 5958
rect 19479 5956 19503 5958
rect 19559 5956 19565 5958
rect 19257 5947 19565 5956
rect 18340 5778 18460 5794
rect 18328 5772 18460 5778
rect 18380 5766 18460 5772
rect 18512 5772 18564 5778
rect 18328 5714 18380 5720
rect 18512 5714 18564 5720
rect 18340 4690 18368 5714
rect 18524 4826 18552 5714
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18340 4282 18368 4626
rect 18524 4282 18552 4762
rect 18800 4690 18828 4966
rect 19257 4924 19565 4933
rect 19257 4922 19263 4924
rect 19319 4922 19343 4924
rect 19399 4922 19423 4924
rect 19479 4922 19503 4924
rect 19559 4922 19565 4924
rect 19319 4870 19321 4922
rect 19501 4870 19503 4922
rect 19257 4868 19263 4870
rect 19319 4868 19343 4870
rect 19399 4868 19423 4870
rect 19479 4868 19503 4870
rect 19559 4868 19565 4870
rect 19257 4859 19565 4868
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18984 3602 19012 4694
rect 19257 3836 19565 3845
rect 19257 3834 19263 3836
rect 19319 3834 19343 3836
rect 19399 3834 19423 3836
rect 19479 3834 19503 3836
rect 19559 3834 19565 3836
rect 19319 3782 19321 3834
rect 19501 3782 19503 3834
rect 19257 3780 19263 3782
rect 19319 3780 19343 3782
rect 19399 3780 19423 3782
rect 19479 3780 19503 3782
rect 19559 3780 19565 3782
rect 19257 3771 19565 3780
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 18984 3058 19012 3538
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18524 1970 18552 2994
rect 19257 2748 19565 2757
rect 19257 2746 19263 2748
rect 19319 2746 19343 2748
rect 19399 2746 19423 2748
rect 19479 2746 19503 2748
rect 19559 2746 19565 2748
rect 19319 2694 19321 2746
rect 19501 2694 19503 2746
rect 19257 2692 19263 2694
rect 19319 2692 19343 2694
rect 19399 2692 19423 2694
rect 19479 2692 19503 2694
rect 19559 2692 19565 2694
rect 19257 2683 19565 2692
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 19076 2145 19104 2246
rect 19062 2136 19118 2145
rect 19062 2071 19118 2080
rect 18512 1964 18564 1970
rect 18512 1906 18564 1912
rect 19064 1896 19116 1902
rect 19064 1838 19116 1844
rect 18236 1556 18288 1562
rect 18236 1498 18288 1504
rect 19076 1465 19104 1838
rect 19257 1660 19565 1669
rect 19257 1658 19263 1660
rect 19319 1658 19343 1660
rect 19399 1658 19423 1660
rect 19479 1658 19503 1660
rect 19559 1658 19565 1660
rect 19319 1606 19321 1658
rect 19501 1606 19503 1658
rect 19257 1604 19263 1606
rect 19319 1604 19343 1606
rect 19399 1604 19423 1606
rect 19479 1604 19503 1606
rect 19559 1604 19565 1606
rect 19257 1595 19565 1604
rect 19062 1456 19118 1465
rect 16396 1420 16448 1426
rect 16396 1362 16448 1368
rect 16488 1420 16540 1426
rect 16488 1362 16540 1368
rect 16580 1420 16632 1426
rect 19062 1391 19118 1400
rect 16580 1362 16632 1368
rect 16304 1012 16356 1018
rect 16304 954 16356 960
rect 16316 814 16344 954
rect 16592 814 16620 1362
rect 16900 1116 17208 1125
rect 16900 1114 16906 1116
rect 16962 1114 16986 1116
rect 17042 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17208 1116
rect 16962 1062 16964 1114
rect 17144 1062 17146 1114
rect 16900 1060 16906 1062
rect 16962 1060 16986 1062
rect 17042 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17208 1062
rect 16900 1051 17208 1060
rect 3608 808 3660 814
rect 3608 750 3660 756
rect 6920 808 6972 814
rect 6920 750 6972 756
rect 10416 808 10468 814
rect 10416 750 10468 756
rect 13176 808 13228 814
rect 13176 750 13228 756
rect 16120 808 16172 814
rect 16120 750 16172 756
rect 16304 808 16356 814
rect 16304 750 16356 756
rect 16580 808 16632 814
rect 16580 750 16632 756
rect 18512 808 18564 814
rect 19064 808 19116 814
rect 18512 750 18564 756
rect 19062 776 19064 785
rect 19116 776 19118 785
rect 5112 572 5420 581
rect 5112 570 5118 572
rect 5174 570 5198 572
rect 5254 570 5278 572
rect 5334 570 5358 572
rect 5414 570 5420 572
rect 5174 518 5176 570
rect 5356 518 5358 570
rect 5112 516 5118 518
rect 5174 516 5198 518
rect 5254 516 5278 518
rect 5334 516 5358 518
rect 5414 516 5420 518
rect 5112 507 5420 516
rect 9827 572 10135 581
rect 9827 570 9833 572
rect 9889 570 9913 572
rect 9969 570 9993 572
rect 10049 570 10073 572
rect 10129 570 10135 572
rect 9889 518 9891 570
rect 10071 518 10073 570
rect 9827 516 9833 518
rect 9889 516 9913 518
rect 9969 516 9993 518
rect 10049 516 10073 518
rect 10129 516 10135 518
rect 9827 507 10135 516
rect 10428 490 10456 750
rect 11796 740 11848 746
rect 11796 682 11848 688
rect 12256 740 12308 746
rect 13084 740 13136 746
rect 12256 682 12308 688
rect 12912 700 13084 728
rect 11808 490 11836 682
rect 10336 462 10456 490
rect 11624 462 11836 490
rect 10336 400 10364 462
rect 11624 400 11652 462
rect 12268 400 12296 682
rect 12912 400 12940 700
rect 13084 682 13136 688
rect 14542 572 14850 581
rect 14542 570 14548 572
rect 14604 570 14628 572
rect 14684 570 14708 572
rect 14764 570 14788 572
rect 14844 570 14850 572
rect 14604 518 14606 570
rect 14786 518 14788 570
rect 14542 516 14548 518
rect 14604 516 14628 518
rect 14684 516 14708 518
rect 14764 516 14788 518
rect 14844 516 14850 518
rect 14542 507 14850 516
rect 18 0 74 400
rect 662 0 718 400
rect 1306 0 1362 400
rect 1950 0 2006 400
rect 2594 0 2650 400
rect 3238 0 3294 400
rect 3882 0 3938 400
rect 4526 0 4582 400
rect 5170 0 5226 400
rect 5814 0 5870 400
rect 6458 0 6514 400
rect 7102 0 7158 400
rect 7746 0 7802 400
rect 8390 0 8446 400
rect 9034 0 9090 400
rect 9678 0 9734 400
rect 10322 0 10378 400
rect 11610 0 11666 400
rect 12254 0 12310 400
rect 12898 0 12954 400
rect 18524 105 18552 750
rect 19062 711 19118 720
rect 19257 572 19565 581
rect 19257 570 19263 572
rect 19319 570 19343 572
rect 19399 570 19423 572
rect 19479 570 19503 572
rect 19559 570 19565 572
rect 19319 518 19321 570
rect 19501 518 19503 570
rect 19257 516 19263 518
rect 19319 516 19343 518
rect 19399 516 19423 518
rect 19479 516 19503 518
rect 19559 516 19565 518
rect 19257 507 19565 516
rect 18510 96 18566 105
rect 18510 31 18566 40
<< via2 >>
rect 1122 19760 1178 19816
rect 754 19080 810 19136
rect 5118 19066 5174 19068
rect 5198 19066 5254 19068
rect 5278 19066 5334 19068
rect 5358 19066 5414 19068
rect 5118 19014 5164 19066
rect 5164 19014 5174 19066
rect 5198 19014 5228 19066
rect 5228 19014 5240 19066
rect 5240 19014 5254 19066
rect 5278 19014 5292 19066
rect 5292 19014 5304 19066
rect 5304 19014 5334 19066
rect 5358 19014 5368 19066
rect 5368 19014 5414 19066
rect 5118 19012 5174 19014
rect 5198 19012 5254 19014
rect 5278 19012 5334 19014
rect 5358 19012 5414 19014
rect 9833 19066 9889 19068
rect 9913 19066 9969 19068
rect 9993 19066 10049 19068
rect 10073 19066 10129 19068
rect 9833 19014 9879 19066
rect 9879 19014 9889 19066
rect 9913 19014 9943 19066
rect 9943 19014 9955 19066
rect 9955 19014 9969 19066
rect 9993 19014 10007 19066
rect 10007 19014 10019 19066
rect 10019 19014 10049 19066
rect 10073 19014 10083 19066
rect 10083 19014 10129 19066
rect 9833 19012 9889 19014
rect 9913 19012 9969 19014
rect 9993 19012 10049 19014
rect 10073 19012 10129 19014
rect 2761 18522 2817 18524
rect 2841 18522 2897 18524
rect 2921 18522 2977 18524
rect 3001 18522 3057 18524
rect 2761 18470 2807 18522
rect 2807 18470 2817 18522
rect 2841 18470 2871 18522
rect 2871 18470 2883 18522
rect 2883 18470 2897 18522
rect 2921 18470 2935 18522
rect 2935 18470 2947 18522
rect 2947 18470 2977 18522
rect 3001 18470 3011 18522
rect 3011 18470 3057 18522
rect 2761 18468 2817 18470
rect 2841 18468 2897 18470
rect 2921 18468 2977 18470
rect 3001 18468 3057 18470
rect 7476 18522 7532 18524
rect 7556 18522 7612 18524
rect 7636 18522 7692 18524
rect 7716 18522 7772 18524
rect 7476 18470 7522 18522
rect 7522 18470 7532 18522
rect 7556 18470 7586 18522
rect 7586 18470 7598 18522
rect 7598 18470 7612 18522
rect 7636 18470 7650 18522
rect 7650 18470 7662 18522
rect 7662 18470 7692 18522
rect 7716 18470 7726 18522
rect 7726 18470 7772 18522
rect 7476 18468 7532 18470
rect 7556 18468 7612 18470
rect 7636 18468 7692 18470
rect 7716 18468 7772 18470
rect 846 18400 902 18456
rect 846 17720 902 17776
rect 846 17076 848 17096
rect 848 17076 900 17096
rect 900 17076 902 17096
rect 846 17040 902 17076
rect 2761 17434 2817 17436
rect 2841 17434 2897 17436
rect 2921 17434 2977 17436
rect 3001 17434 3057 17436
rect 2761 17382 2807 17434
rect 2807 17382 2817 17434
rect 2841 17382 2871 17434
rect 2871 17382 2883 17434
rect 2883 17382 2897 17434
rect 2921 17382 2935 17434
rect 2935 17382 2947 17434
rect 2947 17382 2977 17434
rect 3001 17382 3011 17434
rect 3011 17382 3057 17434
rect 2761 17380 2817 17382
rect 2841 17380 2897 17382
rect 2921 17380 2977 17382
rect 3001 17380 3057 17382
rect 5118 17978 5174 17980
rect 5198 17978 5254 17980
rect 5278 17978 5334 17980
rect 5358 17978 5414 17980
rect 5118 17926 5164 17978
rect 5164 17926 5174 17978
rect 5198 17926 5228 17978
rect 5228 17926 5240 17978
rect 5240 17926 5254 17978
rect 5278 17926 5292 17978
rect 5292 17926 5304 17978
rect 5304 17926 5334 17978
rect 5358 17926 5368 17978
rect 5368 17926 5414 17978
rect 5118 17924 5174 17926
rect 5198 17924 5254 17926
rect 5278 17924 5334 17926
rect 5358 17924 5414 17926
rect 2761 16346 2817 16348
rect 2841 16346 2897 16348
rect 2921 16346 2977 16348
rect 3001 16346 3057 16348
rect 2761 16294 2807 16346
rect 2807 16294 2817 16346
rect 2841 16294 2871 16346
rect 2871 16294 2883 16346
rect 2883 16294 2897 16346
rect 2921 16294 2935 16346
rect 2935 16294 2947 16346
rect 2947 16294 2977 16346
rect 3001 16294 3011 16346
rect 3011 16294 3057 16346
rect 2761 16292 2817 16294
rect 2841 16292 2897 16294
rect 2921 16292 2977 16294
rect 3001 16292 3057 16294
rect 3422 16088 3478 16144
rect 2761 15258 2817 15260
rect 2841 15258 2897 15260
rect 2921 15258 2977 15260
rect 3001 15258 3057 15260
rect 2761 15206 2807 15258
rect 2807 15206 2817 15258
rect 2841 15206 2871 15258
rect 2871 15206 2883 15258
rect 2883 15206 2897 15258
rect 2921 15206 2935 15258
rect 2935 15206 2947 15258
rect 2947 15206 2977 15258
rect 3001 15206 3011 15258
rect 3011 15206 3057 15258
rect 2761 15204 2817 15206
rect 2841 15204 2897 15206
rect 2921 15204 2977 15206
rect 3001 15204 3057 15206
rect 2761 14170 2817 14172
rect 2841 14170 2897 14172
rect 2921 14170 2977 14172
rect 3001 14170 3057 14172
rect 2761 14118 2807 14170
rect 2807 14118 2817 14170
rect 2841 14118 2871 14170
rect 2871 14118 2883 14170
rect 2883 14118 2897 14170
rect 2921 14118 2935 14170
rect 2935 14118 2947 14170
rect 2947 14118 2977 14170
rect 3001 14118 3011 14170
rect 3011 14118 3057 14170
rect 2761 14116 2817 14118
rect 2841 14116 2897 14118
rect 2921 14116 2977 14118
rect 3001 14116 3057 14118
rect 2761 13082 2817 13084
rect 2841 13082 2897 13084
rect 2921 13082 2977 13084
rect 3001 13082 3057 13084
rect 2761 13030 2807 13082
rect 2807 13030 2817 13082
rect 2841 13030 2871 13082
rect 2871 13030 2883 13082
rect 2883 13030 2897 13082
rect 2921 13030 2935 13082
rect 2935 13030 2947 13082
rect 2947 13030 2977 13082
rect 3001 13030 3011 13082
rect 3011 13030 3057 13082
rect 2761 13028 2817 13030
rect 2841 13028 2897 13030
rect 2921 13028 2977 13030
rect 3001 13028 3057 13030
rect 2761 11994 2817 11996
rect 2841 11994 2897 11996
rect 2921 11994 2977 11996
rect 3001 11994 3057 11996
rect 2761 11942 2807 11994
rect 2807 11942 2817 11994
rect 2841 11942 2871 11994
rect 2871 11942 2883 11994
rect 2883 11942 2897 11994
rect 2921 11942 2935 11994
rect 2935 11942 2947 11994
rect 2947 11942 2977 11994
rect 3001 11942 3011 11994
rect 3011 11942 3057 11994
rect 2761 11940 2817 11942
rect 2841 11940 2897 11942
rect 2921 11940 2977 11942
rect 3001 11940 3057 11942
rect 2761 10906 2817 10908
rect 2841 10906 2897 10908
rect 2921 10906 2977 10908
rect 3001 10906 3057 10908
rect 2761 10854 2807 10906
rect 2807 10854 2817 10906
rect 2841 10854 2871 10906
rect 2871 10854 2883 10906
rect 2883 10854 2897 10906
rect 2921 10854 2935 10906
rect 2935 10854 2947 10906
rect 2947 10854 2977 10906
rect 3001 10854 3011 10906
rect 3011 10854 3057 10906
rect 2761 10852 2817 10854
rect 2841 10852 2897 10854
rect 2921 10852 2977 10854
rect 3001 10852 3057 10854
rect 2761 9818 2817 9820
rect 2841 9818 2897 9820
rect 2921 9818 2977 9820
rect 3001 9818 3057 9820
rect 2761 9766 2807 9818
rect 2807 9766 2817 9818
rect 2841 9766 2871 9818
rect 2871 9766 2883 9818
rect 2883 9766 2897 9818
rect 2921 9766 2935 9818
rect 2935 9766 2947 9818
rect 2947 9766 2977 9818
rect 3001 9766 3011 9818
rect 3011 9766 3057 9818
rect 2761 9764 2817 9766
rect 2841 9764 2897 9766
rect 2921 9764 2977 9766
rect 3001 9764 3057 9766
rect 5118 16890 5174 16892
rect 5198 16890 5254 16892
rect 5278 16890 5334 16892
rect 5358 16890 5414 16892
rect 5118 16838 5164 16890
rect 5164 16838 5174 16890
rect 5198 16838 5228 16890
rect 5228 16838 5240 16890
rect 5240 16838 5254 16890
rect 5278 16838 5292 16890
rect 5292 16838 5304 16890
rect 5304 16838 5334 16890
rect 5358 16838 5368 16890
rect 5368 16838 5414 16890
rect 5118 16836 5174 16838
rect 5198 16836 5254 16838
rect 5278 16836 5334 16838
rect 5358 16836 5414 16838
rect 5118 15802 5174 15804
rect 5198 15802 5254 15804
rect 5278 15802 5334 15804
rect 5358 15802 5414 15804
rect 5118 15750 5164 15802
rect 5164 15750 5174 15802
rect 5198 15750 5228 15802
rect 5228 15750 5240 15802
rect 5240 15750 5254 15802
rect 5278 15750 5292 15802
rect 5292 15750 5304 15802
rect 5304 15750 5334 15802
rect 5358 15750 5368 15802
rect 5368 15750 5414 15802
rect 5118 15748 5174 15750
rect 5198 15748 5254 15750
rect 5278 15748 5334 15750
rect 5358 15748 5414 15750
rect 3606 11736 3662 11792
rect 2962 8880 3018 8936
rect 2761 8730 2817 8732
rect 2841 8730 2897 8732
rect 2921 8730 2977 8732
rect 3001 8730 3057 8732
rect 2761 8678 2807 8730
rect 2807 8678 2817 8730
rect 2841 8678 2871 8730
rect 2871 8678 2883 8730
rect 2883 8678 2897 8730
rect 2921 8678 2935 8730
rect 2935 8678 2947 8730
rect 2947 8678 2977 8730
rect 3001 8678 3011 8730
rect 3011 8678 3057 8730
rect 2761 8676 2817 8678
rect 2841 8676 2897 8678
rect 2921 8676 2977 8678
rect 3001 8676 3057 8678
rect 2761 7642 2817 7644
rect 2841 7642 2897 7644
rect 2921 7642 2977 7644
rect 3001 7642 3057 7644
rect 2761 7590 2807 7642
rect 2807 7590 2817 7642
rect 2841 7590 2871 7642
rect 2871 7590 2883 7642
rect 2883 7590 2897 7642
rect 2921 7590 2935 7642
rect 2935 7590 2947 7642
rect 2947 7590 2977 7642
rect 3001 7590 3011 7642
rect 3011 7590 3057 7642
rect 2761 7588 2817 7590
rect 2841 7588 2897 7590
rect 2921 7588 2977 7590
rect 3001 7588 3057 7590
rect 2761 6554 2817 6556
rect 2841 6554 2897 6556
rect 2921 6554 2977 6556
rect 3001 6554 3057 6556
rect 2761 6502 2807 6554
rect 2807 6502 2817 6554
rect 2841 6502 2871 6554
rect 2871 6502 2883 6554
rect 2883 6502 2897 6554
rect 2921 6502 2935 6554
rect 2935 6502 2947 6554
rect 2947 6502 2977 6554
rect 3001 6502 3011 6554
rect 3011 6502 3057 6554
rect 2761 6500 2817 6502
rect 2841 6500 2897 6502
rect 2921 6500 2977 6502
rect 3001 6500 3057 6502
rect 5118 14714 5174 14716
rect 5198 14714 5254 14716
rect 5278 14714 5334 14716
rect 5358 14714 5414 14716
rect 5118 14662 5164 14714
rect 5164 14662 5174 14714
rect 5198 14662 5228 14714
rect 5228 14662 5240 14714
rect 5240 14662 5254 14714
rect 5278 14662 5292 14714
rect 5292 14662 5304 14714
rect 5304 14662 5334 14714
rect 5358 14662 5368 14714
rect 5368 14662 5414 14714
rect 5118 14660 5174 14662
rect 5198 14660 5254 14662
rect 5278 14660 5334 14662
rect 5358 14660 5414 14662
rect 5118 13626 5174 13628
rect 5198 13626 5254 13628
rect 5278 13626 5334 13628
rect 5358 13626 5414 13628
rect 5118 13574 5164 13626
rect 5164 13574 5174 13626
rect 5198 13574 5228 13626
rect 5228 13574 5240 13626
rect 5240 13574 5254 13626
rect 5278 13574 5292 13626
rect 5292 13574 5304 13626
rect 5304 13574 5334 13626
rect 5358 13574 5368 13626
rect 5368 13574 5414 13626
rect 5118 13572 5174 13574
rect 5198 13572 5254 13574
rect 5278 13572 5334 13574
rect 5358 13572 5414 13574
rect 7476 17434 7532 17436
rect 7556 17434 7612 17436
rect 7636 17434 7692 17436
rect 7716 17434 7772 17436
rect 7476 17382 7522 17434
rect 7522 17382 7532 17434
rect 7556 17382 7586 17434
rect 7586 17382 7598 17434
rect 7598 17382 7612 17434
rect 7636 17382 7650 17434
rect 7650 17382 7662 17434
rect 7662 17382 7692 17434
rect 7716 17382 7726 17434
rect 7726 17382 7772 17434
rect 7476 17380 7532 17382
rect 7556 17380 7612 17382
rect 7636 17380 7692 17382
rect 7716 17380 7772 17382
rect 7476 16346 7532 16348
rect 7556 16346 7612 16348
rect 7636 16346 7692 16348
rect 7716 16346 7772 16348
rect 7476 16294 7522 16346
rect 7522 16294 7532 16346
rect 7556 16294 7586 16346
rect 7586 16294 7598 16346
rect 7598 16294 7612 16346
rect 7636 16294 7650 16346
rect 7650 16294 7662 16346
rect 7662 16294 7692 16346
rect 7716 16294 7726 16346
rect 7726 16294 7772 16346
rect 7476 16292 7532 16294
rect 7556 16292 7612 16294
rect 7636 16292 7692 16294
rect 7716 16292 7772 16294
rect 5118 12538 5174 12540
rect 5198 12538 5254 12540
rect 5278 12538 5334 12540
rect 5358 12538 5414 12540
rect 5118 12486 5164 12538
rect 5164 12486 5174 12538
rect 5198 12486 5228 12538
rect 5228 12486 5240 12538
rect 5240 12486 5254 12538
rect 5278 12486 5292 12538
rect 5292 12486 5304 12538
rect 5304 12486 5334 12538
rect 5358 12486 5368 12538
rect 5368 12486 5414 12538
rect 5118 12484 5174 12486
rect 5198 12484 5254 12486
rect 5278 12484 5334 12486
rect 5358 12484 5414 12486
rect 5118 11450 5174 11452
rect 5198 11450 5254 11452
rect 5278 11450 5334 11452
rect 5358 11450 5414 11452
rect 5118 11398 5164 11450
rect 5164 11398 5174 11450
rect 5198 11398 5228 11450
rect 5228 11398 5240 11450
rect 5240 11398 5254 11450
rect 5278 11398 5292 11450
rect 5292 11398 5304 11450
rect 5304 11398 5334 11450
rect 5358 11398 5368 11450
rect 5368 11398 5414 11450
rect 5118 11396 5174 11398
rect 5198 11396 5254 11398
rect 5278 11396 5334 11398
rect 5358 11396 5414 11398
rect 5118 10362 5174 10364
rect 5198 10362 5254 10364
rect 5278 10362 5334 10364
rect 5358 10362 5414 10364
rect 5118 10310 5164 10362
rect 5164 10310 5174 10362
rect 5198 10310 5228 10362
rect 5228 10310 5240 10362
rect 5240 10310 5254 10362
rect 5278 10310 5292 10362
rect 5292 10310 5304 10362
rect 5304 10310 5334 10362
rect 5358 10310 5368 10362
rect 5368 10310 5414 10362
rect 5118 10308 5174 10310
rect 5198 10308 5254 10310
rect 5278 10308 5334 10310
rect 5358 10308 5414 10310
rect 5262 9444 5318 9480
rect 5262 9424 5264 9444
rect 5264 9424 5316 9444
rect 5316 9424 5318 9444
rect 5118 9274 5174 9276
rect 5198 9274 5254 9276
rect 5278 9274 5334 9276
rect 5358 9274 5414 9276
rect 5118 9222 5164 9274
rect 5164 9222 5174 9274
rect 5198 9222 5228 9274
rect 5228 9222 5240 9274
rect 5240 9222 5254 9274
rect 5278 9222 5292 9274
rect 5292 9222 5304 9274
rect 5304 9222 5334 9274
rect 5358 9222 5368 9274
rect 5368 9222 5414 9274
rect 5118 9220 5174 9222
rect 5198 9220 5254 9222
rect 5278 9220 5334 9222
rect 5358 9220 5414 9222
rect 5354 9036 5410 9072
rect 5354 9016 5356 9036
rect 5356 9016 5408 9036
rect 5408 9016 5410 9036
rect 5722 9968 5778 10024
rect 2761 5466 2817 5468
rect 2841 5466 2897 5468
rect 2921 5466 2977 5468
rect 3001 5466 3057 5468
rect 2761 5414 2807 5466
rect 2807 5414 2817 5466
rect 2841 5414 2871 5466
rect 2871 5414 2883 5466
rect 2883 5414 2897 5466
rect 2921 5414 2935 5466
rect 2935 5414 2947 5466
rect 2947 5414 2977 5466
rect 3001 5414 3011 5466
rect 3011 5414 3057 5466
rect 2761 5412 2817 5414
rect 2841 5412 2897 5414
rect 2921 5412 2977 5414
rect 3001 5412 3057 5414
rect 3054 5072 3110 5128
rect 2761 4378 2817 4380
rect 2841 4378 2897 4380
rect 2921 4378 2977 4380
rect 3001 4378 3057 4380
rect 2761 4326 2807 4378
rect 2807 4326 2817 4378
rect 2841 4326 2871 4378
rect 2871 4326 2883 4378
rect 2883 4326 2897 4378
rect 2921 4326 2935 4378
rect 2935 4326 2947 4378
rect 2947 4326 2977 4378
rect 3001 4326 3011 4378
rect 3011 4326 3057 4378
rect 2761 4324 2817 4326
rect 2841 4324 2897 4326
rect 2921 4324 2977 4326
rect 3001 4324 3057 4326
rect 2761 3290 2817 3292
rect 2841 3290 2897 3292
rect 2921 3290 2977 3292
rect 3001 3290 3057 3292
rect 2761 3238 2807 3290
rect 2807 3238 2817 3290
rect 2841 3238 2871 3290
rect 2871 3238 2883 3290
rect 2883 3238 2897 3290
rect 2921 3238 2935 3290
rect 2935 3238 2947 3290
rect 2947 3238 2977 3290
rect 3001 3238 3011 3290
rect 3011 3238 3057 3290
rect 2761 3236 2817 3238
rect 2841 3236 2897 3238
rect 2921 3236 2977 3238
rect 3001 3236 3057 3238
rect 5118 8186 5174 8188
rect 5198 8186 5254 8188
rect 5278 8186 5334 8188
rect 5358 8186 5414 8188
rect 5118 8134 5164 8186
rect 5164 8134 5174 8186
rect 5198 8134 5228 8186
rect 5228 8134 5240 8186
rect 5240 8134 5254 8186
rect 5278 8134 5292 8186
rect 5292 8134 5304 8186
rect 5304 8134 5334 8186
rect 5358 8134 5368 8186
rect 5368 8134 5414 8186
rect 5118 8132 5174 8134
rect 5198 8132 5254 8134
rect 5278 8132 5334 8134
rect 5358 8132 5414 8134
rect 5118 7098 5174 7100
rect 5198 7098 5254 7100
rect 5278 7098 5334 7100
rect 5358 7098 5414 7100
rect 5118 7046 5164 7098
rect 5164 7046 5174 7098
rect 5198 7046 5228 7098
rect 5228 7046 5240 7098
rect 5240 7046 5254 7098
rect 5278 7046 5292 7098
rect 5292 7046 5304 7098
rect 5304 7046 5334 7098
rect 5358 7046 5368 7098
rect 5368 7046 5414 7098
rect 5118 7044 5174 7046
rect 5198 7044 5254 7046
rect 5278 7044 5334 7046
rect 5358 7044 5414 7046
rect 6274 9036 6330 9072
rect 6274 9016 6276 9036
rect 6276 9016 6328 9036
rect 6328 9016 6330 9036
rect 5118 6010 5174 6012
rect 5198 6010 5254 6012
rect 5278 6010 5334 6012
rect 5358 6010 5414 6012
rect 5118 5958 5164 6010
rect 5164 5958 5174 6010
rect 5198 5958 5228 6010
rect 5228 5958 5240 6010
rect 5240 5958 5254 6010
rect 5278 5958 5292 6010
rect 5292 5958 5304 6010
rect 5304 5958 5334 6010
rect 5358 5958 5368 6010
rect 5368 5958 5414 6010
rect 5118 5956 5174 5958
rect 5198 5956 5254 5958
rect 5278 5956 5334 5958
rect 5358 5956 5414 5958
rect 5118 4922 5174 4924
rect 5198 4922 5254 4924
rect 5278 4922 5334 4924
rect 5358 4922 5414 4924
rect 5118 4870 5164 4922
rect 5164 4870 5174 4922
rect 5198 4870 5228 4922
rect 5228 4870 5240 4922
rect 5240 4870 5254 4922
rect 5278 4870 5292 4922
rect 5292 4870 5304 4922
rect 5304 4870 5334 4922
rect 5358 4870 5368 4922
rect 5368 4870 5414 4922
rect 5118 4868 5174 4870
rect 5198 4868 5254 4870
rect 5278 4868 5334 4870
rect 5358 4868 5414 4870
rect 5118 3834 5174 3836
rect 5198 3834 5254 3836
rect 5278 3834 5334 3836
rect 5358 3834 5414 3836
rect 5118 3782 5164 3834
rect 5164 3782 5174 3834
rect 5198 3782 5228 3834
rect 5228 3782 5240 3834
rect 5240 3782 5254 3834
rect 5278 3782 5292 3834
rect 5292 3782 5304 3834
rect 5304 3782 5334 3834
rect 5358 3782 5368 3834
rect 5368 3782 5414 3834
rect 5118 3780 5174 3782
rect 5198 3780 5254 3782
rect 5278 3780 5334 3782
rect 5358 3780 5414 3782
rect 5118 2746 5174 2748
rect 5198 2746 5254 2748
rect 5278 2746 5334 2748
rect 5358 2746 5414 2748
rect 5118 2694 5164 2746
rect 5164 2694 5174 2746
rect 5198 2694 5228 2746
rect 5228 2694 5240 2746
rect 5240 2694 5254 2746
rect 5278 2694 5292 2746
rect 5292 2694 5304 2746
rect 5304 2694 5334 2746
rect 5358 2694 5368 2746
rect 5368 2694 5414 2746
rect 5118 2692 5174 2694
rect 5198 2692 5254 2694
rect 5278 2692 5334 2694
rect 5358 2692 5414 2694
rect 2761 2202 2817 2204
rect 2841 2202 2897 2204
rect 2921 2202 2977 2204
rect 3001 2202 3057 2204
rect 2761 2150 2807 2202
rect 2807 2150 2817 2202
rect 2841 2150 2871 2202
rect 2871 2150 2883 2202
rect 2883 2150 2897 2202
rect 2921 2150 2935 2202
rect 2935 2150 2947 2202
rect 2947 2150 2977 2202
rect 3001 2150 3011 2202
rect 3011 2150 3057 2202
rect 2761 2148 2817 2150
rect 2841 2148 2897 2150
rect 2921 2148 2977 2150
rect 3001 2148 3057 2150
rect 4802 1808 4858 1864
rect 2761 1114 2817 1116
rect 2841 1114 2897 1116
rect 2921 1114 2977 1116
rect 3001 1114 3057 1116
rect 2761 1062 2807 1114
rect 2807 1062 2817 1114
rect 2841 1062 2871 1114
rect 2871 1062 2883 1114
rect 2883 1062 2897 1114
rect 2921 1062 2935 1114
rect 2935 1062 2947 1114
rect 2947 1062 2977 1114
rect 3001 1062 3011 1114
rect 3011 1062 3057 1114
rect 2761 1060 2817 1062
rect 2841 1060 2897 1062
rect 2921 1060 2977 1062
rect 3001 1060 3057 1062
rect 5118 1658 5174 1660
rect 5198 1658 5254 1660
rect 5278 1658 5334 1660
rect 5358 1658 5414 1660
rect 5118 1606 5164 1658
rect 5164 1606 5174 1658
rect 5198 1606 5228 1658
rect 5228 1606 5240 1658
rect 5240 1606 5254 1658
rect 5278 1606 5292 1658
rect 5292 1606 5304 1658
rect 5304 1606 5334 1658
rect 5358 1606 5368 1658
rect 5368 1606 5414 1658
rect 5118 1604 5174 1606
rect 5198 1604 5254 1606
rect 5278 1604 5334 1606
rect 5358 1604 5414 1606
rect 7476 15258 7532 15260
rect 7556 15258 7612 15260
rect 7636 15258 7692 15260
rect 7716 15258 7772 15260
rect 7476 15206 7522 15258
rect 7522 15206 7532 15258
rect 7556 15206 7586 15258
rect 7586 15206 7598 15258
rect 7598 15206 7612 15258
rect 7636 15206 7650 15258
rect 7650 15206 7662 15258
rect 7662 15206 7692 15258
rect 7716 15206 7726 15258
rect 7726 15206 7772 15258
rect 7476 15204 7532 15206
rect 7556 15204 7612 15206
rect 7636 15204 7692 15206
rect 7716 15204 7772 15206
rect 7476 14170 7532 14172
rect 7556 14170 7612 14172
rect 7636 14170 7692 14172
rect 7716 14170 7772 14172
rect 7476 14118 7522 14170
rect 7522 14118 7532 14170
rect 7556 14118 7586 14170
rect 7586 14118 7598 14170
rect 7598 14118 7612 14170
rect 7636 14118 7650 14170
rect 7650 14118 7662 14170
rect 7662 14118 7692 14170
rect 7716 14118 7726 14170
rect 7726 14118 7772 14170
rect 7476 14116 7532 14118
rect 7556 14116 7612 14118
rect 7636 14116 7692 14118
rect 7716 14116 7772 14118
rect 7476 13082 7532 13084
rect 7556 13082 7612 13084
rect 7636 13082 7692 13084
rect 7716 13082 7772 13084
rect 7476 13030 7522 13082
rect 7522 13030 7532 13082
rect 7556 13030 7586 13082
rect 7586 13030 7598 13082
rect 7598 13030 7612 13082
rect 7636 13030 7650 13082
rect 7650 13030 7662 13082
rect 7662 13030 7692 13082
rect 7716 13030 7726 13082
rect 7726 13030 7772 13082
rect 7476 13028 7532 13030
rect 7556 13028 7612 13030
rect 7636 13028 7692 13030
rect 7716 13028 7772 13030
rect 7476 11994 7532 11996
rect 7556 11994 7612 11996
rect 7636 11994 7692 11996
rect 7716 11994 7772 11996
rect 7476 11942 7522 11994
rect 7522 11942 7532 11994
rect 7556 11942 7586 11994
rect 7586 11942 7598 11994
rect 7598 11942 7612 11994
rect 7636 11942 7650 11994
rect 7650 11942 7662 11994
rect 7662 11942 7692 11994
rect 7716 11942 7726 11994
rect 7726 11942 7772 11994
rect 7476 11940 7532 11942
rect 7556 11940 7612 11942
rect 7636 11940 7692 11942
rect 7716 11940 7772 11942
rect 7476 10906 7532 10908
rect 7556 10906 7612 10908
rect 7636 10906 7692 10908
rect 7716 10906 7772 10908
rect 7476 10854 7522 10906
rect 7522 10854 7532 10906
rect 7556 10854 7586 10906
rect 7586 10854 7598 10906
rect 7598 10854 7612 10906
rect 7636 10854 7650 10906
rect 7650 10854 7662 10906
rect 7662 10854 7692 10906
rect 7716 10854 7726 10906
rect 7726 10854 7772 10906
rect 7476 10852 7532 10854
rect 7556 10852 7612 10854
rect 7636 10852 7692 10854
rect 7716 10852 7772 10854
rect 7562 9968 7618 10024
rect 7476 9818 7532 9820
rect 7556 9818 7612 9820
rect 7636 9818 7692 9820
rect 7716 9818 7772 9820
rect 7476 9766 7522 9818
rect 7522 9766 7532 9818
rect 7556 9766 7586 9818
rect 7586 9766 7598 9818
rect 7598 9766 7612 9818
rect 7636 9766 7650 9818
rect 7650 9766 7662 9818
rect 7662 9766 7692 9818
rect 7716 9766 7726 9818
rect 7726 9766 7772 9818
rect 7476 9764 7532 9766
rect 7556 9764 7612 9766
rect 7636 9764 7692 9766
rect 7716 9764 7772 9766
rect 7838 9424 7894 9480
rect 7476 8730 7532 8732
rect 7556 8730 7612 8732
rect 7636 8730 7692 8732
rect 7716 8730 7772 8732
rect 7476 8678 7522 8730
rect 7522 8678 7532 8730
rect 7556 8678 7586 8730
rect 7586 8678 7598 8730
rect 7598 8678 7612 8730
rect 7636 8678 7650 8730
rect 7650 8678 7662 8730
rect 7662 8678 7692 8730
rect 7716 8678 7726 8730
rect 7726 8678 7772 8730
rect 7476 8676 7532 8678
rect 7556 8676 7612 8678
rect 7636 8676 7692 8678
rect 7716 8676 7772 8678
rect 9833 17978 9889 17980
rect 9913 17978 9969 17980
rect 9993 17978 10049 17980
rect 10073 17978 10129 17980
rect 9833 17926 9879 17978
rect 9879 17926 9889 17978
rect 9913 17926 9943 17978
rect 9943 17926 9955 17978
rect 9955 17926 9969 17978
rect 9993 17926 10007 17978
rect 10007 17926 10019 17978
rect 10019 17926 10049 17978
rect 10073 17926 10083 17978
rect 10083 17926 10129 17978
rect 9833 17924 9889 17926
rect 9913 17924 9969 17926
rect 9993 17924 10049 17926
rect 10073 17924 10129 17926
rect 7476 7642 7532 7644
rect 7556 7642 7612 7644
rect 7636 7642 7692 7644
rect 7716 7642 7772 7644
rect 7476 7590 7522 7642
rect 7522 7590 7532 7642
rect 7556 7590 7586 7642
rect 7586 7590 7598 7642
rect 7598 7590 7612 7642
rect 7636 7590 7650 7642
rect 7650 7590 7662 7642
rect 7662 7590 7692 7642
rect 7716 7590 7726 7642
rect 7726 7590 7772 7642
rect 7476 7588 7532 7590
rect 7556 7588 7612 7590
rect 7636 7588 7692 7590
rect 7716 7588 7772 7590
rect 8666 12708 8722 12744
rect 8666 12688 8668 12708
rect 8668 12688 8720 12708
rect 8720 12688 8722 12708
rect 8666 12280 8722 12336
rect 7286 6296 7342 6352
rect 7476 6554 7532 6556
rect 7556 6554 7612 6556
rect 7636 6554 7692 6556
rect 7716 6554 7772 6556
rect 7476 6502 7522 6554
rect 7522 6502 7532 6554
rect 7556 6502 7586 6554
rect 7586 6502 7598 6554
rect 7598 6502 7612 6554
rect 7636 6502 7650 6554
rect 7650 6502 7662 6554
rect 7662 6502 7692 6554
rect 7716 6502 7726 6554
rect 7726 6502 7772 6554
rect 7476 6500 7532 6502
rect 7556 6500 7612 6502
rect 7636 6500 7692 6502
rect 7716 6500 7772 6502
rect 7476 5466 7532 5468
rect 7556 5466 7612 5468
rect 7636 5466 7692 5468
rect 7716 5466 7772 5468
rect 7476 5414 7522 5466
rect 7522 5414 7532 5466
rect 7556 5414 7586 5466
rect 7586 5414 7598 5466
rect 7598 5414 7612 5466
rect 7636 5414 7650 5466
rect 7650 5414 7662 5466
rect 7662 5414 7692 5466
rect 7716 5414 7726 5466
rect 7726 5414 7772 5466
rect 7476 5412 7532 5414
rect 7556 5412 7612 5414
rect 7636 5412 7692 5414
rect 7716 5412 7772 5414
rect 7476 4378 7532 4380
rect 7556 4378 7612 4380
rect 7636 4378 7692 4380
rect 7716 4378 7772 4380
rect 7476 4326 7522 4378
rect 7522 4326 7532 4378
rect 7556 4326 7586 4378
rect 7586 4326 7598 4378
rect 7598 4326 7612 4378
rect 7636 4326 7650 4378
rect 7650 4326 7662 4378
rect 7662 4326 7692 4378
rect 7716 4326 7726 4378
rect 7726 4326 7772 4378
rect 7476 4324 7532 4326
rect 7556 4324 7612 4326
rect 7636 4324 7692 4326
rect 7716 4324 7772 4326
rect 7476 3290 7532 3292
rect 7556 3290 7612 3292
rect 7636 3290 7692 3292
rect 7716 3290 7772 3292
rect 7476 3238 7522 3290
rect 7522 3238 7532 3290
rect 7556 3238 7586 3290
rect 7586 3238 7598 3290
rect 7598 3238 7612 3290
rect 7636 3238 7650 3290
rect 7650 3238 7662 3290
rect 7662 3238 7692 3290
rect 7716 3238 7726 3290
rect 7726 3238 7772 3290
rect 7476 3236 7532 3238
rect 7556 3236 7612 3238
rect 7636 3236 7692 3238
rect 7716 3236 7772 3238
rect 7476 2202 7532 2204
rect 7556 2202 7612 2204
rect 7636 2202 7692 2204
rect 7716 2202 7772 2204
rect 7476 2150 7522 2202
rect 7522 2150 7532 2202
rect 7556 2150 7586 2202
rect 7586 2150 7598 2202
rect 7598 2150 7612 2202
rect 7636 2150 7650 2202
rect 7650 2150 7662 2202
rect 7662 2150 7692 2202
rect 7716 2150 7726 2202
rect 7726 2150 7772 2202
rect 7476 2148 7532 2150
rect 7556 2148 7612 2150
rect 7636 2148 7692 2150
rect 7716 2148 7772 2150
rect 9833 16890 9889 16892
rect 9913 16890 9969 16892
rect 9993 16890 10049 16892
rect 10073 16890 10129 16892
rect 9833 16838 9879 16890
rect 9879 16838 9889 16890
rect 9913 16838 9943 16890
rect 9943 16838 9955 16890
rect 9955 16838 9969 16890
rect 9993 16838 10007 16890
rect 10007 16838 10019 16890
rect 10019 16838 10049 16890
rect 10073 16838 10083 16890
rect 10083 16838 10129 16890
rect 9833 16836 9889 16838
rect 9913 16836 9969 16838
rect 9993 16836 10049 16838
rect 10073 16836 10129 16838
rect 9833 15802 9889 15804
rect 9913 15802 9969 15804
rect 9993 15802 10049 15804
rect 10073 15802 10129 15804
rect 9833 15750 9879 15802
rect 9879 15750 9889 15802
rect 9913 15750 9943 15802
rect 9943 15750 9955 15802
rect 9955 15750 9969 15802
rect 9993 15750 10007 15802
rect 10007 15750 10019 15802
rect 10019 15750 10049 15802
rect 10073 15750 10083 15802
rect 10083 15750 10129 15802
rect 9833 15748 9889 15750
rect 9913 15748 9969 15750
rect 9993 15748 10049 15750
rect 10073 15748 10129 15750
rect 9833 14714 9889 14716
rect 9913 14714 9969 14716
rect 9993 14714 10049 14716
rect 10073 14714 10129 14716
rect 9833 14662 9879 14714
rect 9879 14662 9889 14714
rect 9913 14662 9943 14714
rect 9943 14662 9955 14714
rect 9955 14662 9969 14714
rect 9993 14662 10007 14714
rect 10007 14662 10019 14714
rect 10019 14662 10049 14714
rect 10073 14662 10083 14714
rect 10083 14662 10129 14714
rect 9833 14660 9889 14662
rect 9913 14660 9969 14662
rect 9993 14660 10049 14662
rect 10073 14660 10129 14662
rect 9833 13626 9889 13628
rect 9913 13626 9969 13628
rect 9993 13626 10049 13628
rect 10073 13626 10129 13628
rect 9833 13574 9879 13626
rect 9879 13574 9889 13626
rect 9913 13574 9943 13626
rect 9943 13574 9955 13626
rect 9955 13574 9969 13626
rect 9993 13574 10007 13626
rect 10007 13574 10019 13626
rect 10019 13574 10049 13626
rect 10073 13574 10083 13626
rect 10083 13574 10129 13626
rect 9833 13572 9889 13574
rect 9913 13572 9969 13574
rect 9993 13572 10049 13574
rect 10073 13572 10129 13574
rect 10138 12860 10140 12880
rect 10140 12860 10192 12880
rect 10192 12860 10194 12880
rect 10138 12824 10194 12860
rect 9833 12538 9889 12540
rect 9913 12538 9969 12540
rect 9993 12538 10049 12540
rect 10073 12538 10129 12540
rect 9833 12486 9879 12538
rect 9879 12486 9889 12538
rect 9913 12486 9943 12538
rect 9943 12486 9955 12538
rect 9955 12486 9969 12538
rect 9993 12486 10007 12538
rect 10007 12486 10019 12538
rect 10019 12486 10049 12538
rect 10073 12486 10083 12538
rect 10083 12486 10129 12538
rect 9833 12484 9889 12486
rect 9913 12484 9969 12486
rect 9993 12484 10049 12486
rect 10073 12484 10129 12486
rect 14548 19066 14604 19068
rect 14628 19066 14684 19068
rect 14708 19066 14764 19068
rect 14788 19066 14844 19068
rect 14548 19014 14594 19066
rect 14594 19014 14604 19066
rect 14628 19014 14658 19066
rect 14658 19014 14670 19066
rect 14670 19014 14684 19066
rect 14708 19014 14722 19066
rect 14722 19014 14734 19066
rect 14734 19014 14764 19066
rect 14788 19014 14798 19066
rect 14798 19014 14844 19066
rect 14548 19012 14604 19014
rect 14628 19012 14684 19014
rect 14708 19012 14764 19014
rect 14788 19012 14844 19014
rect 19263 19066 19319 19068
rect 19343 19066 19399 19068
rect 19423 19066 19479 19068
rect 19503 19066 19559 19068
rect 19263 19014 19309 19066
rect 19309 19014 19319 19066
rect 19343 19014 19373 19066
rect 19373 19014 19385 19066
rect 19385 19014 19399 19066
rect 19423 19014 19437 19066
rect 19437 19014 19449 19066
rect 19449 19014 19479 19066
rect 19503 19014 19513 19066
rect 19513 19014 19559 19066
rect 19263 19012 19319 19014
rect 19343 19012 19399 19014
rect 19423 19012 19479 19014
rect 19503 19012 19559 19014
rect 11150 15988 11152 16008
rect 11152 15988 11204 16008
rect 11204 15988 11206 16008
rect 11150 15952 11206 15988
rect 9770 11600 9826 11656
rect 10322 11736 10378 11792
rect 9833 11450 9889 11452
rect 9913 11450 9969 11452
rect 9993 11450 10049 11452
rect 10073 11450 10129 11452
rect 9833 11398 9879 11450
rect 9879 11398 9889 11450
rect 9913 11398 9943 11450
rect 9943 11398 9955 11450
rect 9955 11398 9969 11450
rect 9993 11398 10007 11450
rect 10007 11398 10019 11450
rect 10019 11398 10049 11450
rect 10073 11398 10083 11450
rect 10083 11398 10129 11450
rect 9833 11396 9889 11398
rect 9913 11396 9969 11398
rect 9993 11396 10049 11398
rect 10073 11396 10129 11398
rect 9034 7268 9090 7304
rect 9034 7248 9036 7268
rect 9036 7248 9088 7268
rect 9088 7248 9090 7268
rect 9126 6976 9182 7032
rect 9586 9016 9642 9072
rect 9770 10532 9826 10568
rect 9770 10512 9772 10532
rect 9772 10512 9824 10532
rect 9824 10512 9826 10532
rect 9833 10362 9889 10364
rect 9913 10362 9969 10364
rect 9993 10362 10049 10364
rect 10073 10362 10129 10364
rect 9833 10310 9879 10362
rect 9879 10310 9889 10362
rect 9913 10310 9943 10362
rect 9943 10310 9955 10362
rect 9955 10310 9969 10362
rect 9993 10310 10007 10362
rect 10007 10310 10019 10362
rect 10019 10310 10049 10362
rect 10073 10310 10083 10362
rect 10083 10310 10129 10362
rect 9833 10308 9889 10310
rect 9913 10308 9969 10310
rect 9993 10308 10049 10310
rect 10073 10308 10129 10310
rect 10690 12552 10746 12608
rect 9833 9274 9889 9276
rect 9913 9274 9969 9276
rect 9993 9274 10049 9276
rect 10073 9274 10129 9276
rect 9833 9222 9879 9274
rect 9879 9222 9889 9274
rect 9913 9222 9943 9274
rect 9943 9222 9955 9274
rect 9955 9222 9969 9274
rect 9993 9222 10007 9274
rect 10007 9222 10019 9274
rect 10019 9222 10049 9274
rect 10073 9222 10083 9274
rect 10083 9222 10129 9274
rect 9833 9220 9889 9222
rect 9913 9220 9969 9222
rect 9993 9220 10049 9222
rect 10073 9220 10129 9222
rect 9770 8508 9772 8528
rect 9772 8508 9824 8528
rect 9824 8508 9826 8528
rect 9770 8472 9826 8508
rect 9833 8186 9889 8188
rect 9913 8186 9969 8188
rect 9993 8186 10049 8188
rect 10073 8186 10129 8188
rect 9833 8134 9879 8186
rect 9879 8134 9889 8186
rect 9913 8134 9943 8186
rect 9943 8134 9955 8186
rect 9955 8134 9969 8186
rect 9993 8134 10007 8186
rect 10007 8134 10019 8186
rect 10019 8134 10049 8186
rect 10073 8134 10083 8186
rect 10083 8134 10129 8186
rect 9833 8132 9889 8134
rect 9913 8132 9969 8134
rect 9993 8132 10049 8134
rect 10073 8132 10129 8134
rect 9586 7248 9642 7304
rect 9494 6976 9550 7032
rect 9833 7098 9889 7100
rect 9913 7098 9969 7100
rect 9993 7098 10049 7100
rect 10073 7098 10129 7100
rect 9833 7046 9879 7098
rect 9879 7046 9889 7098
rect 9913 7046 9943 7098
rect 9943 7046 9955 7098
rect 9955 7046 9969 7098
rect 9993 7046 10007 7098
rect 10007 7046 10019 7098
rect 10019 7046 10049 7098
rect 10073 7046 10083 7098
rect 10083 7046 10129 7098
rect 9833 7044 9889 7046
rect 9913 7044 9969 7046
rect 9993 7044 10049 7046
rect 10073 7044 10129 7046
rect 8850 5752 8906 5808
rect 9034 5616 9090 5672
rect 9402 5772 9458 5808
rect 9402 5752 9404 5772
rect 9404 5752 9456 5772
rect 9456 5752 9458 5772
rect 9310 5616 9366 5672
rect 9586 6840 9642 6896
rect 9833 6010 9889 6012
rect 9913 6010 9969 6012
rect 9993 6010 10049 6012
rect 10073 6010 10129 6012
rect 9833 5958 9879 6010
rect 9879 5958 9889 6010
rect 9913 5958 9943 6010
rect 9943 5958 9955 6010
rect 9955 5958 9969 6010
rect 9993 5958 10007 6010
rect 10007 5958 10019 6010
rect 10019 5958 10049 6010
rect 10073 5958 10083 6010
rect 10083 5958 10129 6010
rect 9833 5956 9889 5958
rect 9913 5956 9969 5958
rect 9993 5956 10049 5958
rect 10073 5956 10129 5958
rect 9678 5636 9734 5672
rect 9678 5616 9680 5636
rect 9680 5616 9732 5636
rect 9732 5616 9734 5636
rect 9833 4922 9889 4924
rect 9913 4922 9969 4924
rect 9993 4922 10049 4924
rect 10073 4922 10129 4924
rect 9833 4870 9879 4922
rect 9879 4870 9889 4922
rect 9913 4870 9943 4922
rect 9943 4870 9955 4922
rect 9955 4870 9969 4922
rect 9993 4870 10007 4922
rect 10007 4870 10019 4922
rect 10019 4870 10049 4922
rect 10073 4870 10083 4922
rect 10083 4870 10129 4922
rect 9833 4868 9889 4870
rect 9913 4868 9969 4870
rect 9993 4868 10049 4870
rect 10073 4868 10129 4870
rect 9833 3834 9889 3836
rect 9913 3834 9969 3836
rect 9993 3834 10049 3836
rect 10073 3834 10129 3836
rect 9833 3782 9879 3834
rect 9879 3782 9889 3834
rect 9913 3782 9943 3834
rect 9943 3782 9955 3834
rect 9955 3782 9969 3834
rect 9993 3782 10007 3834
rect 10007 3782 10019 3834
rect 10019 3782 10049 3834
rect 10073 3782 10083 3834
rect 10083 3782 10129 3834
rect 9833 3780 9889 3782
rect 9913 3780 9969 3782
rect 9993 3780 10049 3782
rect 10073 3780 10129 3782
rect 10690 9968 10746 10024
rect 10690 9460 10692 9480
rect 10692 9460 10744 9480
rect 10744 9460 10746 9480
rect 10690 9424 10746 9460
rect 10782 5752 10838 5808
rect 11242 9696 11298 9752
rect 12191 18522 12247 18524
rect 12271 18522 12327 18524
rect 12351 18522 12407 18524
rect 12431 18522 12487 18524
rect 12191 18470 12237 18522
rect 12237 18470 12247 18522
rect 12271 18470 12301 18522
rect 12301 18470 12313 18522
rect 12313 18470 12327 18522
rect 12351 18470 12365 18522
rect 12365 18470 12377 18522
rect 12377 18470 12407 18522
rect 12431 18470 12441 18522
rect 12441 18470 12487 18522
rect 12191 18468 12247 18470
rect 12271 18468 12327 18470
rect 12351 18468 12407 18470
rect 12431 18468 12487 18470
rect 12191 17434 12247 17436
rect 12271 17434 12327 17436
rect 12351 17434 12407 17436
rect 12431 17434 12487 17436
rect 12191 17382 12237 17434
rect 12237 17382 12247 17434
rect 12271 17382 12301 17434
rect 12301 17382 12313 17434
rect 12313 17382 12327 17434
rect 12351 17382 12365 17434
rect 12365 17382 12377 17434
rect 12377 17382 12407 17434
rect 12431 17382 12441 17434
rect 12441 17382 12487 17434
rect 12191 17380 12247 17382
rect 12271 17380 12327 17382
rect 12351 17380 12407 17382
rect 12431 17380 12487 17382
rect 12191 16346 12247 16348
rect 12271 16346 12327 16348
rect 12351 16346 12407 16348
rect 12431 16346 12487 16348
rect 12191 16294 12237 16346
rect 12237 16294 12247 16346
rect 12271 16294 12301 16346
rect 12301 16294 12313 16346
rect 12313 16294 12327 16346
rect 12351 16294 12365 16346
rect 12365 16294 12377 16346
rect 12377 16294 12407 16346
rect 12431 16294 12441 16346
rect 12441 16294 12487 16346
rect 12191 16292 12247 16294
rect 12271 16292 12327 16294
rect 12351 16292 12407 16294
rect 12431 16292 12487 16294
rect 11702 11736 11758 11792
rect 12070 15408 12126 15464
rect 12191 15258 12247 15260
rect 12271 15258 12327 15260
rect 12351 15258 12407 15260
rect 12431 15258 12487 15260
rect 12191 15206 12237 15258
rect 12237 15206 12247 15258
rect 12271 15206 12301 15258
rect 12301 15206 12313 15258
rect 12313 15206 12327 15258
rect 12351 15206 12365 15258
rect 12365 15206 12377 15258
rect 12377 15206 12407 15258
rect 12431 15206 12441 15258
rect 12441 15206 12487 15258
rect 12191 15204 12247 15206
rect 12271 15204 12327 15206
rect 12351 15204 12407 15206
rect 12431 15204 12487 15206
rect 12191 14170 12247 14172
rect 12271 14170 12327 14172
rect 12351 14170 12407 14172
rect 12431 14170 12487 14172
rect 12191 14118 12237 14170
rect 12237 14118 12247 14170
rect 12271 14118 12301 14170
rect 12301 14118 12313 14170
rect 12313 14118 12327 14170
rect 12351 14118 12365 14170
rect 12365 14118 12377 14170
rect 12377 14118 12407 14170
rect 12431 14118 12441 14170
rect 12441 14118 12487 14170
rect 12191 14116 12247 14118
rect 12271 14116 12327 14118
rect 12351 14116 12407 14118
rect 12431 14116 12487 14118
rect 12191 13082 12247 13084
rect 12271 13082 12327 13084
rect 12351 13082 12407 13084
rect 12431 13082 12487 13084
rect 12191 13030 12237 13082
rect 12237 13030 12247 13082
rect 12271 13030 12301 13082
rect 12301 13030 12313 13082
rect 12313 13030 12327 13082
rect 12351 13030 12365 13082
rect 12365 13030 12377 13082
rect 12377 13030 12407 13082
rect 12431 13030 12441 13082
rect 12441 13030 12487 13082
rect 12191 13028 12247 13030
rect 12271 13028 12327 13030
rect 12351 13028 12407 13030
rect 12431 13028 12487 13030
rect 10966 8064 11022 8120
rect 11242 8880 11298 8936
rect 14548 17978 14604 17980
rect 14628 17978 14684 17980
rect 14708 17978 14764 17980
rect 14788 17978 14844 17980
rect 14548 17926 14594 17978
rect 14594 17926 14604 17978
rect 14628 17926 14658 17978
rect 14658 17926 14670 17978
rect 14670 17926 14684 17978
rect 14708 17926 14722 17978
rect 14722 17926 14734 17978
rect 14734 17926 14764 17978
rect 14788 17926 14798 17978
rect 14798 17926 14844 17978
rect 14548 17924 14604 17926
rect 14628 17924 14684 17926
rect 14708 17924 14764 17926
rect 14788 17924 14844 17926
rect 13266 15408 13322 15464
rect 14548 16890 14604 16892
rect 14628 16890 14684 16892
rect 14708 16890 14764 16892
rect 14788 16890 14844 16892
rect 14548 16838 14594 16890
rect 14594 16838 14604 16890
rect 14628 16838 14658 16890
rect 14658 16838 14670 16890
rect 14670 16838 14684 16890
rect 14708 16838 14722 16890
rect 14722 16838 14734 16890
rect 14734 16838 14764 16890
rect 14788 16838 14798 16890
rect 14798 16838 14844 16890
rect 14548 16836 14604 16838
rect 14628 16836 14684 16838
rect 14708 16836 14764 16838
rect 14788 16836 14844 16838
rect 14548 15802 14604 15804
rect 14628 15802 14684 15804
rect 14708 15802 14764 15804
rect 14788 15802 14844 15804
rect 14548 15750 14594 15802
rect 14594 15750 14604 15802
rect 14628 15750 14658 15802
rect 14658 15750 14670 15802
rect 14670 15750 14684 15802
rect 14708 15750 14722 15802
rect 14722 15750 14734 15802
rect 14734 15750 14764 15802
rect 14788 15750 14798 15802
rect 14798 15750 14844 15802
rect 14548 15748 14604 15750
rect 14628 15748 14684 15750
rect 14708 15748 14764 15750
rect 14788 15748 14844 15750
rect 18510 18828 18566 18864
rect 18510 18808 18512 18828
rect 18512 18808 18564 18828
rect 18564 18808 18566 18828
rect 16906 18522 16962 18524
rect 16986 18522 17042 18524
rect 17066 18522 17122 18524
rect 17146 18522 17202 18524
rect 16906 18470 16952 18522
rect 16952 18470 16962 18522
rect 16986 18470 17016 18522
rect 17016 18470 17028 18522
rect 17028 18470 17042 18522
rect 17066 18470 17080 18522
rect 17080 18470 17092 18522
rect 17092 18470 17122 18522
rect 17146 18470 17156 18522
rect 17156 18470 17202 18522
rect 16906 18468 16962 18470
rect 16986 18468 17042 18470
rect 17066 18468 17122 18470
rect 17146 18468 17202 18470
rect 19062 18400 19118 18456
rect 12990 12588 12992 12608
rect 12992 12588 13044 12608
rect 13044 12588 13046 12608
rect 12990 12552 13046 12588
rect 12191 11994 12247 11996
rect 12271 11994 12327 11996
rect 12351 11994 12407 11996
rect 12431 11994 12487 11996
rect 12191 11942 12237 11994
rect 12237 11942 12247 11994
rect 12271 11942 12301 11994
rect 12301 11942 12313 11994
rect 12313 11942 12327 11994
rect 12351 11942 12365 11994
rect 12365 11942 12377 11994
rect 12377 11942 12407 11994
rect 12431 11942 12441 11994
rect 12441 11942 12487 11994
rect 12191 11940 12247 11942
rect 12271 11940 12327 11942
rect 12351 11940 12407 11942
rect 12431 11940 12487 11942
rect 12530 11736 12586 11792
rect 12191 10906 12247 10908
rect 12271 10906 12327 10908
rect 12351 10906 12407 10908
rect 12431 10906 12487 10908
rect 12191 10854 12237 10906
rect 12237 10854 12247 10906
rect 12271 10854 12301 10906
rect 12301 10854 12313 10906
rect 12313 10854 12327 10906
rect 12351 10854 12365 10906
rect 12365 10854 12377 10906
rect 12377 10854 12407 10906
rect 12431 10854 12441 10906
rect 12441 10854 12487 10906
rect 12191 10852 12247 10854
rect 12271 10852 12327 10854
rect 12351 10852 12407 10854
rect 12431 10852 12487 10854
rect 11150 8200 11206 8256
rect 11058 7792 11114 7848
rect 11610 8472 11666 8528
rect 11426 8336 11482 8392
rect 11150 7268 11206 7304
rect 11150 7248 11152 7268
rect 11152 7248 11204 7268
rect 11204 7248 11206 7268
rect 10966 6432 11022 6488
rect 10966 4684 11022 4720
rect 9833 2746 9889 2748
rect 9913 2746 9969 2748
rect 9993 2746 10049 2748
rect 10073 2746 10129 2748
rect 9833 2694 9879 2746
rect 9879 2694 9889 2746
rect 9913 2694 9943 2746
rect 9943 2694 9955 2746
rect 9955 2694 9969 2746
rect 9993 2694 10007 2746
rect 10007 2694 10019 2746
rect 10019 2694 10049 2746
rect 10073 2694 10083 2746
rect 10083 2694 10129 2746
rect 9833 2692 9889 2694
rect 9913 2692 9969 2694
rect 9993 2692 10049 2694
rect 10073 2692 10129 2694
rect 10598 2644 10654 2680
rect 10598 2624 10600 2644
rect 10600 2624 10652 2644
rect 10652 2624 10654 2644
rect 9954 2488 10010 2544
rect 10966 4664 10968 4684
rect 10968 4664 11020 4684
rect 11020 4664 11022 4684
rect 9833 1658 9889 1660
rect 9913 1658 9969 1660
rect 9993 1658 10049 1660
rect 10073 1658 10129 1660
rect 9833 1606 9879 1658
rect 9879 1606 9889 1658
rect 9913 1606 9943 1658
rect 9943 1606 9955 1658
rect 9955 1606 9969 1658
rect 9993 1606 10007 1658
rect 10007 1606 10019 1658
rect 10019 1606 10049 1658
rect 10073 1606 10083 1658
rect 10083 1606 10129 1658
rect 9833 1604 9889 1606
rect 9913 1604 9969 1606
rect 9993 1604 10049 1606
rect 10073 1604 10129 1606
rect 7476 1114 7532 1116
rect 7556 1114 7612 1116
rect 7636 1114 7692 1116
rect 7716 1114 7772 1116
rect 7476 1062 7522 1114
rect 7522 1062 7532 1114
rect 7556 1062 7586 1114
rect 7586 1062 7598 1114
rect 7598 1062 7612 1114
rect 7636 1062 7650 1114
rect 7650 1062 7662 1114
rect 7662 1062 7692 1114
rect 7716 1062 7726 1114
rect 7726 1062 7772 1114
rect 7476 1060 7532 1062
rect 7556 1060 7612 1062
rect 7636 1060 7692 1062
rect 7716 1060 7772 1062
rect 12191 9818 12247 9820
rect 12271 9818 12327 9820
rect 12351 9818 12407 9820
rect 12431 9818 12487 9820
rect 12191 9766 12237 9818
rect 12237 9766 12247 9818
rect 12271 9766 12301 9818
rect 12301 9766 12313 9818
rect 12313 9766 12327 9818
rect 12351 9766 12365 9818
rect 12365 9766 12377 9818
rect 12377 9766 12407 9818
rect 12431 9766 12441 9818
rect 12441 9766 12487 9818
rect 12191 9764 12247 9766
rect 12271 9764 12327 9766
rect 12351 9764 12407 9766
rect 12431 9764 12487 9766
rect 12714 9968 12770 10024
rect 12191 8730 12247 8732
rect 12271 8730 12327 8732
rect 12351 8730 12407 8732
rect 12431 8730 12487 8732
rect 12191 8678 12237 8730
rect 12237 8678 12247 8730
rect 12271 8678 12301 8730
rect 12301 8678 12313 8730
rect 12313 8678 12327 8730
rect 12351 8678 12365 8730
rect 12365 8678 12377 8730
rect 12377 8678 12407 8730
rect 12431 8678 12441 8730
rect 12441 8678 12487 8730
rect 12191 8676 12247 8678
rect 12271 8676 12327 8678
rect 12351 8676 12407 8678
rect 12431 8676 12487 8678
rect 12162 8064 12218 8120
rect 12346 8084 12402 8120
rect 12346 8064 12348 8084
rect 12348 8064 12400 8084
rect 12400 8064 12402 8084
rect 12254 7812 12310 7848
rect 12254 7792 12256 7812
rect 12256 7792 12308 7812
rect 12308 7792 12310 7812
rect 13082 10648 13138 10704
rect 12990 9424 13046 9480
rect 12191 7642 12247 7644
rect 12271 7642 12327 7644
rect 12351 7642 12407 7644
rect 12431 7642 12487 7644
rect 12191 7590 12237 7642
rect 12237 7590 12247 7642
rect 12271 7590 12301 7642
rect 12301 7590 12313 7642
rect 12313 7590 12327 7642
rect 12351 7590 12365 7642
rect 12365 7590 12377 7642
rect 12377 7590 12407 7642
rect 12431 7590 12441 7642
rect 12441 7590 12487 7642
rect 12191 7588 12247 7590
rect 12271 7588 12327 7590
rect 12351 7588 12407 7590
rect 12431 7588 12487 7590
rect 12191 6554 12247 6556
rect 12271 6554 12327 6556
rect 12351 6554 12407 6556
rect 12431 6554 12487 6556
rect 12191 6502 12237 6554
rect 12237 6502 12247 6554
rect 12271 6502 12301 6554
rect 12301 6502 12313 6554
rect 12313 6502 12327 6554
rect 12351 6502 12365 6554
rect 12365 6502 12377 6554
rect 12377 6502 12407 6554
rect 12431 6502 12441 6554
rect 12441 6502 12487 6554
rect 12191 6500 12247 6502
rect 12271 6500 12327 6502
rect 12351 6500 12407 6502
rect 12431 6500 12487 6502
rect 13082 8336 13138 8392
rect 12191 5466 12247 5468
rect 12271 5466 12327 5468
rect 12351 5466 12407 5468
rect 12431 5466 12487 5468
rect 12191 5414 12237 5466
rect 12237 5414 12247 5466
rect 12271 5414 12301 5466
rect 12301 5414 12313 5466
rect 12313 5414 12327 5466
rect 12351 5414 12365 5466
rect 12365 5414 12377 5466
rect 12377 5414 12407 5466
rect 12431 5414 12441 5466
rect 12441 5414 12487 5466
rect 12191 5412 12247 5414
rect 12271 5412 12327 5414
rect 12351 5412 12407 5414
rect 12431 5412 12487 5414
rect 12191 4378 12247 4380
rect 12271 4378 12327 4380
rect 12351 4378 12407 4380
rect 12431 4378 12487 4380
rect 12191 4326 12237 4378
rect 12237 4326 12247 4378
rect 12271 4326 12301 4378
rect 12301 4326 12313 4378
rect 12313 4326 12327 4378
rect 12351 4326 12365 4378
rect 12365 4326 12377 4378
rect 12377 4326 12407 4378
rect 12431 4326 12441 4378
rect 12441 4326 12487 4378
rect 12191 4324 12247 4326
rect 12271 4324 12327 4326
rect 12351 4324 12407 4326
rect 12431 4324 12487 4326
rect 12806 6296 12862 6352
rect 12714 4664 12770 4720
rect 12191 3290 12247 3292
rect 12271 3290 12327 3292
rect 12351 3290 12407 3292
rect 12431 3290 12487 3292
rect 12191 3238 12237 3290
rect 12237 3238 12247 3290
rect 12271 3238 12301 3290
rect 12301 3238 12313 3290
rect 12313 3238 12327 3290
rect 12351 3238 12365 3290
rect 12365 3238 12377 3290
rect 12377 3238 12407 3290
rect 12431 3238 12441 3290
rect 12441 3238 12487 3290
rect 12191 3236 12247 3238
rect 12271 3236 12327 3238
rect 12351 3236 12407 3238
rect 12431 3236 12487 3238
rect 12191 2202 12247 2204
rect 12271 2202 12327 2204
rect 12351 2202 12407 2204
rect 12431 2202 12487 2204
rect 12191 2150 12237 2202
rect 12237 2150 12247 2202
rect 12271 2150 12301 2202
rect 12301 2150 12313 2202
rect 12313 2150 12327 2202
rect 12351 2150 12365 2202
rect 12365 2150 12377 2202
rect 12377 2150 12407 2202
rect 12431 2150 12441 2202
rect 12441 2150 12487 2202
rect 12191 2148 12247 2150
rect 12271 2148 12327 2150
rect 12351 2148 12407 2150
rect 12431 2148 12487 2150
rect 12191 1114 12247 1116
rect 12271 1114 12327 1116
rect 12351 1114 12407 1116
rect 12431 1114 12487 1116
rect 12191 1062 12237 1114
rect 12237 1062 12247 1114
rect 12271 1062 12301 1114
rect 12301 1062 12313 1114
rect 12313 1062 12327 1114
rect 12351 1062 12365 1114
rect 12365 1062 12377 1114
rect 12377 1062 12407 1114
rect 12431 1062 12441 1114
rect 12441 1062 12487 1114
rect 12191 1060 12247 1062
rect 12271 1060 12327 1062
rect 12351 1060 12407 1062
rect 12431 1060 12487 1062
rect 13266 7248 13322 7304
rect 13634 8472 13690 8528
rect 14548 14714 14604 14716
rect 14628 14714 14684 14716
rect 14708 14714 14764 14716
rect 14788 14714 14844 14716
rect 14548 14662 14594 14714
rect 14594 14662 14604 14714
rect 14628 14662 14658 14714
rect 14658 14662 14670 14714
rect 14670 14662 14684 14714
rect 14708 14662 14722 14714
rect 14722 14662 14734 14714
rect 14734 14662 14764 14714
rect 14788 14662 14798 14714
rect 14798 14662 14844 14714
rect 14548 14660 14604 14662
rect 14628 14660 14684 14662
rect 14708 14660 14764 14662
rect 14788 14660 14844 14662
rect 14548 13626 14604 13628
rect 14628 13626 14684 13628
rect 14708 13626 14764 13628
rect 14788 13626 14844 13628
rect 14548 13574 14594 13626
rect 14594 13574 14604 13626
rect 14628 13574 14658 13626
rect 14658 13574 14670 13626
rect 14670 13574 14684 13626
rect 14708 13574 14722 13626
rect 14722 13574 14734 13626
rect 14734 13574 14764 13626
rect 14788 13574 14798 13626
rect 14798 13574 14844 13626
rect 14548 13572 14604 13574
rect 14628 13572 14684 13574
rect 14708 13572 14764 13574
rect 14788 13572 14844 13574
rect 14830 12824 14886 12880
rect 14186 12552 14242 12608
rect 14094 9560 14150 9616
rect 14002 6296 14058 6352
rect 14548 12538 14604 12540
rect 14628 12538 14684 12540
rect 14708 12538 14764 12540
rect 14788 12538 14844 12540
rect 14548 12486 14594 12538
rect 14594 12486 14604 12538
rect 14628 12486 14658 12538
rect 14658 12486 14670 12538
rect 14670 12486 14684 12538
rect 14708 12486 14722 12538
rect 14722 12486 14734 12538
rect 14734 12486 14764 12538
rect 14788 12486 14798 12538
rect 14798 12486 14844 12538
rect 14548 12484 14604 12486
rect 14628 12484 14684 12486
rect 14708 12484 14764 12486
rect 14788 12484 14844 12486
rect 14462 11736 14518 11792
rect 14278 9460 14280 9480
rect 14280 9460 14332 9480
rect 14332 9460 14334 9480
rect 14278 9424 14334 9460
rect 14548 11450 14604 11452
rect 14628 11450 14684 11452
rect 14708 11450 14764 11452
rect 14788 11450 14844 11452
rect 14548 11398 14594 11450
rect 14594 11398 14604 11450
rect 14628 11398 14658 11450
rect 14658 11398 14670 11450
rect 14670 11398 14684 11450
rect 14708 11398 14722 11450
rect 14722 11398 14734 11450
rect 14734 11398 14764 11450
rect 14788 11398 14798 11450
rect 14798 11398 14844 11450
rect 14548 11396 14604 11398
rect 14628 11396 14684 11398
rect 14708 11396 14764 11398
rect 14788 11396 14844 11398
rect 14548 10362 14604 10364
rect 14628 10362 14684 10364
rect 14708 10362 14764 10364
rect 14788 10362 14844 10364
rect 14548 10310 14594 10362
rect 14594 10310 14604 10362
rect 14628 10310 14658 10362
rect 14658 10310 14670 10362
rect 14670 10310 14684 10362
rect 14708 10310 14722 10362
rect 14722 10310 14734 10362
rect 14734 10310 14764 10362
rect 14788 10310 14798 10362
rect 14798 10310 14844 10362
rect 14548 10308 14604 10310
rect 14628 10308 14684 10310
rect 14708 10308 14764 10310
rect 14788 10308 14844 10310
rect 14548 9274 14604 9276
rect 14628 9274 14684 9276
rect 14708 9274 14764 9276
rect 14788 9274 14844 9276
rect 14548 9222 14594 9274
rect 14594 9222 14604 9274
rect 14628 9222 14658 9274
rect 14658 9222 14670 9274
rect 14670 9222 14684 9274
rect 14708 9222 14722 9274
rect 14722 9222 14734 9274
rect 14734 9222 14764 9274
rect 14788 9222 14798 9274
rect 14798 9222 14844 9274
rect 14548 9220 14604 9222
rect 14628 9220 14684 9222
rect 14708 9220 14764 9222
rect 14788 9220 14844 9222
rect 14548 8186 14604 8188
rect 14628 8186 14684 8188
rect 14708 8186 14764 8188
rect 14788 8186 14844 8188
rect 14548 8134 14594 8186
rect 14594 8134 14604 8186
rect 14628 8134 14658 8186
rect 14658 8134 14670 8186
rect 14670 8134 14684 8186
rect 14708 8134 14722 8186
rect 14722 8134 14734 8186
rect 14734 8134 14764 8186
rect 14788 8134 14798 8186
rect 14798 8134 14844 8186
rect 14548 8132 14604 8134
rect 14628 8132 14684 8134
rect 14708 8132 14764 8134
rect 14788 8132 14844 8134
rect 14922 7948 14978 7984
rect 14922 7928 14924 7948
rect 14924 7928 14976 7948
rect 14976 7928 14978 7948
rect 16210 15952 16266 16008
rect 15290 9036 15346 9072
rect 15290 9016 15292 9036
rect 15292 9016 15344 9036
rect 15344 9016 15346 9036
rect 14548 7098 14604 7100
rect 14628 7098 14684 7100
rect 14708 7098 14764 7100
rect 14788 7098 14844 7100
rect 14548 7046 14594 7098
rect 14594 7046 14604 7098
rect 14628 7046 14658 7098
rect 14658 7046 14670 7098
rect 14670 7046 14684 7098
rect 14708 7046 14722 7098
rect 14722 7046 14734 7098
rect 14734 7046 14764 7098
rect 14788 7046 14798 7098
rect 14798 7046 14844 7098
rect 14548 7044 14604 7046
rect 14628 7044 14684 7046
rect 14708 7044 14764 7046
rect 14788 7044 14844 7046
rect 14462 6296 14518 6352
rect 14548 6010 14604 6012
rect 14628 6010 14684 6012
rect 14708 6010 14764 6012
rect 14788 6010 14844 6012
rect 14548 5958 14594 6010
rect 14594 5958 14604 6010
rect 14628 5958 14658 6010
rect 14658 5958 14670 6010
rect 14670 5958 14684 6010
rect 14708 5958 14722 6010
rect 14722 5958 14734 6010
rect 14734 5958 14764 6010
rect 14788 5958 14798 6010
rect 14798 5958 14844 6010
rect 14548 5956 14604 5958
rect 14628 5956 14684 5958
rect 14708 5956 14764 5958
rect 14788 5956 14844 5958
rect 14548 4922 14604 4924
rect 14628 4922 14684 4924
rect 14708 4922 14764 4924
rect 14788 4922 14844 4924
rect 14548 4870 14594 4922
rect 14594 4870 14604 4922
rect 14628 4870 14658 4922
rect 14658 4870 14670 4922
rect 14670 4870 14684 4922
rect 14708 4870 14722 4922
rect 14722 4870 14734 4922
rect 14734 4870 14764 4922
rect 14788 4870 14798 4922
rect 14798 4870 14844 4922
rect 14548 4868 14604 4870
rect 14628 4868 14684 4870
rect 14708 4868 14764 4870
rect 14788 4868 14844 4870
rect 14548 3834 14604 3836
rect 14628 3834 14684 3836
rect 14708 3834 14764 3836
rect 14788 3834 14844 3836
rect 14548 3782 14594 3834
rect 14594 3782 14604 3834
rect 14628 3782 14658 3834
rect 14658 3782 14670 3834
rect 14670 3782 14684 3834
rect 14708 3782 14722 3834
rect 14722 3782 14734 3834
rect 14734 3782 14764 3834
rect 14788 3782 14798 3834
rect 14798 3782 14844 3834
rect 14548 3780 14604 3782
rect 14628 3780 14684 3782
rect 14708 3780 14764 3782
rect 14788 3780 14844 3782
rect 14548 2746 14604 2748
rect 14628 2746 14684 2748
rect 14708 2746 14764 2748
rect 14788 2746 14844 2748
rect 14548 2694 14594 2746
rect 14594 2694 14604 2746
rect 14628 2694 14658 2746
rect 14658 2694 14670 2746
rect 14670 2694 14684 2746
rect 14708 2694 14722 2746
rect 14722 2694 14734 2746
rect 14734 2694 14764 2746
rect 14788 2694 14798 2746
rect 14798 2694 14844 2746
rect 14548 2692 14604 2694
rect 14628 2692 14684 2694
rect 14708 2692 14764 2694
rect 14788 2692 14844 2694
rect 13634 1808 13690 1864
rect 14548 1658 14604 1660
rect 14628 1658 14684 1660
rect 14708 1658 14764 1660
rect 14788 1658 14844 1660
rect 14548 1606 14594 1658
rect 14594 1606 14604 1658
rect 14628 1606 14658 1658
rect 14658 1606 14670 1658
rect 14670 1606 14684 1658
rect 14708 1606 14722 1658
rect 14722 1606 14734 1658
rect 14734 1606 14764 1658
rect 14788 1606 14798 1658
rect 14798 1606 14844 1658
rect 14548 1604 14604 1606
rect 14628 1604 14684 1606
rect 14708 1604 14764 1606
rect 14788 1604 14844 1606
rect 15290 7928 15346 7984
rect 16906 17434 16962 17436
rect 16986 17434 17042 17436
rect 17066 17434 17122 17436
rect 17146 17434 17202 17436
rect 16906 17382 16952 17434
rect 16952 17382 16962 17434
rect 16986 17382 17016 17434
rect 17016 17382 17028 17434
rect 17028 17382 17042 17434
rect 17066 17382 17080 17434
rect 17080 17382 17092 17434
rect 17092 17382 17122 17434
rect 17146 17382 17156 17434
rect 17156 17382 17202 17434
rect 16906 17380 16962 17382
rect 16986 17380 17042 17382
rect 17066 17380 17122 17382
rect 17146 17380 17202 17382
rect 16906 16346 16962 16348
rect 16986 16346 17042 16348
rect 17066 16346 17122 16348
rect 17146 16346 17202 16348
rect 16906 16294 16952 16346
rect 16952 16294 16962 16346
rect 16986 16294 17016 16346
rect 17016 16294 17028 16346
rect 17028 16294 17042 16346
rect 17066 16294 17080 16346
rect 17080 16294 17092 16346
rect 17092 16294 17122 16346
rect 17146 16294 17156 16346
rect 17156 16294 17202 16346
rect 16906 16292 16962 16294
rect 16986 16292 17042 16294
rect 17066 16292 17122 16294
rect 17146 16292 17202 16294
rect 15934 8916 15936 8936
rect 15936 8916 15988 8936
rect 15988 8916 15990 8936
rect 15934 8880 15990 8916
rect 15842 5752 15898 5808
rect 15290 5616 15346 5672
rect 15106 3732 15162 3768
rect 15106 3712 15108 3732
rect 15108 3712 15160 3732
rect 15160 3712 15162 3732
rect 16906 15258 16962 15260
rect 16986 15258 17042 15260
rect 17066 15258 17122 15260
rect 17146 15258 17202 15260
rect 16906 15206 16952 15258
rect 16952 15206 16962 15258
rect 16986 15206 17016 15258
rect 17016 15206 17028 15258
rect 17028 15206 17042 15258
rect 17066 15206 17080 15258
rect 17080 15206 17092 15258
rect 17092 15206 17122 15258
rect 17146 15206 17156 15258
rect 17156 15206 17202 15258
rect 16906 15204 16962 15206
rect 16986 15204 17042 15206
rect 17066 15204 17122 15206
rect 17146 15204 17202 15206
rect 16906 14170 16962 14172
rect 16986 14170 17042 14172
rect 17066 14170 17122 14172
rect 17146 14170 17202 14172
rect 16906 14118 16952 14170
rect 16952 14118 16962 14170
rect 16986 14118 17016 14170
rect 17016 14118 17028 14170
rect 17028 14118 17042 14170
rect 17066 14118 17080 14170
rect 17080 14118 17092 14170
rect 17092 14118 17122 14170
rect 17146 14118 17156 14170
rect 17156 14118 17202 14170
rect 16906 14116 16962 14118
rect 16986 14116 17042 14118
rect 17066 14116 17122 14118
rect 17146 14116 17202 14118
rect 19263 17978 19319 17980
rect 19343 17978 19399 17980
rect 19423 17978 19479 17980
rect 19503 17978 19559 17980
rect 19263 17926 19309 17978
rect 19309 17926 19319 17978
rect 19343 17926 19373 17978
rect 19373 17926 19385 17978
rect 19385 17926 19399 17978
rect 19423 17926 19437 17978
rect 19437 17926 19449 17978
rect 19449 17926 19479 17978
rect 19503 17926 19513 17978
rect 19513 17926 19559 17978
rect 19263 17924 19319 17926
rect 19343 17924 19399 17926
rect 19423 17924 19479 17926
rect 19503 17924 19559 17926
rect 19062 17720 19118 17776
rect 19062 17040 19118 17096
rect 19263 16890 19319 16892
rect 19343 16890 19399 16892
rect 19423 16890 19479 16892
rect 19503 16890 19559 16892
rect 19263 16838 19309 16890
rect 19309 16838 19319 16890
rect 19343 16838 19373 16890
rect 19373 16838 19385 16890
rect 19385 16838 19399 16890
rect 19423 16838 19437 16890
rect 19437 16838 19449 16890
rect 19449 16838 19479 16890
rect 19503 16838 19513 16890
rect 19513 16838 19559 16890
rect 19263 16836 19319 16838
rect 19343 16836 19399 16838
rect 19423 16836 19479 16838
rect 19503 16836 19559 16838
rect 19263 15802 19319 15804
rect 19343 15802 19399 15804
rect 19423 15802 19479 15804
rect 19503 15802 19559 15804
rect 19263 15750 19309 15802
rect 19309 15750 19319 15802
rect 19343 15750 19373 15802
rect 19373 15750 19385 15802
rect 19385 15750 19399 15802
rect 19423 15750 19437 15802
rect 19437 15750 19449 15802
rect 19449 15750 19479 15802
rect 19503 15750 19513 15802
rect 19513 15750 19559 15802
rect 19263 15748 19319 15750
rect 19343 15748 19399 15750
rect 19423 15748 19479 15750
rect 19503 15748 19559 15750
rect 16906 13082 16962 13084
rect 16986 13082 17042 13084
rect 17066 13082 17122 13084
rect 17146 13082 17202 13084
rect 16906 13030 16952 13082
rect 16952 13030 16962 13082
rect 16986 13030 17016 13082
rect 17016 13030 17028 13082
rect 17028 13030 17042 13082
rect 17066 13030 17080 13082
rect 17080 13030 17092 13082
rect 17092 13030 17122 13082
rect 17146 13030 17156 13082
rect 17156 13030 17202 13082
rect 16906 13028 16962 13030
rect 16986 13028 17042 13030
rect 17066 13028 17122 13030
rect 17146 13028 17202 13030
rect 17590 12980 17646 13016
rect 17590 12960 17592 12980
rect 17592 12960 17644 12980
rect 17644 12960 17646 12980
rect 17590 12688 17646 12744
rect 16578 12280 16634 12336
rect 17314 12300 17370 12336
rect 17314 12280 17316 12300
rect 17316 12280 17368 12300
rect 17368 12280 17370 12300
rect 16906 11994 16962 11996
rect 16986 11994 17042 11996
rect 17066 11994 17122 11996
rect 17146 11994 17202 11996
rect 16906 11942 16952 11994
rect 16952 11942 16962 11994
rect 16986 11942 17016 11994
rect 17016 11942 17028 11994
rect 17028 11942 17042 11994
rect 17066 11942 17080 11994
rect 17080 11942 17092 11994
rect 17092 11942 17122 11994
rect 17146 11942 17156 11994
rect 17156 11942 17202 11994
rect 16906 11940 16962 11942
rect 16986 11940 17042 11942
rect 17066 11940 17122 11942
rect 17146 11940 17202 11942
rect 19263 14714 19319 14716
rect 19343 14714 19399 14716
rect 19423 14714 19479 14716
rect 19503 14714 19559 14716
rect 19263 14662 19309 14714
rect 19309 14662 19319 14714
rect 19343 14662 19373 14714
rect 19373 14662 19385 14714
rect 19385 14662 19399 14714
rect 19423 14662 19437 14714
rect 19437 14662 19449 14714
rect 19449 14662 19479 14714
rect 19503 14662 19513 14714
rect 19513 14662 19559 14714
rect 19263 14660 19319 14662
rect 19343 14660 19399 14662
rect 19423 14660 19479 14662
rect 19503 14660 19559 14662
rect 16906 10906 16962 10908
rect 16986 10906 17042 10908
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 16906 10854 16952 10906
rect 16952 10854 16962 10906
rect 16986 10854 17016 10906
rect 17016 10854 17028 10906
rect 17028 10854 17042 10906
rect 17066 10854 17080 10906
rect 17080 10854 17092 10906
rect 17092 10854 17122 10906
rect 17146 10854 17156 10906
rect 17156 10854 17202 10906
rect 16906 10852 16962 10854
rect 16986 10852 17042 10854
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 16670 10512 16726 10568
rect 17314 10004 17316 10024
rect 17316 10004 17368 10024
rect 17368 10004 17370 10024
rect 17314 9968 17370 10004
rect 16906 9818 16962 9820
rect 16986 9818 17042 9820
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 16906 9766 16952 9818
rect 16952 9766 16962 9818
rect 16986 9766 17016 9818
rect 17016 9766 17028 9818
rect 17028 9766 17042 9818
rect 17066 9766 17080 9818
rect 17080 9766 17092 9818
rect 17092 9766 17122 9818
rect 17146 9766 17156 9818
rect 17156 9766 17202 9818
rect 16906 9764 16962 9766
rect 16986 9764 17042 9766
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 16906 8730 16962 8732
rect 16986 8730 17042 8732
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 16906 8678 16952 8730
rect 16952 8678 16962 8730
rect 16986 8678 17016 8730
rect 17016 8678 17028 8730
rect 17028 8678 17042 8730
rect 17066 8678 17080 8730
rect 17080 8678 17092 8730
rect 17092 8678 17122 8730
rect 17146 8678 17156 8730
rect 17156 8678 17202 8730
rect 16906 8676 16962 8678
rect 16986 8676 17042 8678
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 17866 7928 17922 7984
rect 16906 7642 16962 7644
rect 16986 7642 17042 7644
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 16906 7590 16952 7642
rect 16952 7590 16962 7642
rect 16986 7590 17016 7642
rect 17016 7590 17028 7642
rect 17028 7590 17042 7642
rect 17066 7590 17080 7642
rect 17080 7590 17092 7642
rect 17092 7590 17122 7642
rect 17146 7590 17156 7642
rect 17156 7590 17202 7642
rect 16906 7588 16962 7590
rect 16986 7588 17042 7590
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 16906 6554 16962 6556
rect 16986 6554 17042 6556
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 16906 6502 16952 6554
rect 16952 6502 16962 6554
rect 16986 6502 17016 6554
rect 17016 6502 17028 6554
rect 17028 6502 17042 6554
rect 17066 6502 17080 6554
rect 17080 6502 17092 6554
rect 17092 6502 17122 6554
rect 17146 6502 17156 6554
rect 17156 6502 17202 6554
rect 16906 6500 16962 6502
rect 16986 6500 17042 6502
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 17498 6840 17554 6896
rect 16906 5466 16962 5468
rect 16986 5466 17042 5468
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 16906 5414 16952 5466
rect 16952 5414 16962 5466
rect 16986 5414 17016 5466
rect 17016 5414 17028 5466
rect 17028 5414 17042 5466
rect 17066 5414 17080 5466
rect 17080 5414 17092 5466
rect 17092 5414 17122 5466
rect 17146 5414 17156 5466
rect 17156 5414 17202 5466
rect 16906 5412 16962 5414
rect 16986 5412 17042 5414
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 16906 4378 16962 4380
rect 16986 4378 17042 4380
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 16906 4326 16952 4378
rect 16952 4326 16962 4378
rect 16986 4326 17016 4378
rect 17016 4326 17028 4378
rect 17028 4326 17042 4378
rect 17066 4326 17080 4378
rect 17080 4326 17092 4378
rect 17092 4326 17122 4378
rect 17146 4326 17156 4378
rect 17156 4326 17202 4378
rect 16906 4324 16962 4326
rect 16986 4324 17042 4326
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 16762 3732 16818 3768
rect 16762 3712 16764 3732
rect 16764 3712 16816 3732
rect 16816 3712 16818 3732
rect 16906 3290 16962 3292
rect 16986 3290 17042 3292
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 16906 3238 16952 3290
rect 16952 3238 16962 3290
rect 16986 3238 17016 3290
rect 17016 3238 17028 3290
rect 17028 3238 17042 3290
rect 17066 3238 17080 3290
rect 17080 3238 17092 3290
rect 17092 3238 17122 3290
rect 17146 3238 17156 3290
rect 17156 3238 17202 3290
rect 16906 3236 16962 3238
rect 16986 3236 17042 3238
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 16906 2202 16962 2204
rect 16986 2202 17042 2204
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 16906 2150 16952 2202
rect 16952 2150 16962 2202
rect 16986 2150 17016 2202
rect 17016 2150 17028 2202
rect 17028 2150 17042 2202
rect 17066 2150 17080 2202
rect 17080 2150 17092 2202
rect 17092 2150 17122 2202
rect 17146 2150 17156 2202
rect 17156 2150 17202 2202
rect 16906 2148 16962 2150
rect 16986 2148 17042 2150
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 19263 13626 19319 13628
rect 19343 13626 19399 13628
rect 19423 13626 19479 13628
rect 19503 13626 19559 13628
rect 19263 13574 19309 13626
rect 19309 13574 19319 13626
rect 19343 13574 19373 13626
rect 19373 13574 19385 13626
rect 19385 13574 19399 13626
rect 19423 13574 19437 13626
rect 19437 13574 19449 13626
rect 19449 13574 19479 13626
rect 19503 13574 19513 13626
rect 19513 13574 19559 13626
rect 19263 13572 19319 13574
rect 19343 13572 19399 13574
rect 19423 13572 19479 13574
rect 19503 13572 19559 13574
rect 19263 12538 19319 12540
rect 19343 12538 19399 12540
rect 19423 12538 19479 12540
rect 19503 12538 19559 12540
rect 19263 12486 19309 12538
rect 19309 12486 19319 12538
rect 19343 12486 19373 12538
rect 19373 12486 19385 12538
rect 19385 12486 19399 12538
rect 19423 12486 19437 12538
rect 19437 12486 19449 12538
rect 19449 12486 19479 12538
rect 19503 12486 19513 12538
rect 19513 12486 19559 12538
rect 19263 12484 19319 12486
rect 19343 12484 19399 12486
rect 19423 12484 19479 12486
rect 19503 12484 19559 12486
rect 19062 11600 19118 11656
rect 19263 11450 19319 11452
rect 19343 11450 19399 11452
rect 19423 11450 19479 11452
rect 19503 11450 19559 11452
rect 19263 11398 19309 11450
rect 19309 11398 19319 11450
rect 19343 11398 19373 11450
rect 19373 11398 19385 11450
rect 19385 11398 19399 11450
rect 19423 11398 19437 11450
rect 19437 11398 19449 11450
rect 19449 11398 19479 11450
rect 19503 11398 19513 11450
rect 19513 11398 19559 11450
rect 19263 11396 19319 11398
rect 19343 11396 19399 11398
rect 19423 11396 19479 11398
rect 19503 11396 19559 11398
rect 19263 10362 19319 10364
rect 19343 10362 19399 10364
rect 19423 10362 19479 10364
rect 19503 10362 19559 10364
rect 19263 10310 19309 10362
rect 19309 10310 19319 10362
rect 19343 10310 19373 10362
rect 19373 10310 19385 10362
rect 19385 10310 19399 10362
rect 19423 10310 19437 10362
rect 19437 10310 19449 10362
rect 19449 10310 19479 10362
rect 19503 10310 19513 10362
rect 19513 10310 19559 10362
rect 19263 10308 19319 10310
rect 19343 10308 19399 10310
rect 19423 10308 19479 10310
rect 19503 10308 19559 10310
rect 19263 9274 19319 9276
rect 19343 9274 19399 9276
rect 19423 9274 19479 9276
rect 19503 9274 19559 9276
rect 19263 9222 19309 9274
rect 19309 9222 19319 9274
rect 19343 9222 19373 9274
rect 19373 9222 19385 9274
rect 19385 9222 19399 9274
rect 19423 9222 19437 9274
rect 19437 9222 19449 9274
rect 19449 9222 19479 9274
rect 19503 9222 19513 9274
rect 19513 9222 19559 9274
rect 19263 9220 19319 9222
rect 19343 9220 19399 9222
rect 19423 9220 19479 9222
rect 19503 9220 19559 9222
rect 19263 8186 19319 8188
rect 19343 8186 19399 8188
rect 19423 8186 19479 8188
rect 19503 8186 19559 8188
rect 19263 8134 19309 8186
rect 19309 8134 19319 8186
rect 19343 8134 19373 8186
rect 19373 8134 19385 8186
rect 19385 8134 19399 8186
rect 19423 8134 19437 8186
rect 19437 8134 19449 8186
rect 19449 8134 19479 8186
rect 19503 8134 19513 8186
rect 19513 8134 19559 8186
rect 19263 8132 19319 8134
rect 19343 8132 19399 8134
rect 19423 8132 19479 8134
rect 19503 8132 19559 8134
rect 19263 7098 19319 7100
rect 19343 7098 19399 7100
rect 19423 7098 19479 7100
rect 19503 7098 19559 7100
rect 19263 7046 19309 7098
rect 19309 7046 19319 7098
rect 19343 7046 19373 7098
rect 19373 7046 19385 7098
rect 19385 7046 19399 7098
rect 19423 7046 19437 7098
rect 19437 7046 19449 7098
rect 19449 7046 19479 7098
rect 19503 7046 19513 7098
rect 19513 7046 19559 7098
rect 19263 7044 19319 7046
rect 19343 7044 19399 7046
rect 19423 7044 19479 7046
rect 19503 7044 19559 7046
rect 19263 6010 19319 6012
rect 19343 6010 19399 6012
rect 19423 6010 19479 6012
rect 19503 6010 19559 6012
rect 19263 5958 19309 6010
rect 19309 5958 19319 6010
rect 19343 5958 19373 6010
rect 19373 5958 19385 6010
rect 19385 5958 19399 6010
rect 19423 5958 19437 6010
rect 19437 5958 19449 6010
rect 19449 5958 19479 6010
rect 19503 5958 19513 6010
rect 19513 5958 19559 6010
rect 19263 5956 19319 5958
rect 19343 5956 19399 5958
rect 19423 5956 19479 5958
rect 19503 5956 19559 5958
rect 19263 4922 19319 4924
rect 19343 4922 19399 4924
rect 19423 4922 19479 4924
rect 19503 4922 19559 4924
rect 19263 4870 19309 4922
rect 19309 4870 19319 4922
rect 19343 4870 19373 4922
rect 19373 4870 19385 4922
rect 19385 4870 19399 4922
rect 19423 4870 19437 4922
rect 19437 4870 19449 4922
rect 19449 4870 19479 4922
rect 19503 4870 19513 4922
rect 19513 4870 19559 4922
rect 19263 4868 19319 4870
rect 19343 4868 19399 4870
rect 19423 4868 19479 4870
rect 19503 4868 19559 4870
rect 19263 3834 19319 3836
rect 19343 3834 19399 3836
rect 19423 3834 19479 3836
rect 19503 3834 19559 3836
rect 19263 3782 19309 3834
rect 19309 3782 19319 3834
rect 19343 3782 19373 3834
rect 19373 3782 19385 3834
rect 19385 3782 19399 3834
rect 19423 3782 19437 3834
rect 19437 3782 19449 3834
rect 19449 3782 19479 3834
rect 19503 3782 19513 3834
rect 19513 3782 19559 3834
rect 19263 3780 19319 3782
rect 19343 3780 19399 3782
rect 19423 3780 19479 3782
rect 19503 3780 19559 3782
rect 19263 2746 19319 2748
rect 19343 2746 19399 2748
rect 19423 2746 19479 2748
rect 19503 2746 19559 2748
rect 19263 2694 19309 2746
rect 19309 2694 19319 2746
rect 19343 2694 19373 2746
rect 19373 2694 19385 2746
rect 19385 2694 19399 2746
rect 19423 2694 19437 2746
rect 19437 2694 19449 2746
rect 19449 2694 19479 2746
rect 19503 2694 19513 2746
rect 19513 2694 19559 2746
rect 19263 2692 19319 2694
rect 19343 2692 19399 2694
rect 19423 2692 19479 2694
rect 19503 2692 19559 2694
rect 19062 2080 19118 2136
rect 19263 1658 19319 1660
rect 19343 1658 19399 1660
rect 19423 1658 19479 1660
rect 19503 1658 19559 1660
rect 19263 1606 19309 1658
rect 19309 1606 19319 1658
rect 19343 1606 19373 1658
rect 19373 1606 19385 1658
rect 19385 1606 19399 1658
rect 19423 1606 19437 1658
rect 19437 1606 19449 1658
rect 19449 1606 19479 1658
rect 19503 1606 19513 1658
rect 19513 1606 19559 1658
rect 19263 1604 19319 1606
rect 19343 1604 19399 1606
rect 19423 1604 19479 1606
rect 19503 1604 19559 1606
rect 19062 1400 19118 1456
rect 16906 1114 16962 1116
rect 16986 1114 17042 1116
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 16906 1062 16952 1114
rect 16952 1062 16962 1114
rect 16986 1062 17016 1114
rect 17016 1062 17028 1114
rect 17028 1062 17042 1114
rect 17066 1062 17080 1114
rect 17080 1062 17092 1114
rect 17092 1062 17122 1114
rect 17146 1062 17156 1114
rect 17156 1062 17202 1114
rect 16906 1060 16962 1062
rect 16986 1060 17042 1062
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 19062 756 19064 776
rect 19064 756 19116 776
rect 19116 756 19118 776
rect 5118 570 5174 572
rect 5198 570 5254 572
rect 5278 570 5334 572
rect 5358 570 5414 572
rect 5118 518 5164 570
rect 5164 518 5174 570
rect 5198 518 5228 570
rect 5228 518 5240 570
rect 5240 518 5254 570
rect 5278 518 5292 570
rect 5292 518 5304 570
rect 5304 518 5334 570
rect 5358 518 5368 570
rect 5368 518 5414 570
rect 5118 516 5174 518
rect 5198 516 5254 518
rect 5278 516 5334 518
rect 5358 516 5414 518
rect 9833 570 9889 572
rect 9913 570 9969 572
rect 9993 570 10049 572
rect 10073 570 10129 572
rect 9833 518 9879 570
rect 9879 518 9889 570
rect 9913 518 9943 570
rect 9943 518 9955 570
rect 9955 518 9969 570
rect 9993 518 10007 570
rect 10007 518 10019 570
rect 10019 518 10049 570
rect 10073 518 10083 570
rect 10083 518 10129 570
rect 9833 516 9889 518
rect 9913 516 9969 518
rect 9993 516 10049 518
rect 10073 516 10129 518
rect 14548 570 14604 572
rect 14628 570 14684 572
rect 14708 570 14764 572
rect 14788 570 14844 572
rect 14548 518 14594 570
rect 14594 518 14604 570
rect 14628 518 14658 570
rect 14658 518 14670 570
rect 14670 518 14684 570
rect 14708 518 14722 570
rect 14722 518 14734 570
rect 14734 518 14764 570
rect 14788 518 14798 570
rect 14798 518 14844 570
rect 14548 516 14604 518
rect 14628 516 14684 518
rect 14708 516 14764 518
rect 14788 516 14844 518
rect 19062 720 19118 756
rect 19263 570 19319 572
rect 19343 570 19399 572
rect 19423 570 19479 572
rect 19503 570 19559 572
rect 19263 518 19309 570
rect 19309 518 19319 570
rect 19343 518 19373 570
rect 19373 518 19385 570
rect 19385 518 19399 570
rect 19423 518 19437 570
rect 19437 518 19449 570
rect 19449 518 19479 570
rect 19503 518 19513 570
rect 19513 518 19559 570
rect 19263 516 19319 518
rect 19343 516 19399 518
rect 19423 516 19479 518
rect 19503 516 19559 518
rect 18510 40 18566 96
<< metal3 >>
rect 0 19818 400 19848
rect 1117 19818 1183 19821
rect 0 19816 1183 19818
rect 0 19760 1122 19816
rect 1178 19760 1183 19816
rect 0 19758 1183 19760
rect 0 19728 400 19758
rect 1117 19755 1183 19758
rect 0 19138 400 19168
rect 749 19138 815 19141
rect 0 19136 815 19138
rect 0 19080 754 19136
rect 810 19080 815 19136
rect 0 19078 815 19080
rect 0 19048 400 19078
rect 749 19075 815 19078
rect 5108 19072 5424 19073
rect 5108 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5424 19072
rect 5108 19007 5424 19008
rect 9823 19072 10139 19073
rect 9823 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10139 19072
rect 9823 19007 10139 19008
rect 14538 19072 14854 19073
rect 14538 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14854 19072
rect 14538 19007 14854 19008
rect 19253 19072 19569 19073
rect 19253 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19569 19072
rect 19600 19048 20000 19168
rect 19253 19007 19569 19008
rect 18505 18866 18571 18869
rect 19750 18866 19810 19048
rect 18505 18864 19810 18866
rect 18505 18808 18510 18864
rect 18566 18808 19810 18864
rect 18505 18806 19810 18808
rect 18505 18803 18571 18806
rect 2751 18528 3067 18529
rect 0 18458 400 18488
rect 2751 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3067 18528
rect 2751 18463 3067 18464
rect 7466 18528 7782 18529
rect 7466 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7782 18528
rect 7466 18463 7782 18464
rect 12181 18528 12497 18529
rect 12181 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12497 18528
rect 12181 18463 12497 18464
rect 16896 18528 17212 18529
rect 16896 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17212 18528
rect 16896 18463 17212 18464
rect 841 18458 907 18461
rect 0 18456 907 18458
rect 0 18400 846 18456
rect 902 18400 907 18456
rect 0 18398 907 18400
rect 0 18368 400 18398
rect 841 18395 907 18398
rect 19057 18458 19123 18461
rect 19600 18458 20000 18488
rect 19057 18456 20000 18458
rect 19057 18400 19062 18456
rect 19118 18400 20000 18456
rect 19057 18398 20000 18400
rect 19057 18395 19123 18398
rect 19600 18368 20000 18398
rect 5108 17984 5424 17985
rect 5108 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5424 17984
rect 5108 17919 5424 17920
rect 9823 17984 10139 17985
rect 9823 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10139 17984
rect 9823 17919 10139 17920
rect 14538 17984 14854 17985
rect 14538 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14854 17984
rect 14538 17919 14854 17920
rect 19253 17984 19569 17985
rect 19253 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19569 17984
rect 19253 17919 19569 17920
rect 0 17778 400 17808
rect 841 17778 907 17781
rect 0 17776 907 17778
rect 0 17720 846 17776
rect 902 17720 907 17776
rect 0 17718 907 17720
rect 0 17688 400 17718
rect 841 17715 907 17718
rect 19057 17778 19123 17781
rect 19600 17778 20000 17808
rect 19057 17776 20000 17778
rect 19057 17720 19062 17776
rect 19118 17720 20000 17776
rect 19057 17718 20000 17720
rect 19057 17715 19123 17718
rect 19600 17688 20000 17718
rect 2751 17440 3067 17441
rect 2751 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3067 17440
rect 2751 17375 3067 17376
rect 7466 17440 7782 17441
rect 7466 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7782 17440
rect 7466 17375 7782 17376
rect 12181 17440 12497 17441
rect 12181 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12497 17440
rect 12181 17375 12497 17376
rect 16896 17440 17212 17441
rect 16896 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17212 17440
rect 16896 17375 17212 17376
rect 0 17098 400 17128
rect 841 17098 907 17101
rect 0 17096 907 17098
rect 0 17040 846 17096
rect 902 17040 907 17096
rect 0 17038 907 17040
rect 0 17008 400 17038
rect 841 17035 907 17038
rect 19057 17098 19123 17101
rect 19600 17098 20000 17128
rect 19057 17096 20000 17098
rect 19057 17040 19062 17096
rect 19118 17040 20000 17096
rect 19057 17038 20000 17040
rect 19057 17035 19123 17038
rect 19600 17008 20000 17038
rect 5108 16896 5424 16897
rect 5108 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5424 16896
rect 5108 16831 5424 16832
rect 9823 16896 10139 16897
rect 9823 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10139 16896
rect 9823 16831 10139 16832
rect 14538 16896 14854 16897
rect 14538 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14854 16896
rect 14538 16831 14854 16832
rect 19253 16896 19569 16897
rect 19253 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19569 16896
rect 19253 16831 19569 16832
rect 0 16418 400 16448
rect 0 16358 2514 16418
rect 0 16328 400 16358
rect 2454 16146 2514 16358
rect 2751 16352 3067 16353
rect 2751 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3067 16352
rect 2751 16287 3067 16288
rect 7466 16352 7782 16353
rect 7466 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7782 16352
rect 7466 16287 7782 16288
rect 12181 16352 12497 16353
rect 12181 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12497 16352
rect 12181 16287 12497 16288
rect 16896 16352 17212 16353
rect 16896 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17212 16352
rect 16896 16287 17212 16288
rect 3417 16146 3483 16149
rect 2454 16144 3483 16146
rect 2454 16088 3422 16144
rect 3478 16088 3483 16144
rect 2454 16086 3483 16088
rect 3417 16083 3483 16086
rect 11145 16010 11211 16013
rect 16205 16010 16271 16013
rect 11145 16008 16271 16010
rect 11145 15952 11150 16008
rect 11206 15952 16210 16008
rect 16266 15952 16271 16008
rect 11145 15950 16271 15952
rect 11145 15947 11211 15950
rect 16205 15947 16271 15950
rect 5108 15808 5424 15809
rect 5108 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5424 15808
rect 5108 15743 5424 15744
rect 9823 15808 10139 15809
rect 9823 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10139 15808
rect 9823 15743 10139 15744
rect 14538 15808 14854 15809
rect 14538 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14854 15808
rect 14538 15743 14854 15744
rect 19253 15808 19569 15809
rect 19253 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19569 15808
rect 19253 15743 19569 15744
rect 12065 15466 12131 15469
rect 13261 15466 13327 15469
rect 12065 15464 13327 15466
rect 12065 15408 12070 15464
rect 12126 15408 13266 15464
rect 13322 15408 13327 15464
rect 12065 15406 13327 15408
rect 12065 15403 12131 15406
rect 13261 15403 13327 15406
rect 2751 15264 3067 15265
rect 2751 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3067 15264
rect 2751 15199 3067 15200
rect 7466 15264 7782 15265
rect 7466 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7782 15264
rect 7466 15199 7782 15200
rect 12181 15264 12497 15265
rect 12181 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12497 15264
rect 12181 15199 12497 15200
rect 16896 15264 17212 15265
rect 16896 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17212 15264
rect 16896 15199 17212 15200
rect 5108 14720 5424 14721
rect 5108 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5424 14720
rect 5108 14655 5424 14656
rect 9823 14720 10139 14721
rect 9823 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10139 14720
rect 9823 14655 10139 14656
rect 14538 14720 14854 14721
rect 14538 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14854 14720
rect 14538 14655 14854 14656
rect 19253 14720 19569 14721
rect 19253 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19569 14720
rect 19253 14655 19569 14656
rect 2751 14176 3067 14177
rect 2751 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3067 14176
rect 2751 14111 3067 14112
rect 7466 14176 7782 14177
rect 7466 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7782 14176
rect 7466 14111 7782 14112
rect 12181 14176 12497 14177
rect 12181 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12497 14176
rect 12181 14111 12497 14112
rect 16896 14176 17212 14177
rect 16896 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17212 14176
rect 16896 14111 17212 14112
rect 5108 13632 5424 13633
rect 5108 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5424 13632
rect 5108 13567 5424 13568
rect 9823 13632 10139 13633
rect 9823 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10139 13632
rect 9823 13567 10139 13568
rect 14538 13632 14854 13633
rect 14538 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14854 13632
rect 14538 13567 14854 13568
rect 19253 13632 19569 13633
rect 19253 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19569 13632
rect 19253 13567 19569 13568
rect 2751 13088 3067 13089
rect 2751 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3067 13088
rect 2751 13023 3067 13024
rect 7466 13088 7782 13089
rect 7466 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7782 13088
rect 7466 13023 7782 13024
rect 12181 13088 12497 13089
rect 12181 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12497 13088
rect 12181 13023 12497 13024
rect 16896 13088 17212 13089
rect 16896 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17212 13088
rect 16896 13023 17212 13024
rect 17585 13018 17651 13021
rect 19600 13018 20000 13048
rect 17585 13016 20000 13018
rect 17585 12960 17590 13016
rect 17646 12960 20000 13016
rect 17585 12958 20000 12960
rect 17585 12955 17651 12958
rect 19600 12928 20000 12958
rect 10133 12882 10199 12885
rect 14825 12882 14891 12885
rect 10133 12880 14891 12882
rect 10133 12824 10138 12880
rect 10194 12824 14830 12880
rect 14886 12824 14891 12880
rect 10133 12822 14891 12824
rect 10133 12819 10199 12822
rect 14825 12819 14891 12822
rect 8661 12746 8727 12749
rect 17585 12746 17651 12749
rect 8661 12744 17651 12746
rect 8661 12688 8666 12744
rect 8722 12688 17590 12744
rect 17646 12688 17651 12744
rect 8661 12686 17651 12688
rect 8661 12683 8727 12686
rect 17585 12683 17651 12686
rect 10685 12612 10751 12613
rect 10685 12610 10732 12612
rect 10640 12608 10732 12610
rect 10640 12552 10690 12608
rect 10640 12550 10732 12552
rect 10685 12548 10732 12550
rect 10796 12548 10802 12612
rect 12985 12610 13051 12613
rect 14181 12610 14247 12613
rect 12985 12608 14247 12610
rect 12985 12552 12990 12608
rect 13046 12552 14186 12608
rect 14242 12552 14247 12608
rect 12985 12550 14247 12552
rect 10685 12547 10751 12548
rect 12985 12547 13051 12550
rect 14181 12547 14247 12550
rect 5108 12544 5424 12545
rect 5108 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5424 12544
rect 5108 12479 5424 12480
rect 9823 12544 10139 12545
rect 9823 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10139 12544
rect 9823 12479 10139 12480
rect 14538 12544 14854 12545
rect 14538 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14854 12544
rect 14538 12479 14854 12480
rect 19253 12544 19569 12545
rect 19253 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19569 12544
rect 19253 12479 19569 12480
rect 8661 12338 8727 12341
rect 16573 12338 16639 12341
rect 8661 12336 16639 12338
rect 8661 12280 8666 12336
rect 8722 12280 16578 12336
rect 16634 12280 16639 12336
rect 8661 12278 16639 12280
rect 8661 12275 8727 12278
rect 16573 12275 16639 12278
rect 17309 12338 17375 12341
rect 19600 12338 20000 12368
rect 17309 12336 20000 12338
rect 17309 12280 17314 12336
rect 17370 12280 20000 12336
rect 17309 12278 20000 12280
rect 17309 12275 17375 12278
rect 19600 12248 20000 12278
rect 2751 12000 3067 12001
rect 2751 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3067 12000
rect 2751 11935 3067 11936
rect 7466 12000 7782 12001
rect 7466 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7782 12000
rect 7466 11935 7782 11936
rect 12181 12000 12497 12001
rect 12181 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12497 12000
rect 12181 11935 12497 11936
rect 16896 12000 17212 12001
rect 16896 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17212 12000
rect 16896 11935 17212 11936
rect 3601 11794 3667 11797
rect 10317 11794 10383 11797
rect 3601 11792 10383 11794
rect 3601 11736 3606 11792
rect 3662 11736 10322 11792
rect 10378 11736 10383 11792
rect 3601 11734 10383 11736
rect 3601 11731 3667 11734
rect 10317 11731 10383 11734
rect 11697 11794 11763 11797
rect 12525 11794 12591 11797
rect 14457 11794 14523 11797
rect 11697 11792 14523 11794
rect 11697 11736 11702 11792
rect 11758 11736 12530 11792
rect 12586 11736 14462 11792
rect 14518 11736 14523 11792
rect 11697 11734 14523 11736
rect 11697 11731 11763 11734
rect 12525 11731 12591 11734
rect 14457 11731 14523 11734
rect 9622 11596 9628 11660
rect 9692 11658 9698 11660
rect 9765 11658 9831 11661
rect 9692 11656 9831 11658
rect 9692 11600 9770 11656
rect 9826 11600 9831 11656
rect 9692 11598 9831 11600
rect 9692 11596 9698 11598
rect 9765 11595 9831 11598
rect 19057 11658 19123 11661
rect 19600 11658 20000 11688
rect 19057 11656 20000 11658
rect 19057 11600 19062 11656
rect 19118 11600 20000 11656
rect 19057 11598 20000 11600
rect 19057 11595 19123 11598
rect 19600 11568 20000 11598
rect 5108 11456 5424 11457
rect 5108 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5424 11456
rect 5108 11391 5424 11392
rect 9823 11456 10139 11457
rect 9823 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10139 11456
rect 9823 11391 10139 11392
rect 14538 11456 14854 11457
rect 14538 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14854 11456
rect 14538 11391 14854 11392
rect 19253 11456 19569 11457
rect 19253 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19569 11456
rect 19253 11391 19569 11392
rect 19600 10978 20000 11008
rect 17358 10918 20000 10978
rect 2751 10912 3067 10913
rect 2751 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3067 10912
rect 2751 10847 3067 10848
rect 7466 10912 7782 10913
rect 7466 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7782 10912
rect 7466 10847 7782 10848
rect 12181 10912 12497 10913
rect 12181 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12497 10912
rect 12181 10847 12497 10848
rect 16896 10912 17212 10913
rect 16896 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17212 10912
rect 16896 10847 17212 10848
rect 13077 10706 13143 10709
rect 17358 10706 17418 10918
rect 19600 10888 20000 10918
rect 13077 10704 17418 10706
rect 13077 10648 13082 10704
rect 13138 10648 17418 10704
rect 13077 10646 17418 10648
rect 13077 10643 13143 10646
rect 9765 10570 9831 10573
rect 16665 10570 16731 10573
rect 9765 10568 16731 10570
rect 9765 10512 9770 10568
rect 9826 10512 16670 10568
rect 16726 10512 16731 10568
rect 9765 10510 16731 10512
rect 9765 10507 9831 10510
rect 16665 10507 16731 10510
rect 5108 10368 5424 10369
rect 5108 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5424 10368
rect 5108 10303 5424 10304
rect 9823 10368 10139 10369
rect 9823 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10139 10368
rect 9823 10303 10139 10304
rect 14538 10368 14854 10369
rect 14538 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14854 10368
rect 14538 10303 14854 10304
rect 19253 10368 19569 10369
rect 19253 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19569 10368
rect 19253 10303 19569 10304
rect 19600 10208 20000 10328
rect 5717 10026 5783 10029
rect 7557 10026 7623 10029
rect 5717 10024 7623 10026
rect 5717 9968 5722 10024
rect 5778 9968 7562 10024
rect 7618 9968 7623 10024
rect 5717 9966 7623 9968
rect 5717 9963 5783 9966
rect 7557 9963 7623 9966
rect 10685 10026 10751 10029
rect 12709 10026 12775 10029
rect 10685 10024 12775 10026
rect 10685 9968 10690 10024
rect 10746 9968 12714 10024
rect 12770 9968 12775 10024
rect 10685 9966 12775 9968
rect 10685 9963 10751 9966
rect 12709 9963 12775 9966
rect 17309 10026 17375 10029
rect 19934 10026 19994 10208
rect 17309 10024 19994 10026
rect 17309 9968 17314 10024
rect 17370 9968 19994 10024
rect 17309 9966 19994 9968
rect 17309 9963 17375 9966
rect 2751 9824 3067 9825
rect 2751 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3067 9824
rect 2751 9759 3067 9760
rect 7466 9824 7782 9825
rect 7466 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7782 9824
rect 7466 9759 7782 9760
rect 12181 9824 12497 9825
rect 12181 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12497 9824
rect 12181 9759 12497 9760
rect 16896 9824 17212 9825
rect 16896 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17212 9824
rect 16896 9759 17212 9760
rect 11237 9754 11303 9757
rect 11462 9754 11468 9756
rect 11237 9752 11468 9754
rect 11237 9696 11242 9752
rect 11298 9696 11468 9752
rect 11237 9694 11468 9696
rect 11237 9691 11303 9694
rect 11462 9692 11468 9694
rect 11532 9692 11538 9756
rect 14089 9618 14155 9621
rect 19600 9618 20000 9648
rect 14089 9616 20000 9618
rect 14089 9560 14094 9616
rect 14150 9560 20000 9616
rect 14089 9558 20000 9560
rect 14089 9555 14155 9558
rect 19600 9528 20000 9558
rect 5257 9482 5323 9485
rect 7833 9482 7899 9485
rect 5257 9480 7899 9482
rect 5257 9424 5262 9480
rect 5318 9424 7838 9480
rect 7894 9424 7899 9480
rect 5257 9422 7899 9424
rect 5257 9419 5323 9422
rect 7833 9419 7899 9422
rect 10685 9482 10751 9485
rect 12985 9482 13051 9485
rect 14273 9482 14339 9485
rect 10685 9480 14339 9482
rect 10685 9424 10690 9480
rect 10746 9424 12990 9480
rect 13046 9424 14278 9480
rect 14334 9424 14339 9480
rect 10685 9422 14339 9424
rect 10685 9419 10751 9422
rect 12985 9419 13051 9422
rect 14273 9419 14339 9422
rect 5108 9280 5424 9281
rect 5108 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5424 9280
rect 5108 9215 5424 9216
rect 9823 9280 10139 9281
rect 9823 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10139 9280
rect 9823 9215 10139 9216
rect 14538 9280 14854 9281
rect 14538 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14854 9280
rect 14538 9215 14854 9216
rect 19253 9280 19569 9281
rect 19253 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19569 9280
rect 19253 9215 19569 9216
rect 5349 9074 5415 9077
rect 6269 9074 6335 9077
rect 5349 9072 6335 9074
rect 5349 9016 5354 9072
rect 5410 9016 6274 9072
rect 6330 9016 6335 9072
rect 5349 9014 6335 9016
rect 5349 9011 5415 9014
rect 6269 9011 6335 9014
rect 9581 9074 9647 9077
rect 15285 9074 15351 9077
rect 9581 9072 15351 9074
rect 9581 9016 9586 9072
rect 9642 9016 15290 9072
rect 15346 9016 15351 9072
rect 9581 9014 15351 9016
rect 9581 9011 9647 9014
rect 15285 9011 15351 9014
rect 2957 8938 3023 8941
rect 11237 8938 11303 8941
rect 2957 8936 11303 8938
rect 2957 8880 2962 8936
rect 3018 8880 11242 8936
rect 11298 8880 11303 8936
rect 2957 8878 11303 8880
rect 2957 8875 3023 8878
rect 11237 8875 11303 8878
rect 15929 8938 15995 8941
rect 19600 8938 20000 8968
rect 15929 8936 20000 8938
rect 15929 8880 15934 8936
rect 15990 8880 20000 8936
rect 15929 8878 20000 8880
rect 15929 8875 15995 8878
rect 19600 8848 20000 8878
rect 2751 8736 3067 8737
rect 2751 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3067 8736
rect 2751 8671 3067 8672
rect 7466 8736 7782 8737
rect 7466 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7782 8736
rect 7466 8671 7782 8672
rect 12181 8736 12497 8737
rect 12181 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12497 8736
rect 12181 8671 12497 8672
rect 16896 8736 17212 8737
rect 16896 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17212 8736
rect 16896 8671 17212 8672
rect 9765 8530 9831 8533
rect 11605 8530 11671 8533
rect 9765 8528 11671 8530
rect 9765 8472 9770 8528
rect 9826 8472 11610 8528
rect 11666 8472 11671 8528
rect 9765 8470 11671 8472
rect 9765 8467 9831 8470
rect 11605 8467 11671 8470
rect 13629 8528 13695 8533
rect 13629 8472 13634 8528
rect 13690 8472 13695 8528
rect 13629 8467 13695 8472
rect 13770 8470 19994 8530
rect 11421 8394 11487 8397
rect 13077 8394 13143 8397
rect 11421 8392 13143 8394
rect 11421 8336 11426 8392
rect 11482 8336 13082 8392
rect 13138 8336 13143 8392
rect 11421 8334 13143 8336
rect 13632 8394 13692 8467
rect 13770 8394 13830 8470
rect 13632 8334 13830 8394
rect 11421 8331 11487 8334
rect 13077 8331 13143 8334
rect 19934 8288 19994 8470
rect 11145 8260 11211 8261
rect 11094 8258 11100 8260
rect 11054 8198 11100 8258
rect 11164 8256 11211 8260
rect 11206 8200 11211 8256
rect 11094 8196 11100 8198
rect 11164 8196 11211 8200
rect 11145 8195 11211 8196
rect 5108 8192 5424 8193
rect 5108 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5424 8192
rect 5108 8127 5424 8128
rect 9823 8192 10139 8193
rect 9823 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10139 8192
rect 9823 8127 10139 8128
rect 14538 8192 14854 8193
rect 14538 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14854 8192
rect 14538 8127 14854 8128
rect 19253 8192 19569 8193
rect 19253 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19569 8192
rect 19600 8168 20000 8288
rect 19253 8127 19569 8128
rect 10961 8122 11027 8125
rect 12157 8122 12223 8125
rect 10961 8120 12223 8122
rect 10961 8064 10966 8120
rect 11022 8064 12162 8120
rect 12218 8064 12223 8120
rect 10961 8062 12223 8064
rect 10961 8059 11027 8062
rect 12157 8059 12223 8062
rect 12341 8122 12407 8125
rect 12341 8120 13692 8122
rect 12341 8064 12346 8120
rect 12402 8064 13692 8120
rect 12341 8062 13692 8064
rect 12341 8059 12407 8062
rect 13632 7986 13692 8062
rect 14917 7986 14983 7989
rect 15285 7986 15351 7989
rect 17861 7986 17927 7989
rect 13632 7984 17927 7986
rect 13632 7928 14922 7984
rect 14978 7928 15290 7984
rect 15346 7928 17866 7984
rect 17922 7928 17927 7984
rect 13632 7926 17927 7928
rect 14917 7923 14983 7926
rect 15285 7923 15351 7926
rect 17861 7923 17927 7926
rect 11053 7850 11119 7853
rect 12249 7850 12315 7853
rect 11053 7848 12315 7850
rect 11053 7792 11058 7848
rect 11114 7792 12254 7848
rect 12310 7792 12315 7848
rect 11053 7790 12315 7792
rect 11053 7787 11119 7790
rect 12249 7787 12315 7790
rect 2751 7648 3067 7649
rect 2751 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3067 7648
rect 2751 7583 3067 7584
rect 7466 7648 7782 7649
rect 7466 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7782 7648
rect 7466 7583 7782 7584
rect 12181 7648 12497 7649
rect 12181 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12497 7648
rect 12181 7583 12497 7584
rect 16896 7648 17212 7649
rect 16896 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17212 7648
rect 16896 7583 17212 7584
rect 9029 7306 9095 7309
rect 9581 7306 9647 7309
rect 9029 7304 9647 7306
rect 9029 7248 9034 7304
rect 9090 7248 9586 7304
rect 9642 7248 9647 7304
rect 9029 7246 9647 7248
rect 9029 7243 9095 7246
rect 9581 7243 9647 7246
rect 11145 7306 11211 7309
rect 13261 7306 13327 7309
rect 11145 7304 13327 7306
rect 11145 7248 11150 7304
rect 11206 7248 13266 7304
rect 13322 7248 13327 7304
rect 11145 7246 13327 7248
rect 11145 7243 11211 7246
rect 13261 7243 13327 7246
rect 5108 7104 5424 7105
rect 5108 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5424 7104
rect 5108 7039 5424 7040
rect 9823 7104 10139 7105
rect 9823 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10139 7104
rect 9823 7039 10139 7040
rect 14538 7104 14854 7105
rect 14538 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14854 7104
rect 14538 7039 14854 7040
rect 19253 7104 19569 7105
rect 19253 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19569 7104
rect 19253 7039 19569 7040
rect 9121 7034 9187 7037
rect 9489 7034 9555 7037
rect 9121 7032 9555 7034
rect 9121 6976 9126 7032
rect 9182 6976 9494 7032
rect 9550 6976 9555 7032
rect 9121 6974 9555 6976
rect 9121 6971 9187 6974
rect 9489 6971 9555 6974
rect 9581 6898 9647 6901
rect 17493 6898 17559 6901
rect 9581 6896 17559 6898
rect 9581 6840 9586 6896
rect 9642 6840 17498 6896
rect 17554 6840 17559 6896
rect 9581 6838 17559 6840
rect 9581 6835 9647 6838
rect 17493 6835 17559 6838
rect 11094 6700 11100 6764
rect 11164 6700 11170 6764
rect 2751 6560 3067 6561
rect 2751 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3067 6560
rect 2751 6495 3067 6496
rect 7466 6560 7782 6561
rect 7466 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7782 6560
rect 7466 6495 7782 6496
rect 10961 6490 11027 6493
rect 11102 6490 11162 6700
rect 12181 6560 12497 6561
rect 12181 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12497 6560
rect 12181 6495 12497 6496
rect 16896 6560 17212 6561
rect 16896 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17212 6560
rect 16896 6495 17212 6496
rect 10961 6488 11162 6490
rect 10961 6432 10966 6488
rect 11022 6432 11162 6488
rect 10961 6430 11162 6432
rect 10961 6427 11027 6430
rect 7281 6354 7347 6357
rect 12801 6354 12867 6357
rect 7281 6352 12867 6354
rect 7281 6296 7286 6352
rect 7342 6296 12806 6352
rect 12862 6296 12867 6352
rect 7281 6294 12867 6296
rect 7281 6291 7347 6294
rect 12801 6291 12867 6294
rect 13997 6354 14063 6357
rect 14457 6354 14523 6357
rect 13997 6352 14523 6354
rect 13997 6296 14002 6352
rect 14058 6296 14462 6352
rect 14518 6296 14523 6352
rect 13997 6294 14523 6296
rect 13997 6291 14063 6294
rect 14457 6291 14523 6294
rect 5108 6016 5424 6017
rect 5108 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5424 6016
rect 5108 5951 5424 5952
rect 9823 6016 10139 6017
rect 9823 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10139 6016
rect 9823 5951 10139 5952
rect 14538 6016 14854 6017
rect 14538 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14854 6016
rect 14538 5951 14854 5952
rect 19253 6016 19569 6017
rect 19253 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19569 6016
rect 19253 5951 19569 5952
rect 8845 5810 8911 5813
rect 9397 5810 9463 5813
rect 8845 5808 9463 5810
rect 8845 5752 8850 5808
rect 8906 5752 9402 5808
rect 9458 5752 9463 5808
rect 8845 5750 9463 5752
rect 8845 5747 8911 5750
rect 9397 5747 9463 5750
rect 10777 5810 10843 5813
rect 15837 5810 15903 5813
rect 10777 5808 15903 5810
rect 10777 5752 10782 5808
rect 10838 5752 15842 5808
rect 15898 5752 15903 5808
rect 10777 5750 15903 5752
rect 10777 5747 10843 5750
rect 15837 5747 15903 5750
rect 9029 5674 9095 5677
rect 9305 5674 9371 5677
rect 9029 5672 9371 5674
rect 9029 5616 9034 5672
rect 9090 5616 9310 5672
rect 9366 5616 9371 5672
rect 9029 5614 9371 5616
rect 9029 5611 9095 5614
rect 9305 5611 9371 5614
rect 9673 5674 9739 5677
rect 15285 5674 15351 5677
rect 9673 5672 15351 5674
rect 9673 5616 9678 5672
rect 9734 5616 15290 5672
rect 15346 5616 15351 5672
rect 9673 5614 15351 5616
rect 9673 5611 9739 5614
rect 15285 5611 15351 5614
rect 2751 5472 3067 5473
rect 2751 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3067 5472
rect 2751 5407 3067 5408
rect 7466 5472 7782 5473
rect 7466 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7782 5472
rect 7466 5407 7782 5408
rect 12181 5472 12497 5473
rect 12181 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12497 5472
rect 12181 5407 12497 5408
rect 16896 5472 17212 5473
rect 16896 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17212 5472
rect 16896 5407 17212 5408
rect 3049 5130 3115 5133
rect 9622 5130 9628 5132
rect 3049 5128 9628 5130
rect 3049 5072 3054 5128
rect 3110 5072 9628 5128
rect 3049 5070 9628 5072
rect 3049 5067 3115 5070
rect 9622 5068 9628 5070
rect 9692 5068 9698 5132
rect 5108 4928 5424 4929
rect 5108 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5424 4928
rect 5108 4863 5424 4864
rect 9823 4928 10139 4929
rect 9823 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10139 4928
rect 9823 4863 10139 4864
rect 14538 4928 14854 4929
rect 14538 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14854 4928
rect 14538 4863 14854 4864
rect 19253 4928 19569 4929
rect 19253 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19569 4928
rect 19253 4863 19569 4864
rect 10961 4722 11027 4725
rect 12709 4722 12775 4725
rect 10961 4720 12775 4722
rect 10961 4664 10966 4720
rect 11022 4664 12714 4720
rect 12770 4664 12775 4720
rect 10961 4662 12775 4664
rect 10961 4659 11027 4662
rect 12709 4659 12775 4662
rect 2751 4384 3067 4385
rect 2751 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3067 4384
rect 2751 4319 3067 4320
rect 7466 4384 7782 4385
rect 7466 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7782 4384
rect 7466 4319 7782 4320
rect 12181 4384 12497 4385
rect 12181 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12497 4384
rect 12181 4319 12497 4320
rect 16896 4384 17212 4385
rect 16896 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17212 4384
rect 16896 4319 17212 4320
rect 5108 3840 5424 3841
rect 5108 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5424 3840
rect 5108 3775 5424 3776
rect 9823 3840 10139 3841
rect 9823 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10139 3840
rect 9823 3775 10139 3776
rect 14538 3840 14854 3841
rect 14538 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14854 3840
rect 14538 3775 14854 3776
rect 19253 3840 19569 3841
rect 19253 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19569 3840
rect 19253 3775 19569 3776
rect 15101 3770 15167 3773
rect 16757 3770 16823 3773
rect 15101 3768 16823 3770
rect 15101 3712 15106 3768
rect 15162 3712 16762 3768
rect 16818 3712 16823 3768
rect 15101 3710 16823 3712
rect 15101 3707 15167 3710
rect 16757 3707 16823 3710
rect 2751 3296 3067 3297
rect 2751 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3067 3296
rect 2751 3231 3067 3232
rect 7466 3296 7782 3297
rect 7466 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7782 3296
rect 7466 3231 7782 3232
rect 12181 3296 12497 3297
rect 12181 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12497 3296
rect 12181 3231 12497 3232
rect 16896 3296 17212 3297
rect 16896 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17212 3296
rect 16896 3231 17212 3232
rect 5108 2752 5424 2753
rect 5108 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5424 2752
rect 5108 2687 5424 2688
rect 9823 2752 10139 2753
rect 9823 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10139 2752
rect 9823 2687 10139 2688
rect 14538 2752 14854 2753
rect 14538 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14854 2752
rect 14538 2687 14854 2688
rect 19253 2752 19569 2753
rect 19253 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19569 2752
rect 19253 2687 19569 2688
rect 10593 2682 10659 2685
rect 10726 2682 10732 2684
rect 10593 2680 10732 2682
rect 10593 2624 10598 2680
rect 10654 2624 10732 2680
rect 10593 2622 10732 2624
rect 10593 2619 10659 2622
rect 10726 2620 10732 2622
rect 10796 2620 10802 2684
rect 11462 2620 11468 2684
rect 11532 2620 11538 2684
rect 9949 2546 10015 2549
rect 11470 2546 11530 2620
rect 9949 2544 11530 2546
rect 9949 2488 9954 2544
rect 10010 2488 11530 2544
rect 9949 2486 11530 2488
rect 9949 2483 10015 2486
rect 2751 2208 3067 2209
rect 2751 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3067 2208
rect 2751 2143 3067 2144
rect 7466 2208 7782 2209
rect 7466 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7782 2208
rect 7466 2143 7782 2144
rect 12181 2208 12497 2209
rect 12181 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12497 2208
rect 12181 2143 12497 2144
rect 16896 2208 17212 2209
rect 16896 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17212 2208
rect 16896 2143 17212 2144
rect 19057 2138 19123 2141
rect 19600 2138 20000 2168
rect 19057 2136 20000 2138
rect 19057 2080 19062 2136
rect 19118 2080 20000 2136
rect 19057 2078 20000 2080
rect 19057 2075 19123 2078
rect 19600 2048 20000 2078
rect 4797 1866 4863 1869
rect 13629 1866 13695 1869
rect 4797 1864 13695 1866
rect 4797 1808 4802 1864
rect 4858 1808 13634 1864
rect 13690 1808 13695 1864
rect 4797 1806 13695 1808
rect 4797 1803 4863 1806
rect 13629 1803 13695 1806
rect 5108 1664 5424 1665
rect 5108 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5424 1664
rect 5108 1599 5424 1600
rect 9823 1664 10139 1665
rect 9823 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10139 1664
rect 9823 1599 10139 1600
rect 14538 1664 14854 1665
rect 14538 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14854 1664
rect 14538 1599 14854 1600
rect 19253 1664 19569 1665
rect 19253 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19569 1664
rect 19253 1599 19569 1600
rect 19057 1458 19123 1461
rect 19600 1458 20000 1488
rect 19057 1456 20000 1458
rect 19057 1400 19062 1456
rect 19118 1400 20000 1456
rect 19057 1398 20000 1400
rect 19057 1395 19123 1398
rect 19600 1368 20000 1398
rect 2751 1120 3067 1121
rect 2751 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3067 1120
rect 2751 1055 3067 1056
rect 7466 1120 7782 1121
rect 7466 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7782 1120
rect 7466 1055 7782 1056
rect 12181 1120 12497 1121
rect 12181 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12497 1120
rect 12181 1055 12497 1056
rect 16896 1120 17212 1121
rect 16896 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17212 1120
rect 16896 1055 17212 1056
rect 19057 778 19123 781
rect 19600 778 20000 808
rect 19057 776 20000 778
rect 19057 720 19062 776
rect 19118 720 20000 776
rect 19057 718 20000 720
rect 19057 715 19123 718
rect 19600 688 20000 718
rect 5108 576 5424 577
rect 5108 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5424 576
rect 5108 511 5424 512
rect 9823 576 10139 577
rect 9823 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10139 576
rect 9823 511 10139 512
rect 14538 576 14854 577
rect 14538 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14854 576
rect 14538 511 14854 512
rect 19253 576 19569 577
rect 19253 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19569 576
rect 19253 511 19569 512
rect 18505 98 18571 101
rect 19600 98 20000 128
rect 18505 96 20000 98
rect 18505 40 18510 96
rect 18566 40 20000 96
rect 18505 38 20000 40
rect 18505 35 18571 38
rect 19600 8 20000 38
<< via3 >>
rect 5114 19068 5178 19072
rect 5114 19012 5118 19068
rect 5118 19012 5174 19068
rect 5174 19012 5178 19068
rect 5114 19008 5178 19012
rect 5194 19068 5258 19072
rect 5194 19012 5198 19068
rect 5198 19012 5254 19068
rect 5254 19012 5258 19068
rect 5194 19008 5258 19012
rect 5274 19068 5338 19072
rect 5274 19012 5278 19068
rect 5278 19012 5334 19068
rect 5334 19012 5338 19068
rect 5274 19008 5338 19012
rect 5354 19068 5418 19072
rect 5354 19012 5358 19068
rect 5358 19012 5414 19068
rect 5414 19012 5418 19068
rect 5354 19008 5418 19012
rect 9829 19068 9893 19072
rect 9829 19012 9833 19068
rect 9833 19012 9889 19068
rect 9889 19012 9893 19068
rect 9829 19008 9893 19012
rect 9909 19068 9973 19072
rect 9909 19012 9913 19068
rect 9913 19012 9969 19068
rect 9969 19012 9973 19068
rect 9909 19008 9973 19012
rect 9989 19068 10053 19072
rect 9989 19012 9993 19068
rect 9993 19012 10049 19068
rect 10049 19012 10053 19068
rect 9989 19008 10053 19012
rect 10069 19068 10133 19072
rect 10069 19012 10073 19068
rect 10073 19012 10129 19068
rect 10129 19012 10133 19068
rect 10069 19008 10133 19012
rect 14544 19068 14608 19072
rect 14544 19012 14548 19068
rect 14548 19012 14604 19068
rect 14604 19012 14608 19068
rect 14544 19008 14608 19012
rect 14624 19068 14688 19072
rect 14624 19012 14628 19068
rect 14628 19012 14684 19068
rect 14684 19012 14688 19068
rect 14624 19008 14688 19012
rect 14704 19068 14768 19072
rect 14704 19012 14708 19068
rect 14708 19012 14764 19068
rect 14764 19012 14768 19068
rect 14704 19008 14768 19012
rect 14784 19068 14848 19072
rect 14784 19012 14788 19068
rect 14788 19012 14844 19068
rect 14844 19012 14848 19068
rect 14784 19008 14848 19012
rect 19259 19068 19323 19072
rect 19259 19012 19263 19068
rect 19263 19012 19319 19068
rect 19319 19012 19323 19068
rect 19259 19008 19323 19012
rect 19339 19068 19403 19072
rect 19339 19012 19343 19068
rect 19343 19012 19399 19068
rect 19399 19012 19403 19068
rect 19339 19008 19403 19012
rect 19419 19068 19483 19072
rect 19419 19012 19423 19068
rect 19423 19012 19479 19068
rect 19479 19012 19483 19068
rect 19419 19008 19483 19012
rect 19499 19068 19563 19072
rect 19499 19012 19503 19068
rect 19503 19012 19559 19068
rect 19559 19012 19563 19068
rect 19499 19008 19563 19012
rect 2757 18524 2821 18528
rect 2757 18468 2761 18524
rect 2761 18468 2817 18524
rect 2817 18468 2821 18524
rect 2757 18464 2821 18468
rect 2837 18524 2901 18528
rect 2837 18468 2841 18524
rect 2841 18468 2897 18524
rect 2897 18468 2901 18524
rect 2837 18464 2901 18468
rect 2917 18524 2981 18528
rect 2917 18468 2921 18524
rect 2921 18468 2977 18524
rect 2977 18468 2981 18524
rect 2917 18464 2981 18468
rect 2997 18524 3061 18528
rect 2997 18468 3001 18524
rect 3001 18468 3057 18524
rect 3057 18468 3061 18524
rect 2997 18464 3061 18468
rect 7472 18524 7536 18528
rect 7472 18468 7476 18524
rect 7476 18468 7532 18524
rect 7532 18468 7536 18524
rect 7472 18464 7536 18468
rect 7552 18524 7616 18528
rect 7552 18468 7556 18524
rect 7556 18468 7612 18524
rect 7612 18468 7616 18524
rect 7552 18464 7616 18468
rect 7632 18524 7696 18528
rect 7632 18468 7636 18524
rect 7636 18468 7692 18524
rect 7692 18468 7696 18524
rect 7632 18464 7696 18468
rect 7712 18524 7776 18528
rect 7712 18468 7716 18524
rect 7716 18468 7772 18524
rect 7772 18468 7776 18524
rect 7712 18464 7776 18468
rect 12187 18524 12251 18528
rect 12187 18468 12191 18524
rect 12191 18468 12247 18524
rect 12247 18468 12251 18524
rect 12187 18464 12251 18468
rect 12267 18524 12331 18528
rect 12267 18468 12271 18524
rect 12271 18468 12327 18524
rect 12327 18468 12331 18524
rect 12267 18464 12331 18468
rect 12347 18524 12411 18528
rect 12347 18468 12351 18524
rect 12351 18468 12407 18524
rect 12407 18468 12411 18524
rect 12347 18464 12411 18468
rect 12427 18524 12491 18528
rect 12427 18468 12431 18524
rect 12431 18468 12487 18524
rect 12487 18468 12491 18524
rect 12427 18464 12491 18468
rect 16902 18524 16966 18528
rect 16902 18468 16906 18524
rect 16906 18468 16962 18524
rect 16962 18468 16966 18524
rect 16902 18464 16966 18468
rect 16982 18524 17046 18528
rect 16982 18468 16986 18524
rect 16986 18468 17042 18524
rect 17042 18468 17046 18524
rect 16982 18464 17046 18468
rect 17062 18524 17126 18528
rect 17062 18468 17066 18524
rect 17066 18468 17122 18524
rect 17122 18468 17126 18524
rect 17062 18464 17126 18468
rect 17142 18524 17206 18528
rect 17142 18468 17146 18524
rect 17146 18468 17202 18524
rect 17202 18468 17206 18524
rect 17142 18464 17206 18468
rect 5114 17980 5178 17984
rect 5114 17924 5118 17980
rect 5118 17924 5174 17980
rect 5174 17924 5178 17980
rect 5114 17920 5178 17924
rect 5194 17980 5258 17984
rect 5194 17924 5198 17980
rect 5198 17924 5254 17980
rect 5254 17924 5258 17980
rect 5194 17920 5258 17924
rect 5274 17980 5338 17984
rect 5274 17924 5278 17980
rect 5278 17924 5334 17980
rect 5334 17924 5338 17980
rect 5274 17920 5338 17924
rect 5354 17980 5418 17984
rect 5354 17924 5358 17980
rect 5358 17924 5414 17980
rect 5414 17924 5418 17980
rect 5354 17920 5418 17924
rect 9829 17980 9893 17984
rect 9829 17924 9833 17980
rect 9833 17924 9889 17980
rect 9889 17924 9893 17980
rect 9829 17920 9893 17924
rect 9909 17980 9973 17984
rect 9909 17924 9913 17980
rect 9913 17924 9969 17980
rect 9969 17924 9973 17980
rect 9909 17920 9973 17924
rect 9989 17980 10053 17984
rect 9989 17924 9993 17980
rect 9993 17924 10049 17980
rect 10049 17924 10053 17980
rect 9989 17920 10053 17924
rect 10069 17980 10133 17984
rect 10069 17924 10073 17980
rect 10073 17924 10129 17980
rect 10129 17924 10133 17980
rect 10069 17920 10133 17924
rect 14544 17980 14608 17984
rect 14544 17924 14548 17980
rect 14548 17924 14604 17980
rect 14604 17924 14608 17980
rect 14544 17920 14608 17924
rect 14624 17980 14688 17984
rect 14624 17924 14628 17980
rect 14628 17924 14684 17980
rect 14684 17924 14688 17980
rect 14624 17920 14688 17924
rect 14704 17980 14768 17984
rect 14704 17924 14708 17980
rect 14708 17924 14764 17980
rect 14764 17924 14768 17980
rect 14704 17920 14768 17924
rect 14784 17980 14848 17984
rect 14784 17924 14788 17980
rect 14788 17924 14844 17980
rect 14844 17924 14848 17980
rect 14784 17920 14848 17924
rect 19259 17980 19323 17984
rect 19259 17924 19263 17980
rect 19263 17924 19319 17980
rect 19319 17924 19323 17980
rect 19259 17920 19323 17924
rect 19339 17980 19403 17984
rect 19339 17924 19343 17980
rect 19343 17924 19399 17980
rect 19399 17924 19403 17980
rect 19339 17920 19403 17924
rect 19419 17980 19483 17984
rect 19419 17924 19423 17980
rect 19423 17924 19479 17980
rect 19479 17924 19483 17980
rect 19419 17920 19483 17924
rect 19499 17980 19563 17984
rect 19499 17924 19503 17980
rect 19503 17924 19559 17980
rect 19559 17924 19563 17980
rect 19499 17920 19563 17924
rect 2757 17436 2821 17440
rect 2757 17380 2761 17436
rect 2761 17380 2817 17436
rect 2817 17380 2821 17436
rect 2757 17376 2821 17380
rect 2837 17436 2901 17440
rect 2837 17380 2841 17436
rect 2841 17380 2897 17436
rect 2897 17380 2901 17436
rect 2837 17376 2901 17380
rect 2917 17436 2981 17440
rect 2917 17380 2921 17436
rect 2921 17380 2977 17436
rect 2977 17380 2981 17436
rect 2917 17376 2981 17380
rect 2997 17436 3061 17440
rect 2997 17380 3001 17436
rect 3001 17380 3057 17436
rect 3057 17380 3061 17436
rect 2997 17376 3061 17380
rect 7472 17436 7536 17440
rect 7472 17380 7476 17436
rect 7476 17380 7532 17436
rect 7532 17380 7536 17436
rect 7472 17376 7536 17380
rect 7552 17436 7616 17440
rect 7552 17380 7556 17436
rect 7556 17380 7612 17436
rect 7612 17380 7616 17436
rect 7552 17376 7616 17380
rect 7632 17436 7696 17440
rect 7632 17380 7636 17436
rect 7636 17380 7692 17436
rect 7692 17380 7696 17436
rect 7632 17376 7696 17380
rect 7712 17436 7776 17440
rect 7712 17380 7716 17436
rect 7716 17380 7772 17436
rect 7772 17380 7776 17436
rect 7712 17376 7776 17380
rect 12187 17436 12251 17440
rect 12187 17380 12191 17436
rect 12191 17380 12247 17436
rect 12247 17380 12251 17436
rect 12187 17376 12251 17380
rect 12267 17436 12331 17440
rect 12267 17380 12271 17436
rect 12271 17380 12327 17436
rect 12327 17380 12331 17436
rect 12267 17376 12331 17380
rect 12347 17436 12411 17440
rect 12347 17380 12351 17436
rect 12351 17380 12407 17436
rect 12407 17380 12411 17436
rect 12347 17376 12411 17380
rect 12427 17436 12491 17440
rect 12427 17380 12431 17436
rect 12431 17380 12487 17436
rect 12487 17380 12491 17436
rect 12427 17376 12491 17380
rect 16902 17436 16966 17440
rect 16902 17380 16906 17436
rect 16906 17380 16962 17436
rect 16962 17380 16966 17436
rect 16902 17376 16966 17380
rect 16982 17436 17046 17440
rect 16982 17380 16986 17436
rect 16986 17380 17042 17436
rect 17042 17380 17046 17436
rect 16982 17376 17046 17380
rect 17062 17436 17126 17440
rect 17062 17380 17066 17436
rect 17066 17380 17122 17436
rect 17122 17380 17126 17436
rect 17062 17376 17126 17380
rect 17142 17436 17206 17440
rect 17142 17380 17146 17436
rect 17146 17380 17202 17436
rect 17202 17380 17206 17436
rect 17142 17376 17206 17380
rect 5114 16892 5178 16896
rect 5114 16836 5118 16892
rect 5118 16836 5174 16892
rect 5174 16836 5178 16892
rect 5114 16832 5178 16836
rect 5194 16892 5258 16896
rect 5194 16836 5198 16892
rect 5198 16836 5254 16892
rect 5254 16836 5258 16892
rect 5194 16832 5258 16836
rect 5274 16892 5338 16896
rect 5274 16836 5278 16892
rect 5278 16836 5334 16892
rect 5334 16836 5338 16892
rect 5274 16832 5338 16836
rect 5354 16892 5418 16896
rect 5354 16836 5358 16892
rect 5358 16836 5414 16892
rect 5414 16836 5418 16892
rect 5354 16832 5418 16836
rect 9829 16892 9893 16896
rect 9829 16836 9833 16892
rect 9833 16836 9889 16892
rect 9889 16836 9893 16892
rect 9829 16832 9893 16836
rect 9909 16892 9973 16896
rect 9909 16836 9913 16892
rect 9913 16836 9969 16892
rect 9969 16836 9973 16892
rect 9909 16832 9973 16836
rect 9989 16892 10053 16896
rect 9989 16836 9993 16892
rect 9993 16836 10049 16892
rect 10049 16836 10053 16892
rect 9989 16832 10053 16836
rect 10069 16892 10133 16896
rect 10069 16836 10073 16892
rect 10073 16836 10129 16892
rect 10129 16836 10133 16892
rect 10069 16832 10133 16836
rect 14544 16892 14608 16896
rect 14544 16836 14548 16892
rect 14548 16836 14604 16892
rect 14604 16836 14608 16892
rect 14544 16832 14608 16836
rect 14624 16892 14688 16896
rect 14624 16836 14628 16892
rect 14628 16836 14684 16892
rect 14684 16836 14688 16892
rect 14624 16832 14688 16836
rect 14704 16892 14768 16896
rect 14704 16836 14708 16892
rect 14708 16836 14764 16892
rect 14764 16836 14768 16892
rect 14704 16832 14768 16836
rect 14784 16892 14848 16896
rect 14784 16836 14788 16892
rect 14788 16836 14844 16892
rect 14844 16836 14848 16892
rect 14784 16832 14848 16836
rect 19259 16892 19323 16896
rect 19259 16836 19263 16892
rect 19263 16836 19319 16892
rect 19319 16836 19323 16892
rect 19259 16832 19323 16836
rect 19339 16892 19403 16896
rect 19339 16836 19343 16892
rect 19343 16836 19399 16892
rect 19399 16836 19403 16892
rect 19339 16832 19403 16836
rect 19419 16892 19483 16896
rect 19419 16836 19423 16892
rect 19423 16836 19479 16892
rect 19479 16836 19483 16892
rect 19419 16832 19483 16836
rect 19499 16892 19563 16896
rect 19499 16836 19503 16892
rect 19503 16836 19559 16892
rect 19559 16836 19563 16892
rect 19499 16832 19563 16836
rect 2757 16348 2821 16352
rect 2757 16292 2761 16348
rect 2761 16292 2817 16348
rect 2817 16292 2821 16348
rect 2757 16288 2821 16292
rect 2837 16348 2901 16352
rect 2837 16292 2841 16348
rect 2841 16292 2897 16348
rect 2897 16292 2901 16348
rect 2837 16288 2901 16292
rect 2917 16348 2981 16352
rect 2917 16292 2921 16348
rect 2921 16292 2977 16348
rect 2977 16292 2981 16348
rect 2917 16288 2981 16292
rect 2997 16348 3061 16352
rect 2997 16292 3001 16348
rect 3001 16292 3057 16348
rect 3057 16292 3061 16348
rect 2997 16288 3061 16292
rect 7472 16348 7536 16352
rect 7472 16292 7476 16348
rect 7476 16292 7532 16348
rect 7532 16292 7536 16348
rect 7472 16288 7536 16292
rect 7552 16348 7616 16352
rect 7552 16292 7556 16348
rect 7556 16292 7612 16348
rect 7612 16292 7616 16348
rect 7552 16288 7616 16292
rect 7632 16348 7696 16352
rect 7632 16292 7636 16348
rect 7636 16292 7692 16348
rect 7692 16292 7696 16348
rect 7632 16288 7696 16292
rect 7712 16348 7776 16352
rect 7712 16292 7716 16348
rect 7716 16292 7772 16348
rect 7772 16292 7776 16348
rect 7712 16288 7776 16292
rect 12187 16348 12251 16352
rect 12187 16292 12191 16348
rect 12191 16292 12247 16348
rect 12247 16292 12251 16348
rect 12187 16288 12251 16292
rect 12267 16348 12331 16352
rect 12267 16292 12271 16348
rect 12271 16292 12327 16348
rect 12327 16292 12331 16348
rect 12267 16288 12331 16292
rect 12347 16348 12411 16352
rect 12347 16292 12351 16348
rect 12351 16292 12407 16348
rect 12407 16292 12411 16348
rect 12347 16288 12411 16292
rect 12427 16348 12491 16352
rect 12427 16292 12431 16348
rect 12431 16292 12487 16348
rect 12487 16292 12491 16348
rect 12427 16288 12491 16292
rect 16902 16348 16966 16352
rect 16902 16292 16906 16348
rect 16906 16292 16962 16348
rect 16962 16292 16966 16348
rect 16902 16288 16966 16292
rect 16982 16348 17046 16352
rect 16982 16292 16986 16348
rect 16986 16292 17042 16348
rect 17042 16292 17046 16348
rect 16982 16288 17046 16292
rect 17062 16348 17126 16352
rect 17062 16292 17066 16348
rect 17066 16292 17122 16348
rect 17122 16292 17126 16348
rect 17062 16288 17126 16292
rect 17142 16348 17206 16352
rect 17142 16292 17146 16348
rect 17146 16292 17202 16348
rect 17202 16292 17206 16348
rect 17142 16288 17206 16292
rect 5114 15804 5178 15808
rect 5114 15748 5118 15804
rect 5118 15748 5174 15804
rect 5174 15748 5178 15804
rect 5114 15744 5178 15748
rect 5194 15804 5258 15808
rect 5194 15748 5198 15804
rect 5198 15748 5254 15804
rect 5254 15748 5258 15804
rect 5194 15744 5258 15748
rect 5274 15804 5338 15808
rect 5274 15748 5278 15804
rect 5278 15748 5334 15804
rect 5334 15748 5338 15804
rect 5274 15744 5338 15748
rect 5354 15804 5418 15808
rect 5354 15748 5358 15804
rect 5358 15748 5414 15804
rect 5414 15748 5418 15804
rect 5354 15744 5418 15748
rect 9829 15804 9893 15808
rect 9829 15748 9833 15804
rect 9833 15748 9889 15804
rect 9889 15748 9893 15804
rect 9829 15744 9893 15748
rect 9909 15804 9973 15808
rect 9909 15748 9913 15804
rect 9913 15748 9969 15804
rect 9969 15748 9973 15804
rect 9909 15744 9973 15748
rect 9989 15804 10053 15808
rect 9989 15748 9993 15804
rect 9993 15748 10049 15804
rect 10049 15748 10053 15804
rect 9989 15744 10053 15748
rect 10069 15804 10133 15808
rect 10069 15748 10073 15804
rect 10073 15748 10129 15804
rect 10129 15748 10133 15804
rect 10069 15744 10133 15748
rect 14544 15804 14608 15808
rect 14544 15748 14548 15804
rect 14548 15748 14604 15804
rect 14604 15748 14608 15804
rect 14544 15744 14608 15748
rect 14624 15804 14688 15808
rect 14624 15748 14628 15804
rect 14628 15748 14684 15804
rect 14684 15748 14688 15804
rect 14624 15744 14688 15748
rect 14704 15804 14768 15808
rect 14704 15748 14708 15804
rect 14708 15748 14764 15804
rect 14764 15748 14768 15804
rect 14704 15744 14768 15748
rect 14784 15804 14848 15808
rect 14784 15748 14788 15804
rect 14788 15748 14844 15804
rect 14844 15748 14848 15804
rect 14784 15744 14848 15748
rect 19259 15804 19323 15808
rect 19259 15748 19263 15804
rect 19263 15748 19319 15804
rect 19319 15748 19323 15804
rect 19259 15744 19323 15748
rect 19339 15804 19403 15808
rect 19339 15748 19343 15804
rect 19343 15748 19399 15804
rect 19399 15748 19403 15804
rect 19339 15744 19403 15748
rect 19419 15804 19483 15808
rect 19419 15748 19423 15804
rect 19423 15748 19479 15804
rect 19479 15748 19483 15804
rect 19419 15744 19483 15748
rect 19499 15804 19563 15808
rect 19499 15748 19503 15804
rect 19503 15748 19559 15804
rect 19559 15748 19563 15804
rect 19499 15744 19563 15748
rect 2757 15260 2821 15264
rect 2757 15204 2761 15260
rect 2761 15204 2817 15260
rect 2817 15204 2821 15260
rect 2757 15200 2821 15204
rect 2837 15260 2901 15264
rect 2837 15204 2841 15260
rect 2841 15204 2897 15260
rect 2897 15204 2901 15260
rect 2837 15200 2901 15204
rect 2917 15260 2981 15264
rect 2917 15204 2921 15260
rect 2921 15204 2977 15260
rect 2977 15204 2981 15260
rect 2917 15200 2981 15204
rect 2997 15260 3061 15264
rect 2997 15204 3001 15260
rect 3001 15204 3057 15260
rect 3057 15204 3061 15260
rect 2997 15200 3061 15204
rect 7472 15260 7536 15264
rect 7472 15204 7476 15260
rect 7476 15204 7532 15260
rect 7532 15204 7536 15260
rect 7472 15200 7536 15204
rect 7552 15260 7616 15264
rect 7552 15204 7556 15260
rect 7556 15204 7612 15260
rect 7612 15204 7616 15260
rect 7552 15200 7616 15204
rect 7632 15260 7696 15264
rect 7632 15204 7636 15260
rect 7636 15204 7692 15260
rect 7692 15204 7696 15260
rect 7632 15200 7696 15204
rect 7712 15260 7776 15264
rect 7712 15204 7716 15260
rect 7716 15204 7772 15260
rect 7772 15204 7776 15260
rect 7712 15200 7776 15204
rect 12187 15260 12251 15264
rect 12187 15204 12191 15260
rect 12191 15204 12247 15260
rect 12247 15204 12251 15260
rect 12187 15200 12251 15204
rect 12267 15260 12331 15264
rect 12267 15204 12271 15260
rect 12271 15204 12327 15260
rect 12327 15204 12331 15260
rect 12267 15200 12331 15204
rect 12347 15260 12411 15264
rect 12347 15204 12351 15260
rect 12351 15204 12407 15260
rect 12407 15204 12411 15260
rect 12347 15200 12411 15204
rect 12427 15260 12491 15264
rect 12427 15204 12431 15260
rect 12431 15204 12487 15260
rect 12487 15204 12491 15260
rect 12427 15200 12491 15204
rect 16902 15260 16966 15264
rect 16902 15204 16906 15260
rect 16906 15204 16962 15260
rect 16962 15204 16966 15260
rect 16902 15200 16966 15204
rect 16982 15260 17046 15264
rect 16982 15204 16986 15260
rect 16986 15204 17042 15260
rect 17042 15204 17046 15260
rect 16982 15200 17046 15204
rect 17062 15260 17126 15264
rect 17062 15204 17066 15260
rect 17066 15204 17122 15260
rect 17122 15204 17126 15260
rect 17062 15200 17126 15204
rect 17142 15260 17206 15264
rect 17142 15204 17146 15260
rect 17146 15204 17202 15260
rect 17202 15204 17206 15260
rect 17142 15200 17206 15204
rect 5114 14716 5178 14720
rect 5114 14660 5118 14716
rect 5118 14660 5174 14716
rect 5174 14660 5178 14716
rect 5114 14656 5178 14660
rect 5194 14716 5258 14720
rect 5194 14660 5198 14716
rect 5198 14660 5254 14716
rect 5254 14660 5258 14716
rect 5194 14656 5258 14660
rect 5274 14716 5338 14720
rect 5274 14660 5278 14716
rect 5278 14660 5334 14716
rect 5334 14660 5338 14716
rect 5274 14656 5338 14660
rect 5354 14716 5418 14720
rect 5354 14660 5358 14716
rect 5358 14660 5414 14716
rect 5414 14660 5418 14716
rect 5354 14656 5418 14660
rect 9829 14716 9893 14720
rect 9829 14660 9833 14716
rect 9833 14660 9889 14716
rect 9889 14660 9893 14716
rect 9829 14656 9893 14660
rect 9909 14716 9973 14720
rect 9909 14660 9913 14716
rect 9913 14660 9969 14716
rect 9969 14660 9973 14716
rect 9909 14656 9973 14660
rect 9989 14716 10053 14720
rect 9989 14660 9993 14716
rect 9993 14660 10049 14716
rect 10049 14660 10053 14716
rect 9989 14656 10053 14660
rect 10069 14716 10133 14720
rect 10069 14660 10073 14716
rect 10073 14660 10129 14716
rect 10129 14660 10133 14716
rect 10069 14656 10133 14660
rect 14544 14716 14608 14720
rect 14544 14660 14548 14716
rect 14548 14660 14604 14716
rect 14604 14660 14608 14716
rect 14544 14656 14608 14660
rect 14624 14716 14688 14720
rect 14624 14660 14628 14716
rect 14628 14660 14684 14716
rect 14684 14660 14688 14716
rect 14624 14656 14688 14660
rect 14704 14716 14768 14720
rect 14704 14660 14708 14716
rect 14708 14660 14764 14716
rect 14764 14660 14768 14716
rect 14704 14656 14768 14660
rect 14784 14716 14848 14720
rect 14784 14660 14788 14716
rect 14788 14660 14844 14716
rect 14844 14660 14848 14716
rect 14784 14656 14848 14660
rect 19259 14716 19323 14720
rect 19259 14660 19263 14716
rect 19263 14660 19319 14716
rect 19319 14660 19323 14716
rect 19259 14656 19323 14660
rect 19339 14716 19403 14720
rect 19339 14660 19343 14716
rect 19343 14660 19399 14716
rect 19399 14660 19403 14716
rect 19339 14656 19403 14660
rect 19419 14716 19483 14720
rect 19419 14660 19423 14716
rect 19423 14660 19479 14716
rect 19479 14660 19483 14716
rect 19419 14656 19483 14660
rect 19499 14716 19563 14720
rect 19499 14660 19503 14716
rect 19503 14660 19559 14716
rect 19559 14660 19563 14716
rect 19499 14656 19563 14660
rect 2757 14172 2821 14176
rect 2757 14116 2761 14172
rect 2761 14116 2817 14172
rect 2817 14116 2821 14172
rect 2757 14112 2821 14116
rect 2837 14172 2901 14176
rect 2837 14116 2841 14172
rect 2841 14116 2897 14172
rect 2897 14116 2901 14172
rect 2837 14112 2901 14116
rect 2917 14172 2981 14176
rect 2917 14116 2921 14172
rect 2921 14116 2977 14172
rect 2977 14116 2981 14172
rect 2917 14112 2981 14116
rect 2997 14172 3061 14176
rect 2997 14116 3001 14172
rect 3001 14116 3057 14172
rect 3057 14116 3061 14172
rect 2997 14112 3061 14116
rect 7472 14172 7536 14176
rect 7472 14116 7476 14172
rect 7476 14116 7532 14172
rect 7532 14116 7536 14172
rect 7472 14112 7536 14116
rect 7552 14172 7616 14176
rect 7552 14116 7556 14172
rect 7556 14116 7612 14172
rect 7612 14116 7616 14172
rect 7552 14112 7616 14116
rect 7632 14172 7696 14176
rect 7632 14116 7636 14172
rect 7636 14116 7692 14172
rect 7692 14116 7696 14172
rect 7632 14112 7696 14116
rect 7712 14172 7776 14176
rect 7712 14116 7716 14172
rect 7716 14116 7772 14172
rect 7772 14116 7776 14172
rect 7712 14112 7776 14116
rect 12187 14172 12251 14176
rect 12187 14116 12191 14172
rect 12191 14116 12247 14172
rect 12247 14116 12251 14172
rect 12187 14112 12251 14116
rect 12267 14172 12331 14176
rect 12267 14116 12271 14172
rect 12271 14116 12327 14172
rect 12327 14116 12331 14172
rect 12267 14112 12331 14116
rect 12347 14172 12411 14176
rect 12347 14116 12351 14172
rect 12351 14116 12407 14172
rect 12407 14116 12411 14172
rect 12347 14112 12411 14116
rect 12427 14172 12491 14176
rect 12427 14116 12431 14172
rect 12431 14116 12487 14172
rect 12487 14116 12491 14172
rect 12427 14112 12491 14116
rect 16902 14172 16966 14176
rect 16902 14116 16906 14172
rect 16906 14116 16962 14172
rect 16962 14116 16966 14172
rect 16902 14112 16966 14116
rect 16982 14172 17046 14176
rect 16982 14116 16986 14172
rect 16986 14116 17042 14172
rect 17042 14116 17046 14172
rect 16982 14112 17046 14116
rect 17062 14172 17126 14176
rect 17062 14116 17066 14172
rect 17066 14116 17122 14172
rect 17122 14116 17126 14172
rect 17062 14112 17126 14116
rect 17142 14172 17206 14176
rect 17142 14116 17146 14172
rect 17146 14116 17202 14172
rect 17202 14116 17206 14172
rect 17142 14112 17206 14116
rect 5114 13628 5178 13632
rect 5114 13572 5118 13628
rect 5118 13572 5174 13628
rect 5174 13572 5178 13628
rect 5114 13568 5178 13572
rect 5194 13628 5258 13632
rect 5194 13572 5198 13628
rect 5198 13572 5254 13628
rect 5254 13572 5258 13628
rect 5194 13568 5258 13572
rect 5274 13628 5338 13632
rect 5274 13572 5278 13628
rect 5278 13572 5334 13628
rect 5334 13572 5338 13628
rect 5274 13568 5338 13572
rect 5354 13628 5418 13632
rect 5354 13572 5358 13628
rect 5358 13572 5414 13628
rect 5414 13572 5418 13628
rect 5354 13568 5418 13572
rect 9829 13628 9893 13632
rect 9829 13572 9833 13628
rect 9833 13572 9889 13628
rect 9889 13572 9893 13628
rect 9829 13568 9893 13572
rect 9909 13628 9973 13632
rect 9909 13572 9913 13628
rect 9913 13572 9969 13628
rect 9969 13572 9973 13628
rect 9909 13568 9973 13572
rect 9989 13628 10053 13632
rect 9989 13572 9993 13628
rect 9993 13572 10049 13628
rect 10049 13572 10053 13628
rect 9989 13568 10053 13572
rect 10069 13628 10133 13632
rect 10069 13572 10073 13628
rect 10073 13572 10129 13628
rect 10129 13572 10133 13628
rect 10069 13568 10133 13572
rect 14544 13628 14608 13632
rect 14544 13572 14548 13628
rect 14548 13572 14604 13628
rect 14604 13572 14608 13628
rect 14544 13568 14608 13572
rect 14624 13628 14688 13632
rect 14624 13572 14628 13628
rect 14628 13572 14684 13628
rect 14684 13572 14688 13628
rect 14624 13568 14688 13572
rect 14704 13628 14768 13632
rect 14704 13572 14708 13628
rect 14708 13572 14764 13628
rect 14764 13572 14768 13628
rect 14704 13568 14768 13572
rect 14784 13628 14848 13632
rect 14784 13572 14788 13628
rect 14788 13572 14844 13628
rect 14844 13572 14848 13628
rect 14784 13568 14848 13572
rect 19259 13628 19323 13632
rect 19259 13572 19263 13628
rect 19263 13572 19319 13628
rect 19319 13572 19323 13628
rect 19259 13568 19323 13572
rect 19339 13628 19403 13632
rect 19339 13572 19343 13628
rect 19343 13572 19399 13628
rect 19399 13572 19403 13628
rect 19339 13568 19403 13572
rect 19419 13628 19483 13632
rect 19419 13572 19423 13628
rect 19423 13572 19479 13628
rect 19479 13572 19483 13628
rect 19419 13568 19483 13572
rect 19499 13628 19563 13632
rect 19499 13572 19503 13628
rect 19503 13572 19559 13628
rect 19559 13572 19563 13628
rect 19499 13568 19563 13572
rect 2757 13084 2821 13088
rect 2757 13028 2761 13084
rect 2761 13028 2817 13084
rect 2817 13028 2821 13084
rect 2757 13024 2821 13028
rect 2837 13084 2901 13088
rect 2837 13028 2841 13084
rect 2841 13028 2897 13084
rect 2897 13028 2901 13084
rect 2837 13024 2901 13028
rect 2917 13084 2981 13088
rect 2917 13028 2921 13084
rect 2921 13028 2977 13084
rect 2977 13028 2981 13084
rect 2917 13024 2981 13028
rect 2997 13084 3061 13088
rect 2997 13028 3001 13084
rect 3001 13028 3057 13084
rect 3057 13028 3061 13084
rect 2997 13024 3061 13028
rect 7472 13084 7536 13088
rect 7472 13028 7476 13084
rect 7476 13028 7532 13084
rect 7532 13028 7536 13084
rect 7472 13024 7536 13028
rect 7552 13084 7616 13088
rect 7552 13028 7556 13084
rect 7556 13028 7612 13084
rect 7612 13028 7616 13084
rect 7552 13024 7616 13028
rect 7632 13084 7696 13088
rect 7632 13028 7636 13084
rect 7636 13028 7692 13084
rect 7692 13028 7696 13084
rect 7632 13024 7696 13028
rect 7712 13084 7776 13088
rect 7712 13028 7716 13084
rect 7716 13028 7772 13084
rect 7772 13028 7776 13084
rect 7712 13024 7776 13028
rect 12187 13084 12251 13088
rect 12187 13028 12191 13084
rect 12191 13028 12247 13084
rect 12247 13028 12251 13084
rect 12187 13024 12251 13028
rect 12267 13084 12331 13088
rect 12267 13028 12271 13084
rect 12271 13028 12327 13084
rect 12327 13028 12331 13084
rect 12267 13024 12331 13028
rect 12347 13084 12411 13088
rect 12347 13028 12351 13084
rect 12351 13028 12407 13084
rect 12407 13028 12411 13084
rect 12347 13024 12411 13028
rect 12427 13084 12491 13088
rect 12427 13028 12431 13084
rect 12431 13028 12487 13084
rect 12487 13028 12491 13084
rect 12427 13024 12491 13028
rect 16902 13084 16966 13088
rect 16902 13028 16906 13084
rect 16906 13028 16962 13084
rect 16962 13028 16966 13084
rect 16902 13024 16966 13028
rect 16982 13084 17046 13088
rect 16982 13028 16986 13084
rect 16986 13028 17042 13084
rect 17042 13028 17046 13084
rect 16982 13024 17046 13028
rect 17062 13084 17126 13088
rect 17062 13028 17066 13084
rect 17066 13028 17122 13084
rect 17122 13028 17126 13084
rect 17062 13024 17126 13028
rect 17142 13084 17206 13088
rect 17142 13028 17146 13084
rect 17146 13028 17202 13084
rect 17202 13028 17206 13084
rect 17142 13024 17206 13028
rect 10732 12608 10796 12612
rect 10732 12552 10746 12608
rect 10746 12552 10796 12608
rect 10732 12548 10796 12552
rect 5114 12540 5178 12544
rect 5114 12484 5118 12540
rect 5118 12484 5174 12540
rect 5174 12484 5178 12540
rect 5114 12480 5178 12484
rect 5194 12540 5258 12544
rect 5194 12484 5198 12540
rect 5198 12484 5254 12540
rect 5254 12484 5258 12540
rect 5194 12480 5258 12484
rect 5274 12540 5338 12544
rect 5274 12484 5278 12540
rect 5278 12484 5334 12540
rect 5334 12484 5338 12540
rect 5274 12480 5338 12484
rect 5354 12540 5418 12544
rect 5354 12484 5358 12540
rect 5358 12484 5414 12540
rect 5414 12484 5418 12540
rect 5354 12480 5418 12484
rect 9829 12540 9893 12544
rect 9829 12484 9833 12540
rect 9833 12484 9889 12540
rect 9889 12484 9893 12540
rect 9829 12480 9893 12484
rect 9909 12540 9973 12544
rect 9909 12484 9913 12540
rect 9913 12484 9969 12540
rect 9969 12484 9973 12540
rect 9909 12480 9973 12484
rect 9989 12540 10053 12544
rect 9989 12484 9993 12540
rect 9993 12484 10049 12540
rect 10049 12484 10053 12540
rect 9989 12480 10053 12484
rect 10069 12540 10133 12544
rect 10069 12484 10073 12540
rect 10073 12484 10129 12540
rect 10129 12484 10133 12540
rect 10069 12480 10133 12484
rect 14544 12540 14608 12544
rect 14544 12484 14548 12540
rect 14548 12484 14604 12540
rect 14604 12484 14608 12540
rect 14544 12480 14608 12484
rect 14624 12540 14688 12544
rect 14624 12484 14628 12540
rect 14628 12484 14684 12540
rect 14684 12484 14688 12540
rect 14624 12480 14688 12484
rect 14704 12540 14768 12544
rect 14704 12484 14708 12540
rect 14708 12484 14764 12540
rect 14764 12484 14768 12540
rect 14704 12480 14768 12484
rect 14784 12540 14848 12544
rect 14784 12484 14788 12540
rect 14788 12484 14844 12540
rect 14844 12484 14848 12540
rect 14784 12480 14848 12484
rect 19259 12540 19323 12544
rect 19259 12484 19263 12540
rect 19263 12484 19319 12540
rect 19319 12484 19323 12540
rect 19259 12480 19323 12484
rect 19339 12540 19403 12544
rect 19339 12484 19343 12540
rect 19343 12484 19399 12540
rect 19399 12484 19403 12540
rect 19339 12480 19403 12484
rect 19419 12540 19483 12544
rect 19419 12484 19423 12540
rect 19423 12484 19479 12540
rect 19479 12484 19483 12540
rect 19419 12480 19483 12484
rect 19499 12540 19563 12544
rect 19499 12484 19503 12540
rect 19503 12484 19559 12540
rect 19559 12484 19563 12540
rect 19499 12480 19563 12484
rect 2757 11996 2821 12000
rect 2757 11940 2761 11996
rect 2761 11940 2817 11996
rect 2817 11940 2821 11996
rect 2757 11936 2821 11940
rect 2837 11996 2901 12000
rect 2837 11940 2841 11996
rect 2841 11940 2897 11996
rect 2897 11940 2901 11996
rect 2837 11936 2901 11940
rect 2917 11996 2981 12000
rect 2917 11940 2921 11996
rect 2921 11940 2977 11996
rect 2977 11940 2981 11996
rect 2917 11936 2981 11940
rect 2997 11996 3061 12000
rect 2997 11940 3001 11996
rect 3001 11940 3057 11996
rect 3057 11940 3061 11996
rect 2997 11936 3061 11940
rect 7472 11996 7536 12000
rect 7472 11940 7476 11996
rect 7476 11940 7532 11996
rect 7532 11940 7536 11996
rect 7472 11936 7536 11940
rect 7552 11996 7616 12000
rect 7552 11940 7556 11996
rect 7556 11940 7612 11996
rect 7612 11940 7616 11996
rect 7552 11936 7616 11940
rect 7632 11996 7696 12000
rect 7632 11940 7636 11996
rect 7636 11940 7692 11996
rect 7692 11940 7696 11996
rect 7632 11936 7696 11940
rect 7712 11996 7776 12000
rect 7712 11940 7716 11996
rect 7716 11940 7772 11996
rect 7772 11940 7776 11996
rect 7712 11936 7776 11940
rect 12187 11996 12251 12000
rect 12187 11940 12191 11996
rect 12191 11940 12247 11996
rect 12247 11940 12251 11996
rect 12187 11936 12251 11940
rect 12267 11996 12331 12000
rect 12267 11940 12271 11996
rect 12271 11940 12327 11996
rect 12327 11940 12331 11996
rect 12267 11936 12331 11940
rect 12347 11996 12411 12000
rect 12347 11940 12351 11996
rect 12351 11940 12407 11996
rect 12407 11940 12411 11996
rect 12347 11936 12411 11940
rect 12427 11996 12491 12000
rect 12427 11940 12431 11996
rect 12431 11940 12487 11996
rect 12487 11940 12491 11996
rect 12427 11936 12491 11940
rect 16902 11996 16966 12000
rect 16902 11940 16906 11996
rect 16906 11940 16962 11996
rect 16962 11940 16966 11996
rect 16902 11936 16966 11940
rect 16982 11996 17046 12000
rect 16982 11940 16986 11996
rect 16986 11940 17042 11996
rect 17042 11940 17046 11996
rect 16982 11936 17046 11940
rect 17062 11996 17126 12000
rect 17062 11940 17066 11996
rect 17066 11940 17122 11996
rect 17122 11940 17126 11996
rect 17062 11936 17126 11940
rect 17142 11996 17206 12000
rect 17142 11940 17146 11996
rect 17146 11940 17202 11996
rect 17202 11940 17206 11996
rect 17142 11936 17206 11940
rect 9628 11596 9692 11660
rect 5114 11452 5178 11456
rect 5114 11396 5118 11452
rect 5118 11396 5174 11452
rect 5174 11396 5178 11452
rect 5114 11392 5178 11396
rect 5194 11452 5258 11456
rect 5194 11396 5198 11452
rect 5198 11396 5254 11452
rect 5254 11396 5258 11452
rect 5194 11392 5258 11396
rect 5274 11452 5338 11456
rect 5274 11396 5278 11452
rect 5278 11396 5334 11452
rect 5334 11396 5338 11452
rect 5274 11392 5338 11396
rect 5354 11452 5418 11456
rect 5354 11396 5358 11452
rect 5358 11396 5414 11452
rect 5414 11396 5418 11452
rect 5354 11392 5418 11396
rect 9829 11452 9893 11456
rect 9829 11396 9833 11452
rect 9833 11396 9889 11452
rect 9889 11396 9893 11452
rect 9829 11392 9893 11396
rect 9909 11452 9973 11456
rect 9909 11396 9913 11452
rect 9913 11396 9969 11452
rect 9969 11396 9973 11452
rect 9909 11392 9973 11396
rect 9989 11452 10053 11456
rect 9989 11396 9993 11452
rect 9993 11396 10049 11452
rect 10049 11396 10053 11452
rect 9989 11392 10053 11396
rect 10069 11452 10133 11456
rect 10069 11396 10073 11452
rect 10073 11396 10129 11452
rect 10129 11396 10133 11452
rect 10069 11392 10133 11396
rect 14544 11452 14608 11456
rect 14544 11396 14548 11452
rect 14548 11396 14604 11452
rect 14604 11396 14608 11452
rect 14544 11392 14608 11396
rect 14624 11452 14688 11456
rect 14624 11396 14628 11452
rect 14628 11396 14684 11452
rect 14684 11396 14688 11452
rect 14624 11392 14688 11396
rect 14704 11452 14768 11456
rect 14704 11396 14708 11452
rect 14708 11396 14764 11452
rect 14764 11396 14768 11452
rect 14704 11392 14768 11396
rect 14784 11452 14848 11456
rect 14784 11396 14788 11452
rect 14788 11396 14844 11452
rect 14844 11396 14848 11452
rect 14784 11392 14848 11396
rect 19259 11452 19323 11456
rect 19259 11396 19263 11452
rect 19263 11396 19319 11452
rect 19319 11396 19323 11452
rect 19259 11392 19323 11396
rect 19339 11452 19403 11456
rect 19339 11396 19343 11452
rect 19343 11396 19399 11452
rect 19399 11396 19403 11452
rect 19339 11392 19403 11396
rect 19419 11452 19483 11456
rect 19419 11396 19423 11452
rect 19423 11396 19479 11452
rect 19479 11396 19483 11452
rect 19419 11392 19483 11396
rect 19499 11452 19563 11456
rect 19499 11396 19503 11452
rect 19503 11396 19559 11452
rect 19559 11396 19563 11452
rect 19499 11392 19563 11396
rect 2757 10908 2821 10912
rect 2757 10852 2761 10908
rect 2761 10852 2817 10908
rect 2817 10852 2821 10908
rect 2757 10848 2821 10852
rect 2837 10908 2901 10912
rect 2837 10852 2841 10908
rect 2841 10852 2897 10908
rect 2897 10852 2901 10908
rect 2837 10848 2901 10852
rect 2917 10908 2981 10912
rect 2917 10852 2921 10908
rect 2921 10852 2977 10908
rect 2977 10852 2981 10908
rect 2917 10848 2981 10852
rect 2997 10908 3061 10912
rect 2997 10852 3001 10908
rect 3001 10852 3057 10908
rect 3057 10852 3061 10908
rect 2997 10848 3061 10852
rect 7472 10908 7536 10912
rect 7472 10852 7476 10908
rect 7476 10852 7532 10908
rect 7532 10852 7536 10908
rect 7472 10848 7536 10852
rect 7552 10908 7616 10912
rect 7552 10852 7556 10908
rect 7556 10852 7612 10908
rect 7612 10852 7616 10908
rect 7552 10848 7616 10852
rect 7632 10908 7696 10912
rect 7632 10852 7636 10908
rect 7636 10852 7692 10908
rect 7692 10852 7696 10908
rect 7632 10848 7696 10852
rect 7712 10908 7776 10912
rect 7712 10852 7716 10908
rect 7716 10852 7772 10908
rect 7772 10852 7776 10908
rect 7712 10848 7776 10852
rect 12187 10908 12251 10912
rect 12187 10852 12191 10908
rect 12191 10852 12247 10908
rect 12247 10852 12251 10908
rect 12187 10848 12251 10852
rect 12267 10908 12331 10912
rect 12267 10852 12271 10908
rect 12271 10852 12327 10908
rect 12327 10852 12331 10908
rect 12267 10848 12331 10852
rect 12347 10908 12411 10912
rect 12347 10852 12351 10908
rect 12351 10852 12407 10908
rect 12407 10852 12411 10908
rect 12347 10848 12411 10852
rect 12427 10908 12491 10912
rect 12427 10852 12431 10908
rect 12431 10852 12487 10908
rect 12487 10852 12491 10908
rect 12427 10848 12491 10852
rect 16902 10908 16966 10912
rect 16902 10852 16906 10908
rect 16906 10852 16962 10908
rect 16962 10852 16966 10908
rect 16902 10848 16966 10852
rect 16982 10908 17046 10912
rect 16982 10852 16986 10908
rect 16986 10852 17042 10908
rect 17042 10852 17046 10908
rect 16982 10848 17046 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 5114 10364 5178 10368
rect 5114 10308 5118 10364
rect 5118 10308 5174 10364
rect 5174 10308 5178 10364
rect 5114 10304 5178 10308
rect 5194 10364 5258 10368
rect 5194 10308 5198 10364
rect 5198 10308 5254 10364
rect 5254 10308 5258 10364
rect 5194 10304 5258 10308
rect 5274 10364 5338 10368
rect 5274 10308 5278 10364
rect 5278 10308 5334 10364
rect 5334 10308 5338 10364
rect 5274 10304 5338 10308
rect 5354 10364 5418 10368
rect 5354 10308 5358 10364
rect 5358 10308 5414 10364
rect 5414 10308 5418 10364
rect 5354 10304 5418 10308
rect 9829 10364 9893 10368
rect 9829 10308 9833 10364
rect 9833 10308 9889 10364
rect 9889 10308 9893 10364
rect 9829 10304 9893 10308
rect 9909 10364 9973 10368
rect 9909 10308 9913 10364
rect 9913 10308 9969 10364
rect 9969 10308 9973 10364
rect 9909 10304 9973 10308
rect 9989 10364 10053 10368
rect 9989 10308 9993 10364
rect 9993 10308 10049 10364
rect 10049 10308 10053 10364
rect 9989 10304 10053 10308
rect 10069 10364 10133 10368
rect 10069 10308 10073 10364
rect 10073 10308 10129 10364
rect 10129 10308 10133 10364
rect 10069 10304 10133 10308
rect 14544 10364 14608 10368
rect 14544 10308 14548 10364
rect 14548 10308 14604 10364
rect 14604 10308 14608 10364
rect 14544 10304 14608 10308
rect 14624 10364 14688 10368
rect 14624 10308 14628 10364
rect 14628 10308 14684 10364
rect 14684 10308 14688 10364
rect 14624 10304 14688 10308
rect 14704 10364 14768 10368
rect 14704 10308 14708 10364
rect 14708 10308 14764 10364
rect 14764 10308 14768 10364
rect 14704 10304 14768 10308
rect 14784 10364 14848 10368
rect 14784 10308 14788 10364
rect 14788 10308 14844 10364
rect 14844 10308 14848 10364
rect 14784 10304 14848 10308
rect 19259 10364 19323 10368
rect 19259 10308 19263 10364
rect 19263 10308 19319 10364
rect 19319 10308 19323 10364
rect 19259 10304 19323 10308
rect 19339 10364 19403 10368
rect 19339 10308 19343 10364
rect 19343 10308 19399 10364
rect 19399 10308 19403 10364
rect 19339 10304 19403 10308
rect 19419 10364 19483 10368
rect 19419 10308 19423 10364
rect 19423 10308 19479 10364
rect 19479 10308 19483 10364
rect 19419 10304 19483 10308
rect 19499 10364 19563 10368
rect 19499 10308 19503 10364
rect 19503 10308 19559 10364
rect 19559 10308 19563 10364
rect 19499 10304 19563 10308
rect 2757 9820 2821 9824
rect 2757 9764 2761 9820
rect 2761 9764 2817 9820
rect 2817 9764 2821 9820
rect 2757 9760 2821 9764
rect 2837 9820 2901 9824
rect 2837 9764 2841 9820
rect 2841 9764 2897 9820
rect 2897 9764 2901 9820
rect 2837 9760 2901 9764
rect 2917 9820 2981 9824
rect 2917 9764 2921 9820
rect 2921 9764 2977 9820
rect 2977 9764 2981 9820
rect 2917 9760 2981 9764
rect 2997 9820 3061 9824
rect 2997 9764 3001 9820
rect 3001 9764 3057 9820
rect 3057 9764 3061 9820
rect 2997 9760 3061 9764
rect 7472 9820 7536 9824
rect 7472 9764 7476 9820
rect 7476 9764 7532 9820
rect 7532 9764 7536 9820
rect 7472 9760 7536 9764
rect 7552 9820 7616 9824
rect 7552 9764 7556 9820
rect 7556 9764 7612 9820
rect 7612 9764 7616 9820
rect 7552 9760 7616 9764
rect 7632 9820 7696 9824
rect 7632 9764 7636 9820
rect 7636 9764 7692 9820
rect 7692 9764 7696 9820
rect 7632 9760 7696 9764
rect 7712 9820 7776 9824
rect 7712 9764 7716 9820
rect 7716 9764 7772 9820
rect 7772 9764 7776 9820
rect 7712 9760 7776 9764
rect 12187 9820 12251 9824
rect 12187 9764 12191 9820
rect 12191 9764 12247 9820
rect 12247 9764 12251 9820
rect 12187 9760 12251 9764
rect 12267 9820 12331 9824
rect 12267 9764 12271 9820
rect 12271 9764 12327 9820
rect 12327 9764 12331 9820
rect 12267 9760 12331 9764
rect 12347 9820 12411 9824
rect 12347 9764 12351 9820
rect 12351 9764 12407 9820
rect 12407 9764 12411 9820
rect 12347 9760 12411 9764
rect 12427 9820 12491 9824
rect 12427 9764 12431 9820
rect 12431 9764 12487 9820
rect 12487 9764 12491 9820
rect 12427 9760 12491 9764
rect 16902 9820 16966 9824
rect 16902 9764 16906 9820
rect 16906 9764 16962 9820
rect 16962 9764 16966 9820
rect 16902 9760 16966 9764
rect 16982 9820 17046 9824
rect 16982 9764 16986 9820
rect 16986 9764 17042 9820
rect 17042 9764 17046 9820
rect 16982 9760 17046 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 11468 9692 11532 9756
rect 5114 9276 5178 9280
rect 5114 9220 5118 9276
rect 5118 9220 5174 9276
rect 5174 9220 5178 9276
rect 5114 9216 5178 9220
rect 5194 9276 5258 9280
rect 5194 9220 5198 9276
rect 5198 9220 5254 9276
rect 5254 9220 5258 9276
rect 5194 9216 5258 9220
rect 5274 9276 5338 9280
rect 5274 9220 5278 9276
rect 5278 9220 5334 9276
rect 5334 9220 5338 9276
rect 5274 9216 5338 9220
rect 5354 9276 5418 9280
rect 5354 9220 5358 9276
rect 5358 9220 5414 9276
rect 5414 9220 5418 9276
rect 5354 9216 5418 9220
rect 9829 9276 9893 9280
rect 9829 9220 9833 9276
rect 9833 9220 9889 9276
rect 9889 9220 9893 9276
rect 9829 9216 9893 9220
rect 9909 9276 9973 9280
rect 9909 9220 9913 9276
rect 9913 9220 9969 9276
rect 9969 9220 9973 9276
rect 9909 9216 9973 9220
rect 9989 9276 10053 9280
rect 9989 9220 9993 9276
rect 9993 9220 10049 9276
rect 10049 9220 10053 9276
rect 9989 9216 10053 9220
rect 10069 9276 10133 9280
rect 10069 9220 10073 9276
rect 10073 9220 10129 9276
rect 10129 9220 10133 9276
rect 10069 9216 10133 9220
rect 14544 9276 14608 9280
rect 14544 9220 14548 9276
rect 14548 9220 14604 9276
rect 14604 9220 14608 9276
rect 14544 9216 14608 9220
rect 14624 9276 14688 9280
rect 14624 9220 14628 9276
rect 14628 9220 14684 9276
rect 14684 9220 14688 9276
rect 14624 9216 14688 9220
rect 14704 9276 14768 9280
rect 14704 9220 14708 9276
rect 14708 9220 14764 9276
rect 14764 9220 14768 9276
rect 14704 9216 14768 9220
rect 14784 9276 14848 9280
rect 14784 9220 14788 9276
rect 14788 9220 14844 9276
rect 14844 9220 14848 9276
rect 14784 9216 14848 9220
rect 19259 9276 19323 9280
rect 19259 9220 19263 9276
rect 19263 9220 19319 9276
rect 19319 9220 19323 9276
rect 19259 9216 19323 9220
rect 19339 9276 19403 9280
rect 19339 9220 19343 9276
rect 19343 9220 19399 9276
rect 19399 9220 19403 9276
rect 19339 9216 19403 9220
rect 19419 9276 19483 9280
rect 19419 9220 19423 9276
rect 19423 9220 19479 9276
rect 19479 9220 19483 9276
rect 19419 9216 19483 9220
rect 19499 9276 19563 9280
rect 19499 9220 19503 9276
rect 19503 9220 19559 9276
rect 19559 9220 19563 9276
rect 19499 9216 19563 9220
rect 2757 8732 2821 8736
rect 2757 8676 2761 8732
rect 2761 8676 2817 8732
rect 2817 8676 2821 8732
rect 2757 8672 2821 8676
rect 2837 8732 2901 8736
rect 2837 8676 2841 8732
rect 2841 8676 2897 8732
rect 2897 8676 2901 8732
rect 2837 8672 2901 8676
rect 2917 8732 2981 8736
rect 2917 8676 2921 8732
rect 2921 8676 2977 8732
rect 2977 8676 2981 8732
rect 2917 8672 2981 8676
rect 2997 8732 3061 8736
rect 2997 8676 3001 8732
rect 3001 8676 3057 8732
rect 3057 8676 3061 8732
rect 2997 8672 3061 8676
rect 7472 8732 7536 8736
rect 7472 8676 7476 8732
rect 7476 8676 7532 8732
rect 7532 8676 7536 8732
rect 7472 8672 7536 8676
rect 7552 8732 7616 8736
rect 7552 8676 7556 8732
rect 7556 8676 7612 8732
rect 7612 8676 7616 8732
rect 7552 8672 7616 8676
rect 7632 8732 7696 8736
rect 7632 8676 7636 8732
rect 7636 8676 7692 8732
rect 7692 8676 7696 8732
rect 7632 8672 7696 8676
rect 7712 8732 7776 8736
rect 7712 8676 7716 8732
rect 7716 8676 7772 8732
rect 7772 8676 7776 8732
rect 7712 8672 7776 8676
rect 12187 8732 12251 8736
rect 12187 8676 12191 8732
rect 12191 8676 12247 8732
rect 12247 8676 12251 8732
rect 12187 8672 12251 8676
rect 12267 8732 12331 8736
rect 12267 8676 12271 8732
rect 12271 8676 12327 8732
rect 12327 8676 12331 8732
rect 12267 8672 12331 8676
rect 12347 8732 12411 8736
rect 12347 8676 12351 8732
rect 12351 8676 12407 8732
rect 12407 8676 12411 8732
rect 12347 8672 12411 8676
rect 12427 8732 12491 8736
rect 12427 8676 12431 8732
rect 12431 8676 12487 8732
rect 12487 8676 12491 8732
rect 12427 8672 12491 8676
rect 16902 8732 16966 8736
rect 16902 8676 16906 8732
rect 16906 8676 16962 8732
rect 16962 8676 16966 8732
rect 16902 8672 16966 8676
rect 16982 8732 17046 8736
rect 16982 8676 16986 8732
rect 16986 8676 17042 8732
rect 17042 8676 17046 8732
rect 16982 8672 17046 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 11100 8256 11164 8260
rect 11100 8200 11150 8256
rect 11150 8200 11164 8256
rect 11100 8196 11164 8200
rect 5114 8188 5178 8192
rect 5114 8132 5118 8188
rect 5118 8132 5174 8188
rect 5174 8132 5178 8188
rect 5114 8128 5178 8132
rect 5194 8188 5258 8192
rect 5194 8132 5198 8188
rect 5198 8132 5254 8188
rect 5254 8132 5258 8188
rect 5194 8128 5258 8132
rect 5274 8188 5338 8192
rect 5274 8132 5278 8188
rect 5278 8132 5334 8188
rect 5334 8132 5338 8188
rect 5274 8128 5338 8132
rect 5354 8188 5418 8192
rect 5354 8132 5358 8188
rect 5358 8132 5414 8188
rect 5414 8132 5418 8188
rect 5354 8128 5418 8132
rect 9829 8188 9893 8192
rect 9829 8132 9833 8188
rect 9833 8132 9889 8188
rect 9889 8132 9893 8188
rect 9829 8128 9893 8132
rect 9909 8188 9973 8192
rect 9909 8132 9913 8188
rect 9913 8132 9969 8188
rect 9969 8132 9973 8188
rect 9909 8128 9973 8132
rect 9989 8188 10053 8192
rect 9989 8132 9993 8188
rect 9993 8132 10049 8188
rect 10049 8132 10053 8188
rect 9989 8128 10053 8132
rect 10069 8188 10133 8192
rect 10069 8132 10073 8188
rect 10073 8132 10129 8188
rect 10129 8132 10133 8188
rect 10069 8128 10133 8132
rect 14544 8188 14608 8192
rect 14544 8132 14548 8188
rect 14548 8132 14604 8188
rect 14604 8132 14608 8188
rect 14544 8128 14608 8132
rect 14624 8188 14688 8192
rect 14624 8132 14628 8188
rect 14628 8132 14684 8188
rect 14684 8132 14688 8188
rect 14624 8128 14688 8132
rect 14704 8188 14768 8192
rect 14704 8132 14708 8188
rect 14708 8132 14764 8188
rect 14764 8132 14768 8188
rect 14704 8128 14768 8132
rect 14784 8188 14848 8192
rect 14784 8132 14788 8188
rect 14788 8132 14844 8188
rect 14844 8132 14848 8188
rect 14784 8128 14848 8132
rect 19259 8188 19323 8192
rect 19259 8132 19263 8188
rect 19263 8132 19319 8188
rect 19319 8132 19323 8188
rect 19259 8128 19323 8132
rect 19339 8188 19403 8192
rect 19339 8132 19343 8188
rect 19343 8132 19399 8188
rect 19399 8132 19403 8188
rect 19339 8128 19403 8132
rect 19419 8188 19483 8192
rect 19419 8132 19423 8188
rect 19423 8132 19479 8188
rect 19479 8132 19483 8188
rect 19419 8128 19483 8132
rect 19499 8188 19563 8192
rect 19499 8132 19503 8188
rect 19503 8132 19559 8188
rect 19559 8132 19563 8188
rect 19499 8128 19563 8132
rect 2757 7644 2821 7648
rect 2757 7588 2761 7644
rect 2761 7588 2817 7644
rect 2817 7588 2821 7644
rect 2757 7584 2821 7588
rect 2837 7644 2901 7648
rect 2837 7588 2841 7644
rect 2841 7588 2897 7644
rect 2897 7588 2901 7644
rect 2837 7584 2901 7588
rect 2917 7644 2981 7648
rect 2917 7588 2921 7644
rect 2921 7588 2977 7644
rect 2977 7588 2981 7644
rect 2917 7584 2981 7588
rect 2997 7644 3061 7648
rect 2997 7588 3001 7644
rect 3001 7588 3057 7644
rect 3057 7588 3061 7644
rect 2997 7584 3061 7588
rect 7472 7644 7536 7648
rect 7472 7588 7476 7644
rect 7476 7588 7532 7644
rect 7532 7588 7536 7644
rect 7472 7584 7536 7588
rect 7552 7644 7616 7648
rect 7552 7588 7556 7644
rect 7556 7588 7612 7644
rect 7612 7588 7616 7644
rect 7552 7584 7616 7588
rect 7632 7644 7696 7648
rect 7632 7588 7636 7644
rect 7636 7588 7692 7644
rect 7692 7588 7696 7644
rect 7632 7584 7696 7588
rect 7712 7644 7776 7648
rect 7712 7588 7716 7644
rect 7716 7588 7772 7644
rect 7772 7588 7776 7644
rect 7712 7584 7776 7588
rect 12187 7644 12251 7648
rect 12187 7588 12191 7644
rect 12191 7588 12247 7644
rect 12247 7588 12251 7644
rect 12187 7584 12251 7588
rect 12267 7644 12331 7648
rect 12267 7588 12271 7644
rect 12271 7588 12327 7644
rect 12327 7588 12331 7644
rect 12267 7584 12331 7588
rect 12347 7644 12411 7648
rect 12347 7588 12351 7644
rect 12351 7588 12407 7644
rect 12407 7588 12411 7644
rect 12347 7584 12411 7588
rect 12427 7644 12491 7648
rect 12427 7588 12431 7644
rect 12431 7588 12487 7644
rect 12487 7588 12491 7644
rect 12427 7584 12491 7588
rect 16902 7644 16966 7648
rect 16902 7588 16906 7644
rect 16906 7588 16962 7644
rect 16962 7588 16966 7644
rect 16902 7584 16966 7588
rect 16982 7644 17046 7648
rect 16982 7588 16986 7644
rect 16986 7588 17042 7644
rect 17042 7588 17046 7644
rect 16982 7584 17046 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 5114 7100 5178 7104
rect 5114 7044 5118 7100
rect 5118 7044 5174 7100
rect 5174 7044 5178 7100
rect 5114 7040 5178 7044
rect 5194 7100 5258 7104
rect 5194 7044 5198 7100
rect 5198 7044 5254 7100
rect 5254 7044 5258 7100
rect 5194 7040 5258 7044
rect 5274 7100 5338 7104
rect 5274 7044 5278 7100
rect 5278 7044 5334 7100
rect 5334 7044 5338 7100
rect 5274 7040 5338 7044
rect 5354 7100 5418 7104
rect 5354 7044 5358 7100
rect 5358 7044 5414 7100
rect 5414 7044 5418 7100
rect 5354 7040 5418 7044
rect 9829 7100 9893 7104
rect 9829 7044 9833 7100
rect 9833 7044 9889 7100
rect 9889 7044 9893 7100
rect 9829 7040 9893 7044
rect 9909 7100 9973 7104
rect 9909 7044 9913 7100
rect 9913 7044 9969 7100
rect 9969 7044 9973 7100
rect 9909 7040 9973 7044
rect 9989 7100 10053 7104
rect 9989 7044 9993 7100
rect 9993 7044 10049 7100
rect 10049 7044 10053 7100
rect 9989 7040 10053 7044
rect 10069 7100 10133 7104
rect 10069 7044 10073 7100
rect 10073 7044 10129 7100
rect 10129 7044 10133 7100
rect 10069 7040 10133 7044
rect 14544 7100 14608 7104
rect 14544 7044 14548 7100
rect 14548 7044 14604 7100
rect 14604 7044 14608 7100
rect 14544 7040 14608 7044
rect 14624 7100 14688 7104
rect 14624 7044 14628 7100
rect 14628 7044 14684 7100
rect 14684 7044 14688 7100
rect 14624 7040 14688 7044
rect 14704 7100 14768 7104
rect 14704 7044 14708 7100
rect 14708 7044 14764 7100
rect 14764 7044 14768 7100
rect 14704 7040 14768 7044
rect 14784 7100 14848 7104
rect 14784 7044 14788 7100
rect 14788 7044 14844 7100
rect 14844 7044 14848 7100
rect 14784 7040 14848 7044
rect 19259 7100 19323 7104
rect 19259 7044 19263 7100
rect 19263 7044 19319 7100
rect 19319 7044 19323 7100
rect 19259 7040 19323 7044
rect 19339 7100 19403 7104
rect 19339 7044 19343 7100
rect 19343 7044 19399 7100
rect 19399 7044 19403 7100
rect 19339 7040 19403 7044
rect 19419 7100 19483 7104
rect 19419 7044 19423 7100
rect 19423 7044 19479 7100
rect 19479 7044 19483 7100
rect 19419 7040 19483 7044
rect 19499 7100 19563 7104
rect 19499 7044 19503 7100
rect 19503 7044 19559 7100
rect 19559 7044 19563 7100
rect 19499 7040 19563 7044
rect 11100 6700 11164 6764
rect 2757 6556 2821 6560
rect 2757 6500 2761 6556
rect 2761 6500 2817 6556
rect 2817 6500 2821 6556
rect 2757 6496 2821 6500
rect 2837 6556 2901 6560
rect 2837 6500 2841 6556
rect 2841 6500 2897 6556
rect 2897 6500 2901 6556
rect 2837 6496 2901 6500
rect 2917 6556 2981 6560
rect 2917 6500 2921 6556
rect 2921 6500 2977 6556
rect 2977 6500 2981 6556
rect 2917 6496 2981 6500
rect 2997 6556 3061 6560
rect 2997 6500 3001 6556
rect 3001 6500 3057 6556
rect 3057 6500 3061 6556
rect 2997 6496 3061 6500
rect 7472 6556 7536 6560
rect 7472 6500 7476 6556
rect 7476 6500 7532 6556
rect 7532 6500 7536 6556
rect 7472 6496 7536 6500
rect 7552 6556 7616 6560
rect 7552 6500 7556 6556
rect 7556 6500 7612 6556
rect 7612 6500 7616 6556
rect 7552 6496 7616 6500
rect 7632 6556 7696 6560
rect 7632 6500 7636 6556
rect 7636 6500 7692 6556
rect 7692 6500 7696 6556
rect 7632 6496 7696 6500
rect 7712 6556 7776 6560
rect 7712 6500 7716 6556
rect 7716 6500 7772 6556
rect 7772 6500 7776 6556
rect 7712 6496 7776 6500
rect 12187 6556 12251 6560
rect 12187 6500 12191 6556
rect 12191 6500 12247 6556
rect 12247 6500 12251 6556
rect 12187 6496 12251 6500
rect 12267 6556 12331 6560
rect 12267 6500 12271 6556
rect 12271 6500 12327 6556
rect 12327 6500 12331 6556
rect 12267 6496 12331 6500
rect 12347 6556 12411 6560
rect 12347 6500 12351 6556
rect 12351 6500 12407 6556
rect 12407 6500 12411 6556
rect 12347 6496 12411 6500
rect 12427 6556 12491 6560
rect 12427 6500 12431 6556
rect 12431 6500 12487 6556
rect 12487 6500 12491 6556
rect 12427 6496 12491 6500
rect 16902 6556 16966 6560
rect 16902 6500 16906 6556
rect 16906 6500 16962 6556
rect 16962 6500 16966 6556
rect 16902 6496 16966 6500
rect 16982 6556 17046 6560
rect 16982 6500 16986 6556
rect 16986 6500 17042 6556
rect 17042 6500 17046 6556
rect 16982 6496 17046 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 5114 6012 5178 6016
rect 5114 5956 5118 6012
rect 5118 5956 5174 6012
rect 5174 5956 5178 6012
rect 5114 5952 5178 5956
rect 5194 6012 5258 6016
rect 5194 5956 5198 6012
rect 5198 5956 5254 6012
rect 5254 5956 5258 6012
rect 5194 5952 5258 5956
rect 5274 6012 5338 6016
rect 5274 5956 5278 6012
rect 5278 5956 5334 6012
rect 5334 5956 5338 6012
rect 5274 5952 5338 5956
rect 5354 6012 5418 6016
rect 5354 5956 5358 6012
rect 5358 5956 5414 6012
rect 5414 5956 5418 6012
rect 5354 5952 5418 5956
rect 9829 6012 9893 6016
rect 9829 5956 9833 6012
rect 9833 5956 9889 6012
rect 9889 5956 9893 6012
rect 9829 5952 9893 5956
rect 9909 6012 9973 6016
rect 9909 5956 9913 6012
rect 9913 5956 9969 6012
rect 9969 5956 9973 6012
rect 9909 5952 9973 5956
rect 9989 6012 10053 6016
rect 9989 5956 9993 6012
rect 9993 5956 10049 6012
rect 10049 5956 10053 6012
rect 9989 5952 10053 5956
rect 10069 6012 10133 6016
rect 10069 5956 10073 6012
rect 10073 5956 10129 6012
rect 10129 5956 10133 6012
rect 10069 5952 10133 5956
rect 14544 6012 14608 6016
rect 14544 5956 14548 6012
rect 14548 5956 14604 6012
rect 14604 5956 14608 6012
rect 14544 5952 14608 5956
rect 14624 6012 14688 6016
rect 14624 5956 14628 6012
rect 14628 5956 14684 6012
rect 14684 5956 14688 6012
rect 14624 5952 14688 5956
rect 14704 6012 14768 6016
rect 14704 5956 14708 6012
rect 14708 5956 14764 6012
rect 14764 5956 14768 6012
rect 14704 5952 14768 5956
rect 14784 6012 14848 6016
rect 14784 5956 14788 6012
rect 14788 5956 14844 6012
rect 14844 5956 14848 6012
rect 14784 5952 14848 5956
rect 19259 6012 19323 6016
rect 19259 5956 19263 6012
rect 19263 5956 19319 6012
rect 19319 5956 19323 6012
rect 19259 5952 19323 5956
rect 19339 6012 19403 6016
rect 19339 5956 19343 6012
rect 19343 5956 19399 6012
rect 19399 5956 19403 6012
rect 19339 5952 19403 5956
rect 19419 6012 19483 6016
rect 19419 5956 19423 6012
rect 19423 5956 19479 6012
rect 19479 5956 19483 6012
rect 19419 5952 19483 5956
rect 19499 6012 19563 6016
rect 19499 5956 19503 6012
rect 19503 5956 19559 6012
rect 19559 5956 19563 6012
rect 19499 5952 19563 5956
rect 2757 5468 2821 5472
rect 2757 5412 2761 5468
rect 2761 5412 2817 5468
rect 2817 5412 2821 5468
rect 2757 5408 2821 5412
rect 2837 5468 2901 5472
rect 2837 5412 2841 5468
rect 2841 5412 2897 5468
rect 2897 5412 2901 5468
rect 2837 5408 2901 5412
rect 2917 5468 2981 5472
rect 2917 5412 2921 5468
rect 2921 5412 2977 5468
rect 2977 5412 2981 5468
rect 2917 5408 2981 5412
rect 2997 5468 3061 5472
rect 2997 5412 3001 5468
rect 3001 5412 3057 5468
rect 3057 5412 3061 5468
rect 2997 5408 3061 5412
rect 7472 5468 7536 5472
rect 7472 5412 7476 5468
rect 7476 5412 7532 5468
rect 7532 5412 7536 5468
rect 7472 5408 7536 5412
rect 7552 5468 7616 5472
rect 7552 5412 7556 5468
rect 7556 5412 7612 5468
rect 7612 5412 7616 5468
rect 7552 5408 7616 5412
rect 7632 5468 7696 5472
rect 7632 5412 7636 5468
rect 7636 5412 7692 5468
rect 7692 5412 7696 5468
rect 7632 5408 7696 5412
rect 7712 5468 7776 5472
rect 7712 5412 7716 5468
rect 7716 5412 7772 5468
rect 7772 5412 7776 5468
rect 7712 5408 7776 5412
rect 12187 5468 12251 5472
rect 12187 5412 12191 5468
rect 12191 5412 12247 5468
rect 12247 5412 12251 5468
rect 12187 5408 12251 5412
rect 12267 5468 12331 5472
rect 12267 5412 12271 5468
rect 12271 5412 12327 5468
rect 12327 5412 12331 5468
rect 12267 5408 12331 5412
rect 12347 5468 12411 5472
rect 12347 5412 12351 5468
rect 12351 5412 12407 5468
rect 12407 5412 12411 5468
rect 12347 5408 12411 5412
rect 12427 5468 12491 5472
rect 12427 5412 12431 5468
rect 12431 5412 12487 5468
rect 12487 5412 12491 5468
rect 12427 5408 12491 5412
rect 16902 5468 16966 5472
rect 16902 5412 16906 5468
rect 16906 5412 16962 5468
rect 16962 5412 16966 5468
rect 16902 5408 16966 5412
rect 16982 5468 17046 5472
rect 16982 5412 16986 5468
rect 16986 5412 17042 5468
rect 17042 5412 17046 5468
rect 16982 5408 17046 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 9628 5068 9692 5132
rect 5114 4924 5178 4928
rect 5114 4868 5118 4924
rect 5118 4868 5174 4924
rect 5174 4868 5178 4924
rect 5114 4864 5178 4868
rect 5194 4924 5258 4928
rect 5194 4868 5198 4924
rect 5198 4868 5254 4924
rect 5254 4868 5258 4924
rect 5194 4864 5258 4868
rect 5274 4924 5338 4928
rect 5274 4868 5278 4924
rect 5278 4868 5334 4924
rect 5334 4868 5338 4924
rect 5274 4864 5338 4868
rect 5354 4924 5418 4928
rect 5354 4868 5358 4924
rect 5358 4868 5414 4924
rect 5414 4868 5418 4924
rect 5354 4864 5418 4868
rect 9829 4924 9893 4928
rect 9829 4868 9833 4924
rect 9833 4868 9889 4924
rect 9889 4868 9893 4924
rect 9829 4864 9893 4868
rect 9909 4924 9973 4928
rect 9909 4868 9913 4924
rect 9913 4868 9969 4924
rect 9969 4868 9973 4924
rect 9909 4864 9973 4868
rect 9989 4924 10053 4928
rect 9989 4868 9993 4924
rect 9993 4868 10049 4924
rect 10049 4868 10053 4924
rect 9989 4864 10053 4868
rect 10069 4924 10133 4928
rect 10069 4868 10073 4924
rect 10073 4868 10129 4924
rect 10129 4868 10133 4924
rect 10069 4864 10133 4868
rect 14544 4924 14608 4928
rect 14544 4868 14548 4924
rect 14548 4868 14604 4924
rect 14604 4868 14608 4924
rect 14544 4864 14608 4868
rect 14624 4924 14688 4928
rect 14624 4868 14628 4924
rect 14628 4868 14684 4924
rect 14684 4868 14688 4924
rect 14624 4864 14688 4868
rect 14704 4924 14768 4928
rect 14704 4868 14708 4924
rect 14708 4868 14764 4924
rect 14764 4868 14768 4924
rect 14704 4864 14768 4868
rect 14784 4924 14848 4928
rect 14784 4868 14788 4924
rect 14788 4868 14844 4924
rect 14844 4868 14848 4924
rect 14784 4864 14848 4868
rect 19259 4924 19323 4928
rect 19259 4868 19263 4924
rect 19263 4868 19319 4924
rect 19319 4868 19323 4924
rect 19259 4864 19323 4868
rect 19339 4924 19403 4928
rect 19339 4868 19343 4924
rect 19343 4868 19399 4924
rect 19399 4868 19403 4924
rect 19339 4864 19403 4868
rect 19419 4924 19483 4928
rect 19419 4868 19423 4924
rect 19423 4868 19479 4924
rect 19479 4868 19483 4924
rect 19419 4864 19483 4868
rect 19499 4924 19563 4928
rect 19499 4868 19503 4924
rect 19503 4868 19559 4924
rect 19559 4868 19563 4924
rect 19499 4864 19563 4868
rect 2757 4380 2821 4384
rect 2757 4324 2761 4380
rect 2761 4324 2817 4380
rect 2817 4324 2821 4380
rect 2757 4320 2821 4324
rect 2837 4380 2901 4384
rect 2837 4324 2841 4380
rect 2841 4324 2897 4380
rect 2897 4324 2901 4380
rect 2837 4320 2901 4324
rect 2917 4380 2981 4384
rect 2917 4324 2921 4380
rect 2921 4324 2977 4380
rect 2977 4324 2981 4380
rect 2917 4320 2981 4324
rect 2997 4380 3061 4384
rect 2997 4324 3001 4380
rect 3001 4324 3057 4380
rect 3057 4324 3061 4380
rect 2997 4320 3061 4324
rect 7472 4380 7536 4384
rect 7472 4324 7476 4380
rect 7476 4324 7532 4380
rect 7532 4324 7536 4380
rect 7472 4320 7536 4324
rect 7552 4380 7616 4384
rect 7552 4324 7556 4380
rect 7556 4324 7612 4380
rect 7612 4324 7616 4380
rect 7552 4320 7616 4324
rect 7632 4380 7696 4384
rect 7632 4324 7636 4380
rect 7636 4324 7692 4380
rect 7692 4324 7696 4380
rect 7632 4320 7696 4324
rect 7712 4380 7776 4384
rect 7712 4324 7716 4380
rect 7716 4324 7772 4380
rect 7772 4324 7776 4380
rect 7712 4320 7776 4324
rect 12187 4380 12251 4384
rect 12187 4324 12191 4380
rect 12191 4324 12247 4380
rect 12247 4324 12251 4380
rect 12187 4320 12251 4324
rect 12267 4380 12331 4384
rect 12267 4324 12271 4380
rect 12271 4324 12327 4380
rect 12327 4324 12331 4380
rect 12267 4320 12331 4324
rect 12347 4380 12411 4384
rect 12347 4324 12351 4380
rect 12351 4324 12407 4380
rect 12407 4324 12411 4380
rect 12347 4320 12411 4324
rect 12427 4380 12491 4384
rect 12427 4324 12431 4380
rect 12431 4324 12487 4380
rect 12487 4324 12491 4380
rect 12427 4320 12491 4324
rect 16902 4380 16966 4384
rect 16902 4324 16906 4380
rect 16906 4324 16962 4380
rect 16962 4324 16966 4380
rect 16902 4320 16966 4324
rect 16982 4380 17046 4384
rect 16982 4324 16986 4380
rect 16986 4324 17042 4380
rect 17042 4324 17046 4380
rect 16982 4320 17046 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 5114 3836 5178 3840
rect 5114 3780 5118 3836
rect 5118 3780 5174 3836
rect 5174 3780 5178 3836
rect 5114 3776 5178 3780
rect 5194 3836 5258 3840
rect 5194 3780 5198 3836
rect 5198 3780 5254 3836
rect 5254 3780 5258 3836
rect 5194 3776 5258 3780
rect 5274 3836 5338 3840
rect 5274 3780 5278 3836
rect 5278 3780 5334 3836
rect 5334 3780 5338 3836
rect 5274 3776 5338 3780
rect 5354 3836 5418 3840
rect 5354 3780 5358 3836
rect 5358 3780 5414 3836
rect 5414 3780 5418 3836
rect 5354 3776 5418 3780
rect 9829 3836 9893 3840
rect 9829 3780 9833 3836
rect 9833 3780 9889 3836
rect 9889 3780 9893 3836
rect 9829 3776 9893 3780
rect 9909 3836 9973 3840
rect 9909 3780 9913 3836
rect 9913 3780 9969 3836
rect 9969 3780 9973 3836
rect 9909 3776 9973 3780
rect 9989 3836 10053 3840
rect 9989 3780 9993 3836
rect 9993 3780 10049 3836
rect 10049 3780 10053 3836
rect 9989 3776 10053 3780
rect 10069 3836 10133 3840
rect 10069 3780 10073 3836
rect 10073 3780 10129 3836
rect 10129 3780 10133 3836
rect 10069 3776 10133 3780
rect 14544 3836 14608 3840
rect 14544 3780 14548 3836
rect 14548 3780 14604 3836
rect 14604 3780 14608 3836
rect 14544 3776 14608 3780
rect 14624 3836 14688 3840
rect 14624 3780 14628 3836
rect 14628 3780 14684 3836
rect 14684 3780 14688 3836
rect 14624 3776 14688 3780
rect 14704 3836 14768 3840
rect 14704 3780 14708 3836
rect 14708 3780 14764 3836
rect 14764 3780 14768 3836
rect 14704 3776 14768 3780
rect 14784 3836 14848 3840
rect 14784 3780 14788 3836
rect 14788 3780 14844 3836
rect 14844 3780 14848 3836
rect 14784 3776 14848 3780
rect 19259 3836 19323 3840
rect 19259 3780 19263 3836
rect 19263 3780 19319 3836
rect 19319 3780 19323 3836
rect 19259 3776 19323 3780
rect 19339 3836 19403 3840
rect 19339 3780 19343 3836
rect 19343 3780 19399 3836
rect 19399 3780 19403 3836
rect 19339 3776 19403 3780
rect 19419 3836 19483 3840
rect 19419 3780 19423 3836
rect 19423 3780 19479 3836
rect 19479 3780 19483 3836
rect 19419 3776 19483 3780
rect 19499 3836 19563 3840
rect 19499 3780 19503 3836
rect 19503 3780 19559 3836
rect 19559 3780 19563 3836
rect 19499 3776 19563 3780
rect 2757 3292 2821 3296
rect 2757 3236 2761 3292
rect 2761 3236 2817 3292
rect 2817 3236 2821 3292
rect 2757 3232 2821 3236
rect 2837 3292 2901 3296
rect 2837 3236 2841 3292
rect 2841 3236 2897 3292
rect 2897 3236 2901 3292
rect 2837 3232 2901 3236
rect 2917 3292 2981 3296
rect 2917 3236 2921 3292
rect 2921 3236 2977 3292
rect 2977 3236 2981 3292
rect 2917 3232 2981 3236
rect 2997 3292 3061 3296
rect 2997 3236 3001 3292
rect 3001 3236 3057 3292
rect 3057 3236 3061 3292
rect 2997 3232 3061 3236
rect 7472 3292 7536 3296
rect 7472 3236 7476 3292
rect 7476 3236 7532 3292
rect 7532 3236 7536 3292
rect 7472 3232 7536 3236
rect 7552 3292 7616 3296
rect 7552 3236 7556 3292
rect 7556 3236 7612 3292
rect 7612 3236 7616 3292
rect 7552 3232 7616 3236
rect 7632 3292 7696 3296
rect 7632 3236 7636 3292
rect 7636 3236 7692 3292
rect 7692 3236 7696 3292
rect 7632 3232 7696 3236
rect 7712 3292 7776 3296
rect 7712 3236 7716 3292
rect 7716 3236 7772 3292
rect 7772 3236 7776 3292
rect 7712 3232 7776 3236
rect 12187 3292 12251 3296
rect 12187 3236 12191 3292
rect 12191 3236 12247 3292
rect 12247 3236 12251 3292
rect 12187 3232 12251 3236
rect 12267 3292 12331 3296
rect 12267 3236 12271 3292
rect 12271 3236 12327 3292
rect 12327 3236 12331 3292
rect 12267 3232 12331 3236
rect 12347 3292 12411 3296
rect 12347 3236 12351 3292
rect 12351 3236 12407 3292
rect 12407 3236 12411 3292
rect 12347 3232 12411 3236
rect 12427 3292 12491 3296
rect 12427 3236 12431 3292
rect 12431 3236 12487 3292
rect 12487 3236 12491 3292
rect 12427 3232 12491 3236
rect 16902 3292 16966 3296
rect 16902 3236 16906 3292
rect 16906 3236 16962 3292
rect 16962 3236 16966 3292
rect 16902 3232 16966 3236
rect 16982 3292 17046 3296
rect 16982 3236 16986 3292
rect 16986 3236 17042 3292
rect 17042 3236 17046 3292
rect 16982 3232 17046 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 5114 2748 5178 2752
rect 5114 2692 5118 2748
rect 5118 2692 5174 2748
rect 5174 2692 5178 2748
rect 5114 2688 5178 2692
rect 5194 2748 5258 2752
rect 5194 2692 5198 2748
rect 5198 2692 5254 2748
rect 5254 2692 5258 2748
rect 5194 2688 5258 2692
rect 5274 2748 5338 2752
rect 5274 2692 5278 2748
rect 5278 2692 5334 2748
rect 5334 2692 5338 2748
rect 5274 2688 5338 2692
rect 5354 2748 5418 2752
rect 5354 2692 5358 2748
rect 5358 2692 5414 2748
rect 5414 2692 5418 2748
rect 5354 2688 5418 2692
rect 9829 2748 9893 2752
rect 9829 2692 9833 2748
rect 9833 2692 9889 2748
rect 9889 2692 9893 2748
rect 9829 2688 9893 2692
rect 9909 2748 9973 2752
rect 9909 2692 9913 2748
rect 9913 2692 9969 2748
rect 9969 2692 9973 2748
rect 9909 2688 9973 2692
rect 9989 2748 10053 2752
rect 9989 2692 9993 2748
rect 9993 2692 10049 2748
rect 10049 2692 10053 2748
rect 9989 2688 10053 2692
rect 10069 2748 10133 2752
rect 10069 2692 10073 2748
rect 10073 2692 10129 2748
rect 10129 2692 10133 2748
rect 10069 2688 10133 2692
rect 14544 2748 14608 2752
rect 14544 2692 14548 2748
rect 14548 2692 14604 2748
rect 14604 2692 14608 2748
rect 14544 2688 14608 2692
rect 14624 2748 14688 2752
rect 14624 2692 14628 2748
rect 14628 2692 14684 2748
rect 14684 2692 14688 2748
rect 14624 2688 14688 2692
rect 14704 2748 14768 2752
rect 14704 2692 14708 2748
rect 14708 2692 14764 2748
rect 14764 2692 14768 2748
rect 14704 2688 14768 2692
rect 14784 2748 14848 2752
rect 14784 2692 14788 2748
rect 14788 2692 14844 2748
rect 14844 2692 14848 2748
rect 14784 2688 14848 2692
rect 19259 2748 19323 2752
rect 19259 2692 19263 2748
rect 19263 2692 19319 2748
rect 19319 2692 19323 2748
rect 19259 2688 19323 2692
rect 19339 2748 19403 2752
rect 19339 2692 19343 2748
rect 19343 2692 19399 2748
rect 19399 2692 19403 2748
rect 19339 2688 19403 2692
rect 19419 2748 19483 2752
rect 19419 2692 19423 2748
rect 19423 2692 19479 2748
rect 19479 2692 19483 2748
rect 19419 2688 19483 2692
rect 19499 2748 19563 2752
rect 19499 2692 19503 2748
rect 19503 2692 19559 2748
rect 19559 2692 19563 2748
rect 19499 2688 19563 2692
rect 10732 2620 10796 2684
rect 11468 2620 11532 2684
rect 2757 2204 2821 2208
rect 2757 2148 2761 2204
rect 2761 2148 2817 2204
rect 2817 2148 2821 2204
rect 2757 2144 2821 2148
rect 2837 2204 2901 2208
rect 2837 2148 2841 2204
rect 2841 2148 2897 2204
rect 2897 2148 2901 2204
rect 2837 2144 2901 2148
rect 2917 2204 2981 2208
rect 2917 2148 2921 2204
rect 2921 2148 2977 2204
rect 2977 2148 2981 2204
rect 2917 2144 2981 2148
rect 2997 2204 3061 2208
rect 2997 2148 3001 2204
rect 3001 2148 3057 2204
rect 3057 2148 3061 2204
rect 2997 2144 3061 2148
rect 7472 2204 7536 2208
rect 7472 2148 7476 2204
rect 7476 2148 7532 2204
rect 7532 2148 7536 2204
rect 7472 2144 7536 2148
rect 7552 2204 7616 2208
rect 7552 2148 7556 2204
rect 7556 2148 7612 2204
rect 7612 2148 7616 2204
rect 7552 2144 7616 2148
rect 7632 2204 7696 2208
rect 7632 2148 7636 2204
rect 7636 2148 7692 2204
rect 7692 2148 7696 2204
rect 7632 2144 7696 2148
rect 7712 2204 7776 2208
rect 7712 2148 7716 2204
rect 7716 2148 7772 2204
rect 7772 2148 7776 2204
rect 7712 2144 7776 2148
rect 12187 2204 12251 2208
rect 12187 2148 12191 2204
rect 12191 2148 12247 2204
rect 12247 2148 12251 2204
rect 12187 2144 12251 2148
rect 12267 2204 12331 2208
rect 12267 2148 12271 2204
rect 12271 2148 12327 2204
rect 12327 2148 12331 2204
rect 12267 2144 12331 2148
rect 12347 2204 12411 2208
rect 12347 2148 12351 2204
rect 12351 2148 12407 2204
rect 12407 2148 12411 2204
rect 12347 2144 12411 2148
rect 12427 2204 12491 2208
rect 12427 2148 12431 2204
rect 12431 2148 12487 2204
rect 12487 2148 12491 2204
rect 12427 2144 12491 2148
rect 16902 2204 16966 2208
rect 16902 2148 16906 2204
rect 16906 2148 16962 2204
rect 16962 2148 16966 2204
rect 16902 2144 16966 2148
rect 16982 2204 17046 2208
rect 16982 2148 16986 2204
rect 16986 2148 17042 2204
rect 17042 2148 17046 2204
rect 16982 2144 17046 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 5114 1660 5178 1664
rect 5114 1604 5118 1660
rect 5118 1604 5174 1660
rect 5174 1604 5178 1660
rect 5114 1600 5178 1604
rect 5194 1660 5258 1664
rect 5194 1604 5198 1660
rect 5198 1604 5254 1660
rect 5254 1604 5258 1660
rect 5194 1600 5258 1604
rect 5274 1660 5338 1664
rect 5274 1604 5278 1660
rect 5278 1604 5334 1660
rect 5334 1604 5338 1660
rect 5274 1600 5338 1604
rect 5354 1660 5418 1664
rect 5354 1604 5358 1660
rect 5358 1604 5414 1660
rect 5414 1604 5418 1660
rect 5354 1600 5418 1604
rect 9829 1660 9893 1664
rect 9829 1604 9833 1660
rect 9833 1604 9889 1660
rect 9889 1604 9893 1660
rect 9829 1600 9893 1604
rect 9909 1660 9973 1664
rect 9909 1604 9913 1660
rect 9913 1604 9969 1660
rect 9969 1604 9973 1660
rect 9909 1600 9973 1604
rect 9989 1660 10053 1664
rect 9989 1604 9993 1660
rect 9993 1604 10049 1660
rect 10049 1604 10053 1660
rect 9989 1600 10053 1604
rect 10069 1660 10133 1664
rect 10069 1604 10073 1660
rect 10073 1604 10129 1660
rect 10129 1604 10133 1660
rect 10069 1600 10133 1604
rect 14544 1660 14608 1664
rect 14544 1604 14548 1660
rect 14548 1604 14604 1660
rect 14604 1604 14608 1660
rect 14544 1600 14608 1604
rect 14624 1660 14688 1664
rect 14624 1604 14628 1660
rect 14628 1604 14684 1660
rect 14684 1604 14688 1660
rect 14624 1600 14688 1604
rect 14704 1660 14768 1664
rect 14704 1604 14708 1660
rect 14708 1604 14764 1660
rect 14764 1604 14768 1660
rect 14704 1600 14768 1604
rect 14784 1660 14848 1664
rect 14784 1604 14788 1660
rect 14788 1604 14844 1660
rect 14844 1604 14848 1660
rect 14784 1600 14848 1604
rect 19259 1660 19323 1664
rect 19259 1604 19263 1660
rect 19263 1604 19319 1660
rect 19319 1604 19323 1660
rect 19259 1600 19323 1604
rect 19339 1660 19403 1664
rect 19339 1604 19343 1660
rect 19343 1604 19399 1660
rect 19399 1604 19403 1660
rect 19339 1600 19403 1604
rect 19419 1660 19483 1664
rect 19419 1604 19423 1660
rect 19423 1604 19479 1660
rect 19479 1604 19483 1660
rect 19419 1600 19483 1604
rect 19499 1660 19563 1664
rect 19499 1604 19503 1660
rect 19503 1604 19559 1660
rect 19559 1604 19563 1660
rect 19499 1600 19563 1604
rect 2757 1116 2821 1120
rect 2757 1060 2761 1116
rect 2761 1060 2817 1116
rect 2817 1060 2821 1116
rect 2757 1056 2821 1060
rect 2837 1116 2901 1120
rect 2837 1060 2841 1116
rect 2841 1060 2897 1116
rect 2897 1060 2901 1116
rect 2837 1056 2901 1060
rect 2917 1116 2981 1120
rect 2917 1060 2921 1116
rect 2921 1060 2977 1116
rect 2977 1060 2981 1116
rect 2917 1056 2981 1060
rect 2997 1116 3061 1120
rect 2997 1060 3001 1116
rect 3001 1060 3057 1116
rect 3057 1060 3061 1116
rect 2997 1056 3061 1060
rect 7472 1116 7536 1120
rect 7472 1060 7476 1116
rect 7476 1060 7532 1116
rect 7532 1060 7536 1116
rect 7472 1056 7536 1060
rect 7552 1116 7616 1120
rect 7552 1060 7556 1116
rect 7556 1060 7612 1116
rect 7612 1060 7616 1116
rect 7552 1056 7616 1060
rect 7632 1116 7696 1120
rect 7632 1060 7636 1116
rect 7636 1060 7692 1116
rect 7692 1060 7696 1116
rect 7632 1056 7696 1060
rect 7712 1116 7776 1120
rect 7712 1060 7716 1116
rect 7716 1060 7772 1116
rect 7772 1060 7776 1116
rect 7712 1056 7776 1060
rect 12187 1116 12251 1120
rect 12187 1060 12191 1116
rect 12191 1060 12247 1116
rect 12247 1060 12251 1116
rect 12187 1056 12251 1060
rect 12267 1116 12331 1120
rect 12267 1060 12271 1116
rect 12271 1060 12327 1116
rect 12327 1060 12331 1116
rect 12267 1056 12331 1060
rect 12347 1116 12411 1120
rect 12347 1060 12351 1116
rect 12351 1060 12407 1116
rect 12407 1060 12411 1116
rect 12347 1056 12411 1060
rect 12427 1116 12491 1120
rect 12427 1060 12431 1116
rect 12431 1060 12487 1116
rect 12487 1060 12491 1116
rect 12427 1056 12491 1060
rect 16902 1116 16966 1120
rect 16902 1060 16906 1116
rect 16906 1060 16962 1116
rect 16962 1060 16966 1116
rect 16902 1056 16966 1060
rect 16982 1116 17046 1120
rect 16982 1060 16986 1116
rect 16986 1060 17042 1116
rect 17042 1060 17046 1116
rect 16982 1056 17046 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 5114 572 5178 576
rect 5114 516 5118 572
rect 5118 516 5174 572
rect 5174 516 5178 572
rect 5114 512 5178 516
rect 5194 572 5258 576
rect 5194 516 5198 572
rect 5198 516 5254 572
rect 5254 516 5258 572
rect 5194 512 5258 516
rect 5274 572 5338 576
rect 5274 516 5278 572
rect 5278 516 5334 572
rect 5334 516 5338 572
rect 5274 512 5338 516
rect 5354 572 5418 576
rect 5354 516 5358 572
rect 5358 516 5414 572
rect 5414 516 5418 572
rect 5354 512 5418 516
rect 9829 572 9893 576
rect 9829 516 9833 572
rect 9833 516 9889 572
rect 9889 516 9893 572
rect 9829 512 9893 516
rect 9909 572 9973 576
rect 9909 516 9913 572
rect 9913 516 9969 572
rect 9969 516 9973 572
rect 9909 512 9973 516
rect 9989 572 10053 576
rect 9989 516 9993 572
rect 9993 516 10049 572
rect 10049 516 10053 572
rect 9989 512 10053 516
rect 10069 572 10133 576
rect 10069 516 10073 572
rect 10073 516 10129 572
rect 10129 516 10133 572
rect 10069 512 10133 516
rect 14544 572 14608 576
rect 14544 516 14548 572
rect 14548 516 14604 572
rect 14604 516 14608 572
rect 14544 512 14608 516
rect 14624 572 14688 576
rect 14624 516 14628 572
rect 14628 516 14684 572
rect 14684 516 14688 572
rect 14624 512 14688 516
rect 14704 572 14768 576
rect 14704 516 14708 572
rect 14708 516 14764 572
rect 14764 516 14768 572
rect 14704 512 14768 516
rect 14784 572 14848 576
rect 14784 516 14788 572
rect 14788 516 14844 572
rect 14844 516 14848 572
rect 14784 512 14848 516
rect 19259 572 19323 576
rect 19259 516 19263 572
rect 19263 516 19319 572
rect 19319 516 19323 572
rect 19259 512 19323 516
rect 19339 572 19403 576
rect 19339 516 19343 572
rect 19343 516 19399 572
rect 19399 516 19403 572
rect 19339 512 19403 516
rect 19419 572 19483 576
rect 19419 516 19423 572
rect 19423 516 19479 572
rect 19479 516 19483 572
rect 19419 512 19483 516
rect 19499 572 19563 576
rect 19499 516 19503 572
rect 19503 516 19559 572
rect 19559 516 19563 572
rect 19499 512 19563 516
<< metal4 >>
rect 2749 18528 3069 19088
rect 2749 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3069 18528
rect 2749 17440 3069 18464
rect 2749 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3069 17440
rect 2749 16352 3069 17376
rect 2749 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3069 16352
rect 2749 15264 3069 16288
rect 2749 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3069 15264
rect 2749 14176 3069 15200
rect 2749 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3069 14176
rect 2749 13088 3069 14112
rect 2749 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3069 13088
rect 2749 12000 3069 13024
rect 2749 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3069 12000
rect 2749 10912 3069 11936
rect 2749 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3069 10912
rect 2749 9824 3069 10848
rect 2749 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3069 9824
rect 2749 8736 3069 9760
rect 2749 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3069 8736
rect 2749 7648 3069 8672
rect 2749 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3069 7648
rect 2749 6560 3069 7584
rect 2749 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3069 6560
rect 2749 5472 3069 6496
rect 2749 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3069 5472
rect 2749 4384 3069 5408
rect 2749 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3069 4384
rect 2749 3296 3069 4320
rect 2749 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3069 3296
rect 2749 2208 3069 3232
rect 2749 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3069 2208
rect 2749 1120 3069 2144
rect 2749 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3069 1120
rect 2749 496 3069 1056
rect 5106 19072 5426 19088
rect 5106 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5426 19072
rect 5106 17984 5426 19008
rect 5106 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5426 17984
rect 5106 16896 5426 17920
rect 5106 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5426 16896
rect 5106 15808 5426 16832
rect 5106 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5426 15808
rect 5106 14720 5426 15744
rect 5106 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5426 14720
rect 5106 13632 5426 14656
rect 5106 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5426 13632
rect 5106 12544 5426 13568
rect 5106 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5426 12544
rect 5106 11456 5426 12480
rect 5106 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5426 11456
rect 5106 10368 5426 11392
rect 5106 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5426 10368
rect 5106 9280 5426 10304
rect 5106 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5426 9280
rect 5106 8192 5426 9216
rect 5106 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5426 8192
rect 5106 7104 5426 8128
rect 5106 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5426 7104
rect 5106 6016 5426 7040
rect 5106 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5426 6016
rect 5106 4928 5426 5952
rect 5106 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5426 4928
rect 5106 3840 5426 4864
rect 5106 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5426 3840
rect 5106 2752 5426 3776
rect 5106 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5426 2752
rect 5106 1664 5426 2688
rect 5106 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5426 1664
rect 5106 576 5426 1600
rect 5106 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5426 576
rect 5106 496 5426 512
rect 7464 18528 7784 19088
rect 7464 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7784 18528
rect 7464 17440 7784 18464
rect 7464 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7784 17440
rect 7464 16352 7784 17376
rect 7464 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7784 16352
rect 7464 15264 7784 16288
rect 7464 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7784 15264
rect 7464 14176 7784 15200
rect 7464 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7784 14176
rect 7464 13088 7784 14112
rect 7464 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7784 13088
rect 7464 12000 7784 13024
rect 7464 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7784 12000
rect 7464 10912 7784 11936
rect 9821 19072 10141 19088
rect 9821 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10141 19072
rect 9821 17984 10141 19008
rect 9821 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10141 17984
rect 9821 16896 10141 17920
rect 9821 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10141 16896
rect 9821 15808 10141 16832
rect 9821 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10141 15808
rect 9821 14720 10141 15744
rect 9821 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10141 14720
rect 9821 13632 10141 14656
rect 9821 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10141 13632
rect 9821 12544 10141 13568
rect 12179 18528 12499 19088
rect 12179 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12499 18528
rect 12179 17440 12499 18464
rect 12179 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12499 17440
rect 12179 16352 12499 17376
rect 12179 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12499 16352
rect 12179 15264 12499 16288
rect 12179 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12499 15264
rect 12179 14176 12499 15200
rect 12179 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12499 14176
rect 12179 13088 12499 14112
rect 12179 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12499 13088
rect 10731 12612 10797 12613
rect 10731 12548 10732 12612
rect 10796 12548 10797 12612
rect 10731 12547 10797 12548
rect 9821 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10141 12544
rect 9627 11660 9693 11661
rect 9627 11596 9628 11660
rect 9692 11596 9693 11660
rect 9627 11595 9693 11596
rect 7464 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7784 10912
rect 7464 9824 7784 10848
rect 7464 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7784 9824
rect 7464 8736 7784 9760
rect 7464 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7784 8736
rect 7464 7648 7784 8672
rect 7464 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7784 7648
rect 7464 6560 7784 7584
rect 7464 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7784 6560
rect 7464 5472 7784 6496
rect 7464 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7784 5472
rect 7464 4384 7784 5408
rect 9630 5133 9690 11595
rect 9821 11456 10141 12480
rect 9821 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10141 11456
rect 9821 10368 10141 11392
rect 9821 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10141 10368
rect 9821 9280 10141 10304
rect 9821 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10141 9280
rect 9821 8192 10141 9216
rect 9821 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10141 8192
rect 9821 7104 10141 8128
rect 9821 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10141 7104
rect 9821 6016 10141 7040
rect 9821 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10141 6016
rect 9627 5132 9693 5133
rect 9627 5068 9628 5132
rect 9692 5068 9693 5132
rect 9627 5067 9693 5068
rect 7464 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7784 4384
rect 7464 3296 7784 4320
rect 7464 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7784 3296
rect 7464 2208 7784 3232
rect 7464 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7784 2208
rect 7464 1120 7784 2144
rect 7464 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7784 1120
rect 7464 496 7784 1056
rect 9821 4928 10141 5952
rect 9821 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10141 4928
rect 9821 3840 10141 4864
rect 9821 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10141 3840
rect 9821 2752 10141 3776
rect 9821 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10141 2752
rect 9821 1664 10141 2688
rect 10734 2685 10794 12547
rect 12179 12000 12499 13024
rect 12179 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12499 12000
rect 12179 10912 12499 11936
rect 12179 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12499 10912
rect 12179 9824 12499 10848
rect 12179 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12499 9824
rect 11467 9756 11533 9757
rect 11467 9692 11468 9756
rect 11532 9692 11533 9756
rect 11467 9691 11533 9692
rect 11099 8260 11165 8261
rect 11099 8196 11100 8260
rect 11164 8196 11165 8260
rect 11099 8195 11165 8196
rect 11102 6765 11162 8195
rect 11099 6764 11165 6765
rect 11099 6700 11100 6764
rect 11164 6700 11165 6764
rect 11099 6699 11165 6700
rect 11470 2685 11530 9691
rect 12179 8736 12499 9760
rect 12179 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12499 8736
rect 12179 7648 12499 8672
rect 12179 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12499 7648
rect 12179 6560 12499 7584
rect 12179 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12499 6560
rect 12179 5472 12499 6496
rect 12179 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12499 5472
rect 12179 4384 12499 5408
rect 12179 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12499 4384
rect 12179 3296 12499 4320
rect 12179 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12499 3296
rect 10731 2684 10797 2685
rect 10731 2620 10732 2684
rect 10796 2620 10797 2684
rect 10731 2619 10797 2620
rect 11467 2684 11533 2685
rect 11467 2620 11468 2684
rect 11532 2620 11533 2684
rect 11467 2619 11533 2620
rect 9821 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10141 1664
rect 9821 576 10141 1600
rect 9821 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10141 576
rect 9821 496 10141 512
rect 12179 2208 12499 3232
rect 12179 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12499 2208
rect 12179 1120 12499 2144
rect 12179 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12499 1120
rect 12179 496 12499 1056
rect 14536 19072 14856 19088
rect 14536 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14856 19072
rect 14536 17984 14856 19008
rect 14536 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14856 17984
rect 14536 16896 14856 17920
rect 14536 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14856 16896
rect 14536 15808 14856 16832
rect 14536 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14856 15808
rect 14536 14720 14856 15744
rect 14536 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14856 14720
rect 14536 13632 14856 14656
rect 14536 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14856 13632
rect 14536 12544 14856 13568
rect 14536 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14856 12544
rect 14536 11456 14856 12480
rect 14536 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14856 11456
rect 14536 10368 14856 11392
rect 14536 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14856 10368
rect 14536 9280 14856 10304
rect 14536 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14856 9280
rect 14536 8192 14856 9216
rect 14536 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14856 8192
rect 14536 7104 14856 8128
rect 14536 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14856 7104
rect 14536 6016 14856 7040
rect 14536 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14856 6016
rect 14536 4928 14856 5952
rect 14536 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14856 4928
rect 14536 3840 14856 4864
rect 14536 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14856 3840
rect 14536 2752 14856 3776
rect 14536 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14856 2752
rect 14536 1664 14856 2688
rect 14536 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14856 1664
rect 14536 576 14856 1600
rect 14536 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14856 576
rect 14536 496 14856 512
rect 16894 18528 17214 19088
rect 16894 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17214 18528
rect 16894 17440 17214 18464
rect 16894 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17214 17440
rect 16894 16352 17214 17376
rect 16894 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17214 16352
rect 16894 15264 17214 16288
rect 16894 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17214 15264
rect 16894 14176 17214 15200
rect 16894 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17214 14176
rect 16894 13088 17214 14112
rect 16894 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17214 13088
rect 16894 12000 17214 13024
rect 16894 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17214 12000
rect 16894 10912 17214 11936
rect 16894 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17214 10912
rect 16894 9824 17214 10848
rect 16894 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17214 9824
rect 16894 8736 17214 9760
rect 16894 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17214 8736
rect 16894 7648 17214 8672
rect 16894 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17214 7648
rect 16894 6560 17214 7584
rect 16894 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17214 6560
rect 16894 5472 17214 6496
rect 16894 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17214 5472
rect 16894 4384 17214 5408
rect 16894 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17214 4384
rect 16894 3296 17214 4320
rect 16894 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17214 3296
rect 16894 2208 17214 3232
rect 16894 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17214 2208
rect 16894 1120 17214 2144
rect 16894 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17214 1120
rect 16894 496 17214 1056
rect 19251 19072 19571 19088
rect 19251 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19571 19072
rect 19251 17984 19571 19008
rect 19251 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19571 17984
rect 19251 16896 19571 17920
rect 19251 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19571 16896
rect 19251 15808 19571 16832
rect 19251 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19571 15808
rect 19251 14720 19571 15744
rect 19251 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19571 14720
rect 19251 13632 19571 14656
rect 19251 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19571 13632
rect 19251 12544 19571 13568
rect 19251 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19571 12544
rect 19251 11456 19571 12480
rect 19251 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19571 11456
rect 19251 10368 19571 11392
rect 19251 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19571 10368
rect 19251 9280 19571 10304
rect 19251 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19571 9280
rect 19251 8192 19571 9216
rect 19251 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19571 8192
rect 19251 7104 19571 8128
rect 19251 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19571 7104
rect 19251 6016 19571 7040
rect 19251 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19571 6016
rect 19251 4928 19571 5952
rect 19251 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19571 4928
rect 19251 3840 19571 4864
rect 19251 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19571 3840
rect 19251 2752 19571 3776
rect 19251 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19571 2752
rect 19251 1664 19571 2688
rect 19251 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19571 1664
rect 19251 576 19571 1600
rect 19251 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19571 576
rect 19251 496 19571 512
use sky130_fd_sc_hd__buf_2  _102_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1701704242
transform 1 0 13892 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1701704242
transform 1 0 13156 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1701704242
transform 1 0 14260 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _106_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 14168 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _107_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 11224 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_1  _108_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 11960 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _109_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10396 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _110_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15916 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _111_
timestamp 1701704242
transform -1 0 12512 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _112_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11960 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _113_
timestamp 1701704242
transform 1 0 13432 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _114_
timestamp 1701704242
transform -1 0 13432 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__and4b_4  _115_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 12144 0 1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__a22o_1  _116_
timestamp 1701704242
transform 1 0 13708 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _117_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12144 0 -1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_2  _118_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10120 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _119_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14076 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _120_
timestamp 1701704242
transform 1 0 14168 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_2  _121_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_2  _122_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 9292 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _123_
timestamp 1701704242
transform 1 0 8832 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _124_
timestamp 1701704242
transform 1 0 11040 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__nor4b_2  _125_
timestamp 1701704242
transform 1 0 9752 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _126_
timestamp 1701704242
transform 1 0 7452 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_4  _127_
timestamp 1701704242
transform 1 0 9476 0 -1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__and4bb_4  _128_
timestamp 1701704242
transform 1 0 11316 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _129_
timestamp 1701704242
transform 1 0 9016 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _130_
timestamp 1701704242
transform 1 0 9292 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_4  _131_
timestamp 1701704242
transform 1 0 10948 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _132_
timestamp 1701704242
transform 1 0 8372 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _133_
timestamp 1701704242
transform 1 0 9016 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _134_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16008 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _135_
timestamp 1701704242
transform -1 0 10396 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _136_
timestamp 1701704242
transform 1 0 9568 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _137_
timestamp 1701704242
transform 1 0 9660 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _138_
timestamp 1701704242
transform -1 0 10120 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _139_
timestamp 1701704242
transform 1 0 9476 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _140_
timestamp 1701704242
transform 1 0 10212 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _141_
timestamp 1701704242
transform 1 0 9384 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _142_
timestamp 1701704242
transform -1 0 18768 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _143_
timestamp 1701704242
transform 1 0 10120 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _144_
timestamp 1701704242
transform 1 0 11408 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _145_
timestamp 1701704242
transform -1 0 12512 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _146_
timestamp 1701704242
transform -1 0 6440 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _147_
timestamp 1701704242
transform 1 0 11040 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _148_
timestamp 1701704242
transform -1 0 11500 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _149_
timestamp 1701704242
transform -1 0 16008 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _150_
timestamp 1701704242
transform 1 0 11960 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _151_
timestamp 1701704242
transform -1 0 16744 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _152_
timestamp 1701704242
transform 1 0 5060 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _153_
timestamp 1701704242
transform 1 0 10212 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _154_
timestamp 1701704242
transform 1 0 11500 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _155_
timestamp 1701704242
transform 1 0 13064 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _156_
timestamp 1701704242
transform -1 0 13432 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _157_
timestamp 1701704242
transform -1 0 18308 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _158_
timestamp 1701704242
transform 1 0 10948 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _159_
timestamp 1701704242
transform -1 0 10580 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _160_
timestamp 1701704242
transform 1 0 10396 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _161_
timestamp 1701704242
transform 1 0 10856 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _162_
timestamp 1701704242
transform 1 0 10212 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _163_
timestamp 1701704242
transform 1 0 9384 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _164_
timestamp 1701704242
transform 1 0 10764 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _165_
timestamp 1701704242
transform 1 0 10028 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _166_
timestamp 1701704242
transform 1 0 10580 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _167_
timestamp 1701704242
transform 1 0 11408 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _168_
timestamp 1701704242
transform 1 0 8464 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _169_
timestamp 1701704242
transform -1 0 16744 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _170_
timestamp 1701704242
transform 1 0 16652 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _171_
timestamp 1701704242
transform 1 0 14536 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _172_
timestamp 1701704242
transform 1 0 15548 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _173_
timestamp 1701704242
transform 1 0 6440 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _174_
timestamp 1701704242
transform 1 0 7544 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _175_
timestamp 1701704242
transform 1 0 8372 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _176_
timestamp 1701704242
transform 1 0 2576 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _177_
timestamp 1701704242
transform 1 0 7728 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _178_
timestamp 1701704242
transform -1 0 17388 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _179_
timestamp 1701704242
transform 1 0 11224 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _180_
timestamp 1701704242
transform 1 0 10948 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _181_
timestamp 1701704242
transform 1 0 13524 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _182_
timestamp 1701704242
transform 1 0 11224 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _183_
timestamp 1701704242
transform 1 0 11592 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _184_
timestamp 1701704242
transform 1 0 4508 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _185_
timestamp 1701704242
transform 1 0 9292 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _186_
timestamp 1701704242
transform 1 0 9016 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _187_
timestamp 1701704242
transform -1 0 12788 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _188_
timestamp 1701704242
transform -1 0 9844 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _189_
timestamp 1701704242
transform -1 0 13340 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _190_
timestamp 1701704242
transform 1 0 9108 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _191_
timestamp 1701704242
transform -1 0 14536 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _192_
timestamp 1701704242
transform 1 0 16100 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _193_
timestamp 1701704242
transform -1 0 15824 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _194_
timestamp 1701704242
transform -1 0 15640 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 1701704242
transform 1 0 5612 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _196_
timestamp 1701704242
transform 1 0 6164 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _197_
timestamp 1701704242
transform -1 0 16744 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _198_
timestamp 1701704242
transform 1 0 3220 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _199_
timestamp 1701704242
transform 1 0 6808 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _200_
timestamp 1701704242
transform -1 0 15732 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _201_
timestamp 1701704242
transform 1 0 8372 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _202_
timestamp 1701704242
transform 1 0 16008 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _203_
timestamp 1701704242
transform -1 0 16376 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _204_
timestamp 1701704242
transform 1 0 14720 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _205_
timestamp 1701704242
transform 1 0 16100 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _206_
timestamp 1701704242
transform 1 0 5796 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _207_
timestamp 1701704242
transform 1 0 6072 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _208_
timestamp 1701704242
transform 1 0 8372 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _209_
timestamp 1701704242
transform 1 0 2484 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _210_
timestamp 1701704242
transform 1 0 6440 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _211_
timestamp 1701704242
transform -1 0 17388 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__dfxtp_1  _212_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17204 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _213_
timestamp 1701704242
transform -1 0 18216 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _214_
timestamp 1701704242
transform -1 0 16008 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _215_
timestamp 1701704242
transform 1 0 15272 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _216_
timestamp 1701704242
transform -1 0 15916 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _217_
timestamp 1701704242
transform -1 0 14168 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _218_
timestamp 1701704242
transform -1 0 14812 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _219_
timestamp 1701704242
transform -1 0 13892 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _220_
timestamp 1701704242
transform 1 0 13616 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _221_
timestamp 1701704242
transform -1 0 12420 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _222_
timestamp 1701704242
transform 1 0 12972 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _223_
timestamp 1701704242
transform 1 0 13524 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _224_
timestamp 1701704242
transform 1 0 13616 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _225_
timestamp 1701704242
transform -1 0 12420 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _226_
timestamp 1701704242
transform -1 0 12420 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _227_
timestamp 1701704242
transform -1 0 11408 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _228_
timestamp 1701704242
transform -1 0 8280 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _229_
timestamp 1701704242
transform 1 0 8280 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _230_
timestamp 1701704242
transform -1 0 7636 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _231_
timestamp 1701704242
transform 1 0 4692 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _232_
timestamp 1701704242
transform -1 0 13340 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _233_
timestamp 1701704242
transform 1 0 8832 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _234_
timestamp 1701704242
transform 1 0 15180 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _235_
timestamp 1701704242
transform -1 0 15180 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _236_
timestamp 1701704242
transform 1 0 14536 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _237_
timestamp 1701704242
transform -1 0 15732 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _238_
timestamp 1701704242
transform 1 0 14536 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _239_
timestamp 1701704242
transform 1 0 14996 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _240_
timestamp 1701704242
transform -1 0 14996 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _241_
timestamp 1701704242
transform 1 0 8740 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _242_
timestamp 1701704242
transform 1 0 9016 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _243_
timestamp 1701704242
transform 1 0 8648 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _244_
timestamp 1701704242
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _245_
timestamp 1701704242
transform 1 0 7544 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _246_
timestamp 1701704242
transform 1 0 6992 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _247_
timestamp 1701704242
transform 1 0 6992 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _248_
timestamp 1701704242
transform 1 0 5612 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _249_
timestamp 1701704242
transform 1 0 8372 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _250_
timestamp 1701704242
transform 1 0 5060 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _251_
timestamp 1701704242
transform 1 0 8096 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _252_
timestamp 1701704242
transform 1 0 5520 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _253_
timestamp 1701704242
transform 1 0 6440 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _254_
timestamp 1701704242
transform 1 0 4140 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _255_
timestamp 1701704242
transform 1 0 3220 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _256_
timestamp 1701704242
transform 1 0 3496 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _257_
timestamp 1701704242
transform 1 0 2392 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _258_
timestamp 1701704242
transform 1 0 3220 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _259_
timestamp 1701704242
transform 1 0 1564 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _260_
timestamp 1701704242
transform 1 0 1196 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _261_
timestamp 1701704242
transform 1 0 2116 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _262_
timestamp 1701704242
transform 1 0 1104 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _263_
timestamp 1701704242
transform 1 0 1472 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _264_
timestamp 1701704242
transform 1 0 3680 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _265_
timestamp 1701704242
transform 1 0 3220 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _266_
timestamp 1701704242
transform 1 0 4232 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _267_
timestamp 1701704242
transform 1 0 3404 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _268_
timestamp 1701704242
transform 1 0 5336 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _269_
timestamp 1701704242
transform 1 0 5796 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _270_
timestamp 1701704242
transform 1 0 5888 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _271_
timestamp 1701704242
transform 1 0 6164 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _272_
timestamp 1701704242
transform 1 0 6624 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _273_
timestamp 1701704242
transform 1 0 7636 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _274_
timestamp 1701704242
transform 1 0 6716 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _275_
timestamp 1701704242
transform 1 0 7820 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _276_
timestamp 1701704242
transform 1 0 4968 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _277_
timestamp 1701704242
transform 1 0 5980 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _278_
timestamp 1701704242
transform 1 0 4140 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _279_
timestamp 1701704242
transform 1 0 3864 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _280_
timestamp 1701704242
transform 1 0 5152 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _281_
timestamp 1701704242
transform 1 0 3680 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _282_
timestamp 1701704242
transform 1 0 3036 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _283_
timestamp 1701704242
transform 1 0 3128 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _284_
timestamp 1701704242
transform 1 0 1012 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _285_
timestamp 1701704242
transform 1 0 1564 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _286_
timestamp 1701704242
transform 1 0 920 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _287_
timestamp 1701704242
transform 1 0 1012 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _288_
timestamp 1701704242
transform 1 0 1380 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _289_
timestamp 1701704242
transform 1 0 1196 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _290_
timestamp 1701704242
transform 1 0 1564 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _291_
timestamp 1701704242
transform 1 0 1656 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _292_
timestamp 1701704242
transform 1 0 1932 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _293_
timestamp 1701704242
transform 1 0 1656 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _294_
timestamp 1701704242
transform 1 0 1656 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _295_
timestamp 1701704242
transform 1 0 3588 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _296_
timestamp 1701704242
transform 1 0 3404 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _297_
timestamp 1701704242
transform 1 0 3864 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _298_
timestamp 1701704242
transform 1 0 5060 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _299_
timestamp 1701704242
transform 1 0 5336 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _300_
timestamp 1701704242
transform 1 0 6072 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _301_
timestamp 1701704242
transform 1 0 6532 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _302_
timestamp 1701704242
transform 1 0 6716 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _303_
timestamp 1701704242
transform 1 0 6900 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _304_
timestamp 1701704242
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _305_
timestamp 1701704242
transform 1 0 8372 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _306_
timestamp 1701704242
transform 1 0 9200 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _307_
timestamp 1701704242
transform 1 0 9016 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _308_
timestamp 1701704242
transform 1 0 13892 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _309_
timestamp 1701704242
transform 1 0 10948 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _310_
timestamp 1701704242
transform 1 0 12420 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _311_
timestamp 1701704242
transform 1 0 13432 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _312_
timestamp 1701704242
transform 1 0 12972 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _313_
timestamp 1701704242
transform 1 0 16468 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _314_
timestamp 1701704242
transform -1 0 12328 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _315_
timestamp 1701704242
transform 1 0 16744 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _316_
timestamp 1701704242
transform 1 0 15272 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _317_
timestamp 1701704242
transform 1 0 11592 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _318_
timestamp 1701704242
transform -1 0 14996 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _319_
timestamp 1701704242
transform 1 0 14536 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _320_
timestamp 1701704242
transform -1 0 9384 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _321_
timestamp 1701704242
transform 1 0 8740 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _322_
timestamp 1701704242
transform -1 0 18584 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _323_
timestamp 1701704242
transform -1 0 10856 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _324_
timestamp 1701704242
transform -1 0 19044 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _325_
timestamp 1701704242
transform -1 0 18216 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _326_
timestamp 1701704242
transform -1 0 19136 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _327_
timestamp 1701704242
transform -1 0 17848 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _328_
timestamp 1701704242
transform -1 0 18952 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _329_
timestamp 1701704242
transform 1 0 16652 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _330_
timestamp 1701704242
transform -1 0 19136 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _331_
timestamp 1701704242
transform 1 0 17112 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _332_
timestamp 1701704242
transform -1 0 19044 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _333_
timestamp 1701704242
transform -1 0 18952 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _334_
timestamp 1701704242
transform -1 0 18860 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _335_
timestamp 1701704242
transform -1 0 18584 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _336_
timestamp 1701704242
transform -1 0 17940 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _337_
timestamp 1701704242
transform -1 0 18584 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _338_
timestamp 1701704242
transform -1 0 18124 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _339_
timestamp 1701704242
transform -1 0 18584 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _356_
timestamp 1701704242
transform -1 0 17020 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1701704242
transform -1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1701704242
transform -1 0 17020 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 5060 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1701704242
transform 1 0 3680 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1701704242
transform -1 0 9384 0 1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1701704242
transform 1 0 7176 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1701704242
transform 1 0 3588 0 1 12512
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1701704242
transform -1 0 4232 0 -1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1701704242
transform 1 0 6440 0 -1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1701704242
transform -1 0 8740 0 -1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1701704242
transform -1 0 13432 0 1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1701704242
transform -1 0 15548 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1701704242
transform -1 0 17296 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1701704242
transform 1 0 16652 0 1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1701704242
transform -1 0 13432 0 -1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1701704242
transform -1 0 15272 0 1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1701704242
transform 1 0 17204 0 1 12512
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1701704242
transform 1 0 16468 0 -1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_6 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1104 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_12 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1656 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_16 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 2024 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_23
timestamp 1701704242
transform 1 0 2668 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 1701704242
transform 1 0 3956 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1701704242
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1701704242
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_69 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6900 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_74
timestamp 1701704242
transform 1 0 7360 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1701704242
transform 1 0 8096 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_97
timestamp 1701704242
transform 1 0 9476 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_105
timestamp 1701704242
transform 1 0 10212 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1701704242
transform 1 0 10764 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1701704242
transform 1 0 10948 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_125 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12052 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1701704242
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_153
timestamp 1701704242
transform 1 0 14628 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_161
timestamp 1701704242
transform 1 0 15364 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1701704242
transform 1 0 15824 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_175
timestamp 1701704242
transform 1 0 16652 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_187
timestamp 1701704242
transform 1 0 17756 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197
timestamp 1701704242
transform 1 0 18676 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_104
timestamp 1701704242
transform 1 0 10120 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_172
timestamp 1701704242
transform 1 0 16376 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_189
timestamp 1701704242
transform 1 0 17940 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_201
timestamp 1701704242
transform 1 0 19044 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1701704242
transform 1 0 828 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_68
timestamp 1701704242
transform 1 0 6808 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_108
timestamp 1701704242
transform 1 0 10488 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_112
timestamp 1701704242
transform 1 0 10856 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_135
timestamp 1701704242
transform 1 0 12972 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_150
timestamp 1701704242
transform 1 0 14352 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_192
timestamp 1701704242
transform 1 0 18216 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_197
timestamp 1701704242
transform 1 0 18676 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_17
timestamp 1701704242
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_22
timestamp 1701704242
transform 1 0 2576 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_30
timestamp 1701704242
transform 1 0 3312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_49
timestamp 1701704242
transform 1 0 5060 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_81
timestamp 1701704242
transform 1 0 8004 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_88
timestamp 1701704242
transform 1 0 8648 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_95
timestamp 1701704242
transform 1 0 9292 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1701704242
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_119
timestamp 1701704242
transform 1 0 11500 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_127
timestamp 1701704242
transform 1 0 12236 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1701704242
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_178
timestamp 1701704242
transform 1 0 16928 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_182
timestamp 1701704242
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_187
timestamp 1701704242
transform 1 0 17756 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_32
timestamp 1701704242
transform 1 0 3496 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_44
timestamp 1701704242
transform 1 0 4600 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_59
timestamp 1701704242
transform 1 0 5980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_67
timestamp 1701704242
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_71
timestamp 1701704242
transform 1 0 7084 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_75
timestamp 1701704242
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp 1701704242
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_91
timestamp 1701704242
transform 1 0 8924 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_103
timestamp 1701704242
transform 1 0 10028 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_111
timestamp 1701704242
transform 1 0 10764 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_128
timestamp 1701704242
transform 1 0 12328 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_132
timestamp 1701704242
transform 1 0 12696 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 1701704242
transform 1 0 13064 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1701704242
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_153
timestamp 1701704242
transform 1 0 14628 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_163
timestamp 1701704242
transform 1 0 15548 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_167
timestamp 1701704242
transform 1 0 15916 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_197
timestamp 1701704242
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_201
timestamp 1701704242
transform 1 0 19044 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_14
timestamp 1701704242
transform 1 0 1840 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_31
timestamp 1701704242
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_49
timestamp 1701704242
transform 1 0 5060 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1701704242
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_61
timestamp 1701704242
transform 1 0 6164 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_65
timestamp 1701704242
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_83
timestamp 1701704242
transform 1 0 8188 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_91
timestamp 1701704242
transform 1 0 8924 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 1701704242
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1701704242
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_125
timestamp 1701704242
transform 1 0 12052 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_133
timestamp 1701704242
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_151
timestamp 1701704242
transform 1 0 14444 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_157
timestamp 1701704242
transform 1 0 14996 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_184
timestamp 1701704242
transform 1 0 17480 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_201
timestamp 1701704242
transform 1 0 19044 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 1701704242
transform 1 0 2208 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1701704242
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_41
timestamp 1701704242
transform 1 0 4324 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_65
timestamp 1701704242
transform 1 0 6532 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_105
timestamp 1701704242
transform 1 0 10212 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_111
timestamp 1701704242
transform 1 0 10764 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_119
timestamp 1701704242
transform 1 0 11500 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_136
timestamp 1701704242
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_157
timestamp 1701704242
transform 1 0 14996 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_166
timestamp 1701704242
transform 1 0 15824 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_182
timestamp 1701704242
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1701704242
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_200
timestamp 1701704242
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 1701704242
transform 1 0 828 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_27
timestamp 1701704242
transform 1 0 3036 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_35
timestamp 1701704242
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_52
timestamp 1701704242
transform 1 0 5336 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_57
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_76
timestamp 1701704242
transform 1 0 7544 0 -1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_133
timestamp 1701704242
transform 1 0 12788 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_145
timestamp 1701704242
transform 1 0 13892 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_151
timestamp 1701704242
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_169
timestamp 1701704242
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_177
timestamp 1701704242
transform 1 0 16836 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_181
timestamp 1701704242
transform 1 0 17204 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_185
timestamp 1701704242
transform 1 0 17572 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_11
timestamp 1701704242
transform 1 0 1564 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_33
timestamp 1701704242
transform 1 0 3588 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_66
timestamp 1701704242
transform 1 0 6624 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_78
timestamp 1701704242
transform 1 0 7728 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_96
timestamp 1701704242
transform 1 0 9384 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_104
timestamp 1701704242
transform 1 0 10120 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_114
timestamp 1701704242
transform 1 0 11040 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_126
timestamp 1701704242
transform 1 0 12144 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_153
timestamp 1701704242
transform 1 0 14628 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_157
timestamp 1701704242
transform 1 0 14996 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_164
timestamp 1701704242
transform 1 0 15640 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1701704242
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_200
timestamp 1701704242
transform 1 0 18952 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_3
timestamp 1701704242
transform 1 0 828 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_7
timestamp 1701704242
transform 1 0 1196 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_17
timestamp 1701704242
transform 1 0 2116 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_47
timestamp 1701704242
transform 1 0 4876 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1701704242
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_64
timestamp 1701704242
transform 1 0 6440 0 -1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_100
timestamp 1701704242
transform 1 0 9752 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_125
timestamp 1701704242
transform 1 0 12052 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_130
timestamp 1701704242
transform 1 0 12512 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_134
timestamp 1701704242
transform 1 0 12880 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_151
timestamp 1701704242
transform 1 0 14444 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1701704242
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_196
timestamp 1701704242
transform 1 0 18584 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_9
timestamp 1701704242
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_20
timestamp 1701704242
transform 1 0 2392 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_24
timestamp 1701704242
transform 1 0 2760 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_34
timestamp 1701704242
transform 1 0 3680 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_52
timestamp 1701704242
transform 1 0 5336 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_62
timestamp 1701704242
transform 1 0 6256 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_85
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_89
timestamp 1701704242
transform 1 0 8740 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1701704242
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_109
timestamp 1701704242
transform 1 0 10580 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_130
timestamp 1701704242
transform 1 0 12512 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1701704242
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1701704242
transform 1 0 13524 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_176
timestamp 1701704242
transform 1 0 16744 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_180
timestamp 1701704242
transform 1 0 17112 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_184
timestamp 1701704242
transform 1 0 17480 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_200
timestamp 1701704242
transform 1 0 18952 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_7
timestamp 1701704242
transform 1 0 1196 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_25
timestamp 1701704242
transform 1 0 2852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_35
timestamp 1701704242
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1701704242
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_74
timestamp 1701704242
transform 1 0 7360 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_78
timestamp 1701704242
transform 1 0 7728 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_84
timestamp 1701704242
transform 1 0 8280 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_99
timestamp 1701704242
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_113
timestamp 1701704242
transform 1 0 10948 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_141
timestamp 1701704242
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_158
timestamp 1701704242
transform 1 0 15088 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1701704242
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_169
timestamp 1701704242
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_182
timestamp 1701704242
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_200
timestamp 1701704242
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_71
timestamp 1701704242
transform 1 0 7084 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1701704242
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1701704242
transform 1 0 8372 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_156
timestamp 1701704242
transform 1 0 14904 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_164
timestamp 1701704242
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 1701704242
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_197
timestamp 1701704242
transform 1 0 18676 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp 1701704242
transform 1 0 19044 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_21
timestamp 1701704242
transform 1 0 2484 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_25
timestamp 1701704242
transform 1 0 2852 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_29
timestamp 1701704242
transform 1 0 3220 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_38
timestamp 1701704242
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1701704242
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1701704242
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_69
timestamp 1701704242
transform 1 0 6900 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_86
timestamp 1701704242
transform 1 0 8464 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_93
timestamp 1701704242
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_152
timestamp 1701704242
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_175
timestamp 1701704242
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_182
timestamp 1701704242
transform 1 0 17296 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_16
timestamp 1701704242
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_21
timestamp 1701704242
transform 1 0 2484 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1701704242
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_41
timestamp 1701704242
transform 1 0 4324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_57
timestamp 1701704242
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_75
timestamp 1701704242
transform 1 0 7452 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1701704242
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_98
timestamp 1701704242
transform 1 0 9568 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_107
timestamp 1701704242
transform 1 0 10396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_157
timestamp 1701704242
transform 1 0 14996 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_165
timestamp 1701704242
transform 1 0 15732 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_200
timestamp 1701704242
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_3
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_7
timestamp 1701704242
transform 1 0 1196 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_66
timestamp 1701704242
transform 1 0 6624 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_74
timestamp 1701704242
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_99
timestamp 1701704242
transform 1 0 9660 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_147
timestamp 1701704242
transform 1 0 14076 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_169
timestamp 1701704242
transform 1 0 16100 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_201
timestamp 1701704242
transform 1 0 19044 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_21
timestamp 1701704242
transform 1 0 2484 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1701704242
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_41
timestamp 1701704242
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_56
timestamp 1701704242
transform 1 0 5704 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_60
timestamp 1701704242
transform 1 0 6072 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_64
timestamp 1701704242
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1701704242
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp 1701704242
transform 1 0 8372 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_91
timestamp 1701704242
transform 1 0 8924 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_108
timestamp 1701704242
transform 1 0 10488 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_121
timestamp 1701704242
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1701704242
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1701704242
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_150
timestamp 1701704242
transform 1 0 14352 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_167
timestamp 1701704242
transform 1 0 15916 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_175
timestamp 1701704242
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_200
timestamp 1701704242
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_23
timestamp 1701704242
transform 1 0 2668 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_35
timestamp 1701704242
transform 1 0 3772 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_47
timestamp 1701704242
transform 1 0 4876 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_66
timestamp 1701704242
transform 1 0 6624 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_83
timestamp 1701704242
transform 1 0 8188 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_101
timestamp 1701704242
transform 1 0 9844 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1701704242
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_133
timestamp 1701704242
transform 1 0 12788 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_155
timestamp 1701704242
transform 1 0 14812 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1701704242
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_183
timestamp 1701704242
transform 1 0 17388 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_200
timestamp 1701704242
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_15
timestamp 1701704242
transform 1 0 1932 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_45
timestamp 1701704242
transform 1 0 4692 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_56
timestamp 1701704242
transform 1 0 5704 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_60
timestamp 1701704242
transform 1 0 6072 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_70
timestamp 1701704242
transform 1 0 6992 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_76
timestamp 1701704242
transform 1 0 7544 0 1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1701704242
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_97
timestamp 1701704242
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_112
timestamp 1701704242
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_116
timestamp 1701704242
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_130
timestamp 1701704242
transform 1 0 12512 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1701704242
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_141
timestamp 1701704242
transform 1 0 13524 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_147
timestamp 1701704242
transform 1 0 14076 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_154
timestamp 1701704242
transform 1 0 14720 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1701704242
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_200
timestamp 1701704242
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_26
timestamp 1701704242
transform 1 0 2944 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_30
timestamp 1701704242
transform 1 0 3312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_57
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_93
timestamp 1701704242
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1701704242
transform 1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 1701704242
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_130
timestamp 1701704242
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_154
timestamp 1701704242
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1701704242
transform 1 0 15732 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_178
timestamp 1701704242
transform 1 0 16928 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_186
timestamp 1701704242
transform 1 0 17664 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_3
timestamp 1701704242
transform 1 0 828 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_24
timestamp 1701704242
transform 1 0 2760 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_29
timestamp 1701704242
transform 1 0 3220 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_33
timestamp 1701704242
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_62
timestamp 1701704242
transform 1 0 6256 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_74
timestamp 1701704242
transform 1 0 7360 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1701704242
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_92
timestamp 1701704242
transform 1 0 9016 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_105
timestamp 1701704242
transform 1 0 10212 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_111
timestamp 1701704242
transform 1 0 10764 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_135
timestamp 1701704242
transform 1 0 12972 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1701704242
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_147
timestamp 1701704242
transform 1 0 14076 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_188
timestamp 1701704242
transform 1 0 17848 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_200
timestamp 1701704242
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_3
timestamp 1701704242
transform 1 0 828 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_20
timestamp 1701704242
transform 1 0 2392 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_39
timestamp 1701704242
transform 1 0 4140 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_43
timestamp 1701704242
transform 1 0 4508 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1701704242
transform 1 0 5428 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_73
timestamp 1701704242
transform 1 0 7268 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_102
timestamp 1701704242
transform 1 0 9936 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_151
timestamp 1701704242
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1701704242
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_183
timestamp 1701704242
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_201
timestamp 1701704242
transform 1 0 19044 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1701704242
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_15
timestamp 1701704242
transform 1 0 1932 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 1701704242
transform 1 0 3220 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_50
timestamp 1701704242
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_74
timestamp 1701704242
transform 1 0 7360 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_92
timestamp 1701704242
transform 1 0 9016 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_103
timestamp 1701704242
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_107
timestamp 1701704242
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_115
timestamp 1701704242
transform 1 0 11132 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_127
timestamp 1701704242
transform 1 0 12236 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_133
timestamp 1701704242
transform 1 0 12788 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_150
timestamp 1701704242
transform 1 0 14352 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1701704242
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_200
timestamp 1701704242
transform 1 0 18952 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_3
timestamp 1701704242
transform 1 0 828 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_22
timestamp 1701704242
transform 1 0 2576 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_82
timestamp 1701704242
transform 1 0 8096 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_104
timestamp 1701704242
transform 1 0 10120 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_129
timestamp 1701704242
transform 1 0 12420 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_151
timestamp 1701704242
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_172
timestamp 1701704242
transform 1 0 16376 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_3
timestamp 1701704242
transform 1 0 828 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_9
timestamp 1701704242
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_29
timestamp 1701704242
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_50
timestamp 1701704242
transform 1 0 5152 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_54
timestamp 1701704242
transform 1 0 5520 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_71
timestamp 1701704242
transform 1 0 7084 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1701704242
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_94
timestamp 1701704242
transform 1 0 9200 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_106
timestamp 1701704242
transform 1 0 10304 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_118
timestamp 1701704242
transform 1 0 11408 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_130
timestamp 1701704242
transform 1 0 12512 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_134
timestamp 1701704242
transform 1 0 12880 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1701704242
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_147
timestamp 1701704242
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_167
timestamp 1701704242
transform 1 0 15916 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_171
timestamp 1701704242
transform 1 0 16284 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_175
timestamp 1701704242
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_200
timestamp 1701704242
transform 1 0 18952 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1701704242
transform 1 0 828 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_33
timestamp 1701704242
transform 1 0 3588 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_45
timestamp 1701704242
transform 1 0 4692 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1701704242
transform 1 0 5428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_105
timestamp 1701704242
transform 1 0 10212 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_140
timestamp 1701704242
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_158
timestamp 1701704242
transform 1 0 15088 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1701704242
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_176
timestamp 1701704242
transform 1 0 16744 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_182
timestamp 1701704242
transform 1 0 17296 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_3
timestamp 1701704242
transform 1 0 828 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1701704242
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_45
timestamp 1701704242
transform 1 0 4692 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1701704242
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_85
timestamp 1701704242
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_98
timestamp 1701704242
transform 1 0 9568 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_118
timestamp 1701704242
transform 1 0 11408 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_122
timestamp 1701704242
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_127
timestamp 1701704242
transform 1 0 12236 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1701704242
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_192
timestamp 1701704242
transform 1 0 18216 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_197
timestamp 1701704242
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_3
timestamp 1701704242
transform 1 0 828 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_7
timestamp 1701704242
transform 1 0 1196 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_26
timestamp 1701704242
transform 1 0 2944 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_48
timestamp 1701704242
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_57
timestamp 1701704242
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_68
timestamp 1701704242
transform 1 0 6808 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_78
timestamp 1701704242
transform 1 0 7728 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_90
timestamp 1701704242
transform 1 0 8832 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_102
timestamp 1701704242
transform 1 0 9936 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 1701704242
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_123
timestamp 1701704242
transform 1 0 11868 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_151
timestamp 1701704242
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1701704242
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_190
timestamp 1701704242
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_198
timestamp 1701704242
transform 1 0 18768 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_3
timestamp 1701704242
transform 1 0 828 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_24
timestamp 1701704242
transform 1 0 2760 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_32
timestamp 1701704242
transform 1 0 3496 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_44
timestamp 1701704242
transform 1 0 4600 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_50
timestamp 1701704242
transform 1 0 5152 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_63
timestamp 1701704242
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1701704242
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_101
timestamp 1701704242
transform 1 0 9844 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_118
timestamp 1701704242
transform 1 0 11408 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_122
timestamp 1701704242
transform 1 0 11776 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_134
timestamp 1701704242
transform 1 0 12880 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_141
timestamp 1701704242
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1701704242
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_177
timestamp 1701704242
transform 1 0 16836 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_183
timestamp 1701704242
transform 1 0 17388 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1701704242
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_201
timestamp 1701704242
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_3
timestamp 1701704242
transform 1 0 828 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_31
timestamp 1701704242
transform 1 0 3404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_35
timestamp 1701704242
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_49
timestamp 1701704242
transform 1 0 5060 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_70
timestamp 1701704242
transform 1 0 6992 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_98
timestamp 1701704242
transform 1 0 9568 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_110
timestamp 1701704242
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1701704242
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_137
timestamp 1701704242
transform 1 0 13156 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_148
timestamp 1701704242
transform 1 0 14168 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1701704242
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_169
timestamp 1701704242
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_173
timestamp 1701704242
transform 1 0 16468 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_6
timestamp 1701704242
transform 1 0 1104 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1701704242
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3220 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_42
timestamp 1701704242
transform 1 0 4416 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_49
timestamp 1701704242
transform 1 0 5060 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_53
timestamp 1701704242
transform 1 0 5428 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_70
timestamp 1701704242
transform 1 0 6992 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1701704242
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_88
timestamp 1701704242
transform 1 0 8648 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_100
timestamp 1701704242
transform 1 0 9752 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_108
timestamp 1701704242
transform 1 0 10488 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_112
timestamp 1701704242
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_126
timestamp 1701704242
transform 1 0 12144 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_134
timestamp 1701704242
transform 1 0 12880 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_144
timestamp 1701704242
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_164
timestamp 1701704242
transform 1 0 15640 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_172
timestamp 1701704242
transform 1 0 16376 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1701704242
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_200
timestamp 1701704242
transform 1 0 18952 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_3
timestamp 1701704242
transform 1 0 828 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_11
timestamp 1701704242
transform 1 0 1564 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1701704242
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_57
timestamp 1701704242
transform 1 0 5796 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_107
timestamp 1701704242
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_142
timestamp 1701704242
transform 1 0 13616 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_176
timestamp 1701704242
transform 1 0 16744 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_199
timestamp 1701704242
transform 1 0 18860 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_6
timestamp 1701704242
transform 1 0 1104 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_18
timestamp 1701704242
transform 1 0 2208 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_24
timestamp 1701704242
transform 1 0 2760 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1701704242
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1701704242
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_85
timestamp 1701704242
transform 1 0 8372 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_89
timestamp 1701704242
transform 1 0 8740 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_109
timestamp 1701704242
transform 1 0 10580 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_116
timestamp 1701704242
transform 1 0 11224 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1701704242
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1701704242
transform 1 0 13524 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_191
timestamp 1701704242
transform 1 0 18124 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1701704242
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_197
timestamp 1701704242
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_12
timestamp 1701704242
transform 1 0 1656 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_24
timestamp 1701704242
transform 1 0 2760 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1701704242
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1701704242
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1701704242
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1701704242
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1701704242
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1701704242
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_85
timestamp 1701704242
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1701704242
transform 1 0 9476 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1701704242
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_113
timestamp 1701704242
transform 1 0 10948 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_117
timestamp 1701704242
transform 1 0 11316 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_121
timestamp 1701704242
transform 1 0 11684 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_128
timestamp 1701704242
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_139
timestamp 1701704242
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_153
timestamp 1701704242
transform 1 0 14628 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1701704242
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1701704242
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1701704242
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_197
timestamp 1701704242
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 19136 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input2 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12972 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1701704242
transform 1 0 10396 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1701704242
transform 1 0 12604 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1701704242
transform 1 0 11684 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  max_cap1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12512 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  max_cap6
timestamp 1701704242
transform -1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap7
timestamp 1701704242
transform -1 0 11316 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  max_cap9 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 9200 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap10
timestamp 1701704242
transform -1 0 13892 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap11
timestamp 1701704242
transform 1 0 14168 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 19412 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 19412 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 19412 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 19412 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 19412 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 19412 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 19412 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 19412 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 19412 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 19412 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 19412 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 19412 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 19412 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 19412 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 19412 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 19412 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1701704242
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1701704242
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 19412 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1701704242
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 19412 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1701704242
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 19412 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1701704242
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 19412 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1701704242
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1701704242
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 19412 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1701704242
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1701704242
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 19412 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1701704242
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 19412 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1701704242
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1701704242
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1701704242
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1701704242
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1701704242
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1701704242
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1701704242
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_77
timestamp 1701704242
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp 1701704242
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp 1701704242
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp 1701704242
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_85
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_86
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp 1701704242
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp 1701704242
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_89
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_90
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_91
timestamp 1701704242
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_92
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_93
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_94
timestamp 1701704242
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_95
timestamp 1701704242
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_96
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_97
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_98
timestamp 1701704242
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp 1701704242
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp 1701704242
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_103
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp 1701704242
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_108
timestamp 1701704242
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_109
timestamp 1701704242
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp 1701704242
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_113
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_114
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_115
timestamp 1701704242
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_116
timestamp 1701704242
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_117
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_118
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_119
timestamp 1701704242
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_120
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_121
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_122
timestamp 1701704242
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_123
timestamp 1701704242
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_124
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_125
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_126
timestamp 1701704242
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_127
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_128
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_129
timestamp 1701704242
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_130
timestamp 1701704242
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_131
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_132
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_133
timestamp 1701704242
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_134
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_135
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_136
timestamp 1701704242
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_137
timestamp 1701704242
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_138
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_139
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_140
timestamp 1701704242
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_141
timestamp 1701704242
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_142
timestamp 1701704242
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_143
timestamp 1701704242
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_144
timestamp 1701704242
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_145
timestamp 1701704242
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_146
timestamp 1701704242
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_147
timestamp 1701704242
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_148
timestamp 1701704242
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_149
timestamp 1701704242
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_150
timestamp 1701704242
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_151
timestamp 1701704242
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_152
timestamp 1701704242
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_153
timestamp 1701704242
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_154
timestamp 1701704242
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_155
timestamp 1701704242
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_156
timestamp 1701704242
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_157
timestamp 1701704242
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_158
timestamp 1701704242
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_159
timestamp 1701704242
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_160
timestamp 1701704242
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_161
timestamp 1701704242
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_162
timestamp 1701704242
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_163
timestamp 1701704242
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_164
timestamp 1701704242
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_165
timestamp 1701704242
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_166
timestamp 1701704242
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_167
timestamp 1701704242
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_168
timestamp 1701704242
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_169
timestamp 1701704242
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_170
timestamp 1701704242
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_171
timestamp 1701704242
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_172
timestamp 1701704242
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_173
timestamp 1701704242
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_174
timestamp 1701704242
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_175
timestamp 1701704242
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_176
timestamp 1701704242
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_177
timestamp 1701704242
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_178
timestamp 1701704242
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_179
timestamp 1701704242
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_180
timestamp 1701704242
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_181
timestamp 1701704242
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_182
timestamp 1701704242
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_183
timestamp 1701704242
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_184
timestamp 1701704242
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_185
timestamp 1701704242
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_186
timestamp 1701704242
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_187
timestamp 1701704242
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_188
timestamp 1701704242
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_189
timestamp 1701704242
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_190
timestamp 1701704242
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_191
timestamp 1701704242
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_192
timestamp 1701704242
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_193
timestamp 1701704242
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  tdc0.g_dly_chain_even\[0\].dly_stg pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 19136 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  tdc0.g_dly_chain_even\[1\].dly_stg pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14628 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[2\].dly_stg pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17572 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[3\].dly_stg
timestamp 1701704242
transform 1 0 15640 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[4\].dly_stg
timestamp 1701704242
transform -1 0 15732 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[5\].dly_stg
timestamp 1701704242
transform 1 0 15548 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[6\].dly_stg
timestamp 1701704242
transform 1 0 14168 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[7\].dly_stg
timestamp 1701704242
transform -1 0 14444 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[8\].dly_stg
timestamp 1701704242
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[9\].dly_stg
timestamp 1701704242
transform -1 0 13800 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[10\].dly_stg
timestamp 1701704242
transform 1 0 13800 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[11\].dly_stg
timestamp 1701704242
transform -1 0 13064 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[12\].dly_stg
timestamp 1701704242
transform -1 0 13248 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[13\].dly_stg
timestamp 1701704242
transform -1 0 12972 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[14\].dly_stg
timestamp 1701704242
transform -1 0 12788 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[15\].dly_stg
timestamp 1701704242
transform 1 0 11500 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[16\].dly_stg
timestamp 1701704242
transform 1 0 11500 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[17\].dly_stg
timestamp 1701704242
transform 1 0 11592 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[18\].dly_stg
timestamp 1701704242
transform 1 0 10948 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[19\].dly_stg
timestamp 1701704242
transform -1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[20\].dly_stg
timestamp 1701704242
transform 1 0 11408 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[21\].dly_stg
timestamp 1701704242
transform 1 0 12972 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[22\].dly_stg
timestamp 1701704242
transform -1 0 13800 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[23\].dly_stg
timestamp 1701704242
transform -1 0 13800 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[24\].dly_stg
timestamp 1701704242
transform -1 0 13432 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[25\].dly_stg
timestamp 1701704242
transform -1 0 15364 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[26\].dly_stg
timestamp 1701704242
transform -1 0 14260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[27\].dly_stg
timestamp 1701704242
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[28\].dly_stg
timestamp 1701704242
transform 1 0 13984 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[29\].dly_stg
timestamp 1701704242
transform 1 0 13064 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[30\].dly_stg
timestamp 1701704242
transform 1 0 9660 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[31\].dly_stg
timestamp 1701704242
transform -1 0 10856 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[32\].dly_stg
timestamp 1701704242
transform -1 0 8740 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[33\].dly_stg
timestamp 1701704242
transform -1 0 8188 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[34\].dly_stg
timestamp 1701704242
transform -1 0 8188 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[35\].dly_stg
timestamp 1701704242
transform 1 0 6348 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[36\].dly_stg
timestamp 1701704242
transform -1 0 7084 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[37\].dly_stg
timestamp 1701704242
transform -1 0 6532 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[38\].dly_stg
timestamp 1701704242
transform -1 0 6256 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[39\].dly_stg
timestamp 1701704242
transform -1 0 5796 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[40\].dly_stg
timestamp 1701704242
transform -1 0 6072 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[41\].dly_stg
timestamp 1701704242
transform -1 0 5060 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[42\].dly_stg
timestamp 1701704242
transform -1 0 4232 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[43\].dly_stg
timestamp 1701704242
transform -1 0 4140 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[44\].dly_stg
timestamp 1701704242
transform -1 0 2576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[45\].dly_stg
timestamp 1701704242
transform -1 0 3128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[46\].dly_stg
timestamp 1701704242
transform -1 0 1564 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[47\].dly_stg
timestamp 1701704242
transform -1 0 2760 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[48\].dly_stg
timestamp 1701704242
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[49\].dly_stg
timestamp 1701704242
transform -1 0 1564 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[50\].dly_stg
timestamp 1701704242
transform -1 0 2116 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[51\].dly_stg
timestamp 1701704242
transform 1 0 1564 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[52\].dly_stg
timestamp 1701704242
transform 1 0 1748 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[53\].dly_stg
timestamp 1701704242
transform -1 0 2944 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[54\].dly_stg
timestamp 1701704242
transform 1 0 2576 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[55\].dly_stg
timestamp 1701704242
transform -1 0 3128 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[56\].dly_stg
timestamp 1701704242
transform -1 0 4048 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[57\].dly_stg
timestamp 1701704242
transform -1 0 5152 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[58\].dly_stg
timestamp 1701704242
transform 1 0 4600 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[59\].dly_stg
timestamp 1701704242
transform -1 0 5704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[60\].dly_stg
timestamp 1701704242
transform -1 0 5704 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[61\].dly_stg
timestamp 1701704242
transform -1 0 6624 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[62\].dly_stg
timestamp 1701704242
transform -1 0 6072 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[63\].dly_stg
timestamp 1701704242
transform -1 0 5060 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[64\].dly_stg
timestamp 1701704242
transform -1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[65\].dly_stg
timestamp 1701704242
transform -1 0 4968 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[66\].dly_stg
timestamp 1701704242
transform -1 0 5244 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[67\].dly_stg
timestamp 1701704242
transform -1 0 4968 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[68\].dly_stg
timestamp 1701704242
transform -1 0 3772 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[69\].dly_stg
timestamp 1701704242
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[70\].dly_stg
timestamp 1701704242
transform -1 0 3128 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[71\].dly_stg
timestamp 1701704242
transform -1 0 2300 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[72\].dly_stg
timestamp 1701704242
transform -1 0 1748 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[73\].dly_stg
timestamp 1701704242
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[74\].dly_stg
timestamp 1701704242
transform -1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[75\].dly_stg
timestamp 1701704242
transform -1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[76\].dly_stg
timestamp 1701704242
transform -1 0 1196 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[77\].dly_stg
timestamp 1701704242
transform 1 0 1288 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[78\].dly_stg
timestamp 1701704242
transform -1 0 1564 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[79\].dly_stg
timestamp 1701704242
transform 1 0 1656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[80\].dly_stg
timestamp 1701704242
transform 1 0 1932 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[81\].dly_stg
timestamp 1701704242
transform -1 0 1288 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[82\].dly_stg
timestamp 1701704242
transform -1 0 1564 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[83\].dly_stg
timestamp 1701704242
transform -1 0 2392 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[84\].dly_stg
timestamp 1701704242
transform 1 0 2760 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[85\].dly_stg
timestamp 1701704242
transform -1 0 2576 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[86\].dly_stg
timestamp 1701704242
transform -1 0 4232 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[87\].dly_stg
timestamp 1701704242
transform 1 0 3588 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[88\].dly_stg
timestamp 1701704242
transform -1 0 5152 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[89\].dly_stg
timestamp 1701704242
transform -1 0 5704 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[90\].dly_stg
timestamp 1701704242
transform 1 0 5980 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[91\].dly_stg
timestamp 1701704242
transform -1 0 7084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[92\].dly_stg
timestamp 1701704242
transform -1 0 7176 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[93\].dly_stg
timestamp 1701704242
transform -1 0 8372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[94\].dly_stg
timestamp 1701704242
transform -1 0 8280 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[95\].dly_stg
timestamp 1701704242
transform -1 0 10120 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[96\].dly_stg
timestamp 1701704242
transform -1 0 10580 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[97\].dly_stg
timestamp 1701704242
transform -1 0 11500 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[98\].dly_stg
timestamp 1701704242
transform -1 0 12328 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[99\].dly_stg
timestamp 1701704242
transform 1 0 12880 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[100\].dly_stg
timestamp 1701704242
transform -1 0 14352 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[101\].dly_stg
timestamp 1701704242
transform 1 0 13800 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[102\].dly_stg
timestamp 1701704242
transform -1 0 15456 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[103\].dly_stg
timestamp 1701704242
transform 1 0 14720 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[104\].dly_stg
timestamp 1701704242
transform -1 0 16560 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[105\].dly_stg
timestamp 1701704242
transform 1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[106\].dly_stg
timestamp 1701704242
transform 1 0 14720 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[107\].dly_stg
timestamp 1701704242
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[108\].dly_stg
timestamp 1701704242
transform 1 0 15640 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[109\].dly_stg
timestamp 1701704242
transform -1 0 16284 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[110\].dly_stg
timestamp 1701704242
transform 1 0 16192 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[111\].dly_stg
timestamp 1701704242
transform 1 0 17020 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[112\].dly_stg
timestamp 1701704242
transform -1 0 17296 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[113\].dly_stg
timestamp 1701704242
transform 1 0 18676 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[114\].dly_stg
timestamp 1701704242
transform 1 0 18216 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[115\].dly_stg
timestamp 1701704242
transform -1 0 18308 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[116\].dly_stg
timestamp 1701704242
transform 1 0 17204 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[117\].dly_stg
timestamp 1701704242
transform -1 0 18308 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[118\].dly_stg
timestamp 1701704242
transform 1 0 18676 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[119\].dly_stg
timestamp 1701704242
transform -1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[120\].dly_stg
timestamp 1701704242
transform 1 0 18676 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[121\].dly_stg
timestamp 1701704242
transform 1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[122\].dly_stg
timestamp 1701704242
transform 1 0 18860 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[123\].dly_stg
timestamp 1701704242
transform -1 0 18492 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[124\].dly_stg
timestamp 1701704242
transform 1 0 18308 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[125\].dly_stg
timestamp 1701704242
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[126\].dly_stg
timestamp 1701704242
transform -1 0 16836 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[127\].dly_stg
timestamp 1701704242
transform 1 0 17020 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_even\[128\].dly_stg
timestamp 1701704242
transform -1 0 17112 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[0\].dly_stg
timestamp 1701704242
transform -1 0 17848 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[1\].dly_stg
timestamp 1701704242
transform -1 0 16652 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[2\].dly_stg
timestamp 1701704242
transform -1 0 16376 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[3\].dly_stg
timestamp 1701704242
transform -1 0 15640 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[4\].dly_stg
timestamp 1701704242
transform -1 0 15180 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[5\].dly_stg
timestamp 1701704242
transform -1 0 14720 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[6\].dly_stg
timestamp 1701704242
transform 1 0 13524 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[7\].dly_stg
timestamp 1701704242
transform 1 0 13800 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[8\].dly_stg
timestamp 1701704242
transform -1 0 12972 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[9\].dly_stg
timestamp 1701704242
transform -1 0 14904 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[10\].dly_stg
timestamp 1701704242
transform 1 0 12880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[11\].dly_stg
timestamp 1701704242
transform -1 0 14444 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[12\].dly_stg
timestamp 1701704242
transform -1 0 12880 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[13\].dly_stg
timestamp 1701704242
transform -1 0 12696 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[14\].dly_stg
timestamp 1701704242
transform -1 0 11224 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[15\].dly_stg
timestamp 1701704242
transform -1 0 11224 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[16\].dly_stg
timestamp 1701704242
transform -1 0 10856 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[17\].dly_stg
timestamp 1701704242
transform -1 0 8648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[18\].dly_stg
timestamp 1701704242
transform -1 0 9752 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[19\].dly_stg
timestamp 1701704242
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[20\].dly_stg
timestamp 1701704242
transform 1 0 10304 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[21\].dly_stg
timestamp 1701704242
transform 1 0 13064 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[22\].dly_stg
timestamp 1701704242
transform 1 0 13800 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[23\].dly_stg
timestamp 1701704242
transform 1 0 15364 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[24\].dly_stg
timestamp 1701704242
transform 1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[25\].dly_stg
timestamp 1701704242
transform 1 0 15640 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[26\].dly_stg
timestamp 1701704242
transform -1 0 15088 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[27\].dly_stg
timestamp 1701704242
transform -1 0 14536 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[28\].dly_stg
timestamp 1701704242
transform -1 0 14168 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[29\].dly_stg
timestamp 1701704242
transform -1 0 11776 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[30\].dly_stg
timestamp 1701704242
transform -1 0 9292 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[31\].dly_stg
timestamp 1701704242
transform -1 0 9200 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[32\].dly_stg
timestamp 1701704242
transform -1 0 8648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[33\].dly_stg
timestamp 1701704242
transform -1 0 7728 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[34\].dly_stg
timestamp 1701704242
transform -1 0 7912 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[35\].dly_stg
timestamp 1701704242
transform -1 0 6348 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[36\].dly_stg
timestamp 1701704242
transform -1 0 7728 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[37\].dly_stg
timestamp 1701704242
transform -1 0 6072 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[38\].dly_stg
timestamp 1701704242
transform -1 0 8188 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[39\].dly_stg
timestamp 1701704242
transform -1 0 5520 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[40\].dly_stg
timestamp 1701704242
transform -1 0 6992 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[41\].dly_stg
timestamp 1701704242
transform -1 0 4784 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[42\].dly_stg
timestamp 1701704242
transform -1 0 4140 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[43\].dly_stg
timestamp 1701704242
transform -1 0 3864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[44\].dly_stg
timestamp 1701704242
transform -1 0 3128 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[45\].dly_stg
timestamp 1701704242
transform 1 0 3220 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[46\].dly_stg
timestamp 1701704242
transform -1 0 2116 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[47\].dly_stg
timestamp 1701704242
transform -1 0 2944 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[48\].dly_stg
timestamp 1701704242
transform 1 0 1932 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[49\].dly_stg
timestamp 1701704242
transform -1 0 1840 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[50\].dly_stg
timestamp 1701704242
transform -1 0 1564 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[51\].dly_stg
timestamp 1701704242
transform 1 0 2024 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[52\].dly_stg
timestamp 1701704242
transform 1 0 2484 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[53\].dly_stg
timestamp 1701704242
transform -1 0 3220 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[54\].dly_stg
timestamp 1701704242
transform 1 0 3312 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[55\].dly_stg
timestamp 1701704242
transform 1 0 4600 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[56\].dly_stg
timestamp 1701704242
transform 1 0 4048 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[57\].dly_stg
timestamp 1701704242
transform 1 0 5152 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[58\].dly_stg
timestamp 1701704242
transform -1 0 5980 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[59\].dly_stg
timestamp 1701704242
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[60\].dly_stg
timestamp 1701704242
transform 1 0 5888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[61\].dly_stg
timestamp 1701704242
transform 1 0 6164 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[62\].dly_stg
timestamp 1701704242
transform 1 0 7268 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[63\].dly_stg
timestamp 1701704242
transform -1 0 5520 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[64\].dly_stg
timestamp 1701704242
transform -1 0 6624 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[65\].dly_stg
timestamp 1701704242
transform -1 0 5520 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[66\].dly_stg
timestamp 1701704242
transform -1 0 4416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[67\].dly_stg
timestamp 1701704242
transform -1 0 5336 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[68\].dly_stg
timestamp 1701704242
transform 1 0 4600 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[69\].dly_stg
timestamp 1701704242
transform -1 0 2852 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[70\].dly_stg
timestamp 1701704242
transform -1 0 3128 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[71\].dly_stg
timestamp 1701704242
transform -1 0 2484 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[72\].dly_stg
timestamp 1701704242
transform -1 0 2484 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[73\].dly_stg
timestamp 1701704242
transform -1 0 1472 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[74\].dly_stg
timestamp 1701704242
transform -1 0 1748 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[75\].dly_stg
timestamp 1701704242
transform 1 0 2116 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[76\].dly_stg
timestamp 1701704242
transform 1 0 1288 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[77\].dly_stg
timestamp 1701704242
transform -1 0 1288 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[78\].dly_stg
timestamp 1701704242
transform 1 0 1840 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[79\].dly_stg
timestamp 1701704242
transform -1 0 1840 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[80\].dly_stg
timestamp 1701704242
transform -1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[81\].dly_stg
timestamp 1701704242
transform -1 0 1196 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[82\].dly_stg
timestamp 1701704242
transform 1 0 2300 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[83\].dly_stg
timestamp 1701704242
transform 1 0 3128 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[84\].dly_stg
timestamp 1701704242
transform 1 0 2852 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[85\].dly_stg
timestamp 1701704242
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[86\].dly_stg
timestamp 1701704242
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[87\].dly_stg
timestamp 1701704242
transform 1 0 5336 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[88\].dly_stg
timestamp 1701704242
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[89\].dly_stg
timestamp 1701704242
transform 1 0 6256 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[90\].dly_stg
timestamp 1701704242
transform 1 0 6348 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[91\].dly_stg
timestamp 1701704242
transform 1 0 7176 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[92\].dly_stg
timestamp 1701704242
transform 1 0 7176 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[93\].dly_stg
timestamp 1701704242
transform 1 0 8648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[94\].dly_stg
timestamp 1701704242
transform 1 0 8740 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[95\].dly_stg
timestamp 1701704242
transform 1 0 10948 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[96\].dly_stg
timestamp 1701704242
transform 1 0 11224 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[97\].dly_stg
timestamp 1701704242
transform 1 0 12420 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[98\].dly_stg
timestamp 1701704242
transform 1 0 12604 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[99\].dly_stg
timestamp 1701704242
transform 1 0 12788 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[100\].dly_stg
timestamp 1701704242
transform 1 0 14352 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[101\].dly_stg
timestamp 1701704242
transform -1 0 13432 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[102\].dly_stg
timestamp 1701704242
transform -1 0 16652 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[103\].dly_stg
timestamp 1701704242
transform 1 0 15640 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[104\].dly_stg
timestamp 1701704242
transform -1 0 15824 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[105\].dly_stg
timestamp 1701704242
transform -1 0 15640 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[106\].dly_stg
timestamp 1701704242
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[107\].dly_stg
timestamp 1701704242
transform 1 0 14720 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[108\].dly_stg
timestamp 1701704242
transform -1 0 15548 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[109\].dly_stg
timestamp 1701704242
transform 1 0 16560 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[110\].dly_stg
timestamp 1701704242
transform 1 0 10488 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[111\].dly_stg
timestamp 1701704242
transform -1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[112\].dly_stg
timestamp 1701704242
transform 1 0 16928 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[113\].dly_stg
timestamp 1701704242
transform -1 0 18492 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[114\].dly_stg
timestamp 1701704242
transform -1 0 17480 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[115\].dly_stg
timestamp 1701704242
transform 1 0 18676 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[116\].dly_stg
timestamp 1701704242
transform -1 0 17296 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[117\].dly_stg
timestamp 1701704242
transform -1 0 18400 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[118\].dly_stg
timestamp 1701704242
transform -1 0 17112 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[119\].dly_stg
timestamp 1701704242
transform -1 0 18952 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[120\].dly_stg
timestamp 1701704242
transform 1 0 18216 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[121\].dly_stg
timestamp 1701704242
transform -1 0 18952 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[122\].dly_stg
timestamp 1701704242
transform -1 0 17112 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[123\].dly_stg
timestamp 1701704242
transform -1 0 17756 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[124\].dly_stg
timestamp 1701704242
transform -1 0 18032 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[125\].dly_stg
timestamp 1701704242
transform -1 0 17112 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[126\].dly_stg
timestamp 1701704242
transform -1 0 17572 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave\[127\].dly_stg
timestamp 1701704242
transform 1 0 18584 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[0\].dly_stg
timestamp 1701704242
transform -1 0 16376 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[1\].dly_stg
timestamp 1701704242
transform -1 0 16652 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[2\].dly_stg
timestamp 1701704242
transform -1 0 17296 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[3\].dly_stg
timestamp 1701704242
transform -1 0 16100 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[4\].dly_stg
timestamp 1701704242
transform -1 0 15548 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[5\].dly_stg
timestamp 1701704242
transform -1 0 14996 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[6\].dly_stg
timestamp 1701704242
transform -1 0 14720 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[7\].dly_stg
timestamp 1701704242
transform -1 0 14076 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[8\].dly_stg
timestamp 1701704242
transform -1 0 14352 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[9\].dly_stg
timestamp 1701704242
transform -1 0 13616 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[10\].dly_stg
timestamp 1701704242
transform -1 0 13340 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[11\].dly_stg
timestamp 1701704242
transform 1 0 13800 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[12\].dly_stg
timestamp 1701704242
transform -1 0 13064 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[13\].dly_stg
timestamp 1701704242
transform -1 0 12236 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[14\].dly_stg
timestamp 1701704242
transform -1 0 12052 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[15\].dly_stg
timestamp 1701704242
transform -1 0 11592 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[16\].dly_stg
timestamp 1701704242
transform -1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[17\].dly_stg
timestamp 1701704242
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[18\].dly_stg
timestamp 1701704242
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[19\].dly_stg
timestamp 1701704242
transform 1 0 12696 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[20\].dly_stg
timestamp 1701704242
transform 1 0 12512 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[21\].dly_stg
timestamp 1701704242
transform 1 0 13340 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[22\].dly_stg
timestamp 1701704242
transform 1 0 13984 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[23\].dly_stg
timestamp 1701704242
transform 1 0 13708 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[24\].dly_stg
timestamp 1701704242
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[25\].dly_stg
timestamp 1701704242
transform 1 0 15088 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[26\].dly_stg
timestamp 1701704242
transform -1 0 14168 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[27\].dly_stg
timestamp 1701704242
transform -1 0 13984 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[28\].dly_stg
timestamp 1701704242
transform -1 0 13892 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[29\].dly_stg
timestamp 1701704242
transform -1 0 12236 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[30\].dly_stg
timestamp 1701704242
transform -1 0 9568 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[31\].dly_stg
timestamp 1701704242
transform -1 0 9016 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[32\].dly_stg
timestamp 1701704242
transform -1 0 7176 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[33\].dly_stg
timestamp 1701704242
transform -1 0 7636 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[34\].dly_stg
timestamp 1701704242
transform -1 0 7912 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[35\].dly_stg
timestamp 1701704242
transform -1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[36\].dly_stg
timestamp 1701704242
transform -1 0 7452 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[37\].dly_stg
timestamp 1701704242
transform -1 0 5704 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[38\].dly_stg
timestamp 1701704242
transform -1 0 6348 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[39\].dly_stg
timestamp 1701704242
transform -1 0 5428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[40\].dly_stg
timestamp 1701704242
transform -1 0 4784 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[41\].dly_stg
timestamp 1701704242
transform -1 0 4416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[42\].dly_stg
timestamp 1701704242
transform -1 0 3588 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[43\].dly_stg
timestamp 1701704242
transform -1 0 2852 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[44\].dly_stg
timestamp 1701704242
transform -1 0 2392 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[45\].dly_stg
timestamp 1701704242
transform -1 0 1748 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[46\].dly_stg
timestamp 1701704242
transform -1 0 2024 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[47\].dly_stg
timestamp 1701704242
transform -1 0 2484 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[48\].dly_stg
timestamp 1701704242
transform 1 0 2392 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[49\].dly_stg
timestamp 1701704242
transform 1 0 2668 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[50\].dly_stg
timestamp 1701704242
transform -1 0 2116 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[51\].dly_stg
timestamp 1701704242
transform -1 0 2852 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[52\].dly_stg
timestamp 1701704242
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[53\].dly_stg
timestamp 1701704242
transform 1 0 4876 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[54\].dly_stg
timestamp 1701704242
transform 1 0 3312 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[55\].dly_stg
timestamp 1701704242
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[56\].dly_stg
timestamp 1701704242
transform 1 0 4600 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[57\].dly_stg
timestamp 1701704242
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[58\].dly_stg
timestamp 1701704242
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[59\].dly_stg
timestamp 1701704242
transform 1 0 5428 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[60\].dly_stg
timestamp 1701704242
transform 1 0 5428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[61\].dly_stg
timestamp 1701704242
transform -1 0 5704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[62\].dly_stg
timestamp 1701704242
transform 1 0 6072 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[63\].dly_stg
timestamp 1701704242
transform -1 0 5244 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[64\].dly_stg
timestamp 1701704242
transform -1 0 4968 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[65\].dly_stg
timestamp 1701704242
transform -1 0 4692 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[66\].dly_stg
timestamp 1701704242
transform -1 0 4140 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[67\].dly_stg
timestamp 1701704242
transform -1 0 3128 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[68\].dly_stg
timestamp 1701704242
transform -1 0 3496 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[69\].dly_stg
timestamp 1701704242
transform -1 0 3220 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[70\].dly_stg
timestamp 1701704242
transform -1 0 2852 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[71\].dly_stg
timestamp 1701704242
transform -1 0 1472 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[72\].dly_stg
timestamp 1701704242
transform -1 0 2024 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[73\].dly_stg
timestamp 1701704242
transform -1 0 1196 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[74\].dly_stg
timestamp 1701704242
transform -1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[75\].dly_stg
timestamp 1701704242
transform 1 0 1564 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[76\].dly_stg
timestamp 1701704242
transform -1 0 1840 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[77\].dly_stg
timestamp 1701704242
transform -1 0 1288 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[78\].dly_stg
timestamp 1701704242
transform -1 0 1288 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[79\].dly_stg
timestamp 1701704242
transform -1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[80\].dly_stg
timestamp 1701704242
transform 1 0 1196 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[81\].dly_stg
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[82\].dly_stg
timestamp 1701704242
transform 1 0 1472 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[83\].dly_stg
timestamp 1701704242
transform 1 0 2024 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[84\].dly_stg
timestamp 1701704242
transform 1 0 2576 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[85\].dly_stg
timestamp 1701704242
transform 1 0 4048 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[86\].dly_stg
timestamp 1701704242
transform 1 0 4508 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[87\].dly_stg
timestamp 1701704242
transform 1 0 5152 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[88\].dly_stg
timestamp 1701704242
transform 1 0 5428 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[89\].dly_stg
timestamp 1701704242
transform 1 0 6072 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[90\].dly_stg
timestamp 1701704242
transform 1 0 6624 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[91\].dly_stg
timestamp 1701704242
transform 1 0 7452 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[92\].dly_stg
timestamp 1701704242
transform 1 0 7728 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[93\].dly_stg
timestamp 1701704242
transform 1 0 9016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[94\].dly_stg
timestamp 1701704242
transform 1 0 8740 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[95\].dly_stg
timestamp 1701704242
transform 1 0 10580 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[96\].dly_stg
timestamp 1701704242
transform 1 0 11500 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[97\].dly_stg
timestamp 1701704242
transform 1 0 12328 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[98\].dly_stg
timestamp 1701704242
transform 1 0 13156 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[99\].dly_stg
timestamp 1701704242
transform 1 0 13800 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[100\].dly_stg
timestamp 1701704242
transform 1 0 14076 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[101\].dly_stg
timestamp 1701704242
transform 1 0 14996 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[102\].dly_stg
timestamp 1701704242
transform 1 0 15732 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[103\].dly_stg
timestamp 1701704242
transform -1 0 15732 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[104\].dly_stg
timestamp 1701704242
transform 1 0 16652 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[105\].dly_stg
timestamp 1701704242
transform -1 0 15272 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[106\].dly_stg
timestamp 1701704242
transform 1 0 15640 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[107\].dly_stg
timestamp 1701704242
transform 1 0 16376 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[108\].dly_stg
timestamp 1701704242
transform 1 0 16928 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[109\].dly_stg
timestamp 1701704242
transform 1 0 17204 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[110\].dly_stg
timestamp 1701704242
transform -1 0 17020 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[111\].dly_stg
timestamp 1701704242
transform 1 0 17940 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[112\].dly_stg
timestamp 1701704242
transform 1 0 17388 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[113\].dly_stg
timestamp 1701704242
transform -1 0 18584 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[114\].dly_stg
timestamp 1701704242
transform -1 0 18032 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[115\].dly_stg
timestamp 1701704242
transform 1 0 18308 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[116\].dly_stg
timestamp 1701704242
transform 1 0 17848 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[117\].dly_stg
timestamp 1701704242
transform -1 0 18032 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[118\].dly_stg
timestamp 1701704242
transform 1 0 18768 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[119\].dly_stg
timestamp 1701704242
transform -1 0 18584 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[120\].dly_stg
timestamp 1701704242
transform -1 0 18584 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[121\].dly_stg
timestamp 1701704242
transform -1 0 18492 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[122\].dly_stg
timestamp 1701704242
transform -1 0 18768 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[123\].dly_stg
timestamp 1701704242
transform -1 0 17480 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[124\].dly_stg
timestamp 1701704242
transform -1 0 17848 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[125\].dly_stg
timestamp 1701704242
transform 1 0 18584 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_interleave_n\[126\].dly_stg
timestamp 1701704242
transform -1 0 16744 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  tdc0.g_dly_chain_odd\[0\].dly_stg
timestamp 1701704242
transform -1 0 18308 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[1\].dly_stg
timestamp 1701704242
transform 1 0 16652 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[2\].dly_stg
timestamp 1701704242
transform -1 0 16652 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[3\].dly_stg
timestamp 1701704242
transform -1 0 16376 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[4\].dly_stg
timestamp 1701704242
transform -1 0 15456 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[5\].dly_stg
timestamp 1701704242
transform -1 0 15272 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[6\].dly_stg
timestamp 1701704242
transform -1 0 14720 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[7\].dly_stg
timestamp 1701704242
transform -1 0 14168 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[8\].dly_stg
timestamp 1701704242
transform 1 0 15088 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[9\].dly_stg
timestamp 1701704242
transform -1 0 13432 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[10\].dly_stg
timestamp 1701704242
transform -1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[11\].dly_stg
timestamp 1701704242
transform 1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[12\].dly_stg
timestamp 1701704242
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[13\].dly_stg
timestamp 1701704242
transform -1 0 13248 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[14\].dly_stg
timestamp 1701704242
transform 1 0 12236 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[15\].dly_stg
timestamp 1701704242
transform -1 0 11500 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[16\].dly_stg
timestamp 1701704242
transform -1 0 11316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[17\].dly_stg
timestamp 1701704242
transform -1 0 10856 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[18\].dly_stg
timestamp 1701704242
transform -1 0 11868 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[19\].dly_stg
timestamp 1701704242
transform -1 0 12144 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[20\].dly_stg
timestamp 1701704242
transform 1 0 12052 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[21\].dly_stg
timestamp 1701704242
transform -1 0 13064 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[22\].dly_stg
timestamp 1701704242
transform 1 0 14076 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[23\].dly_stg
timestamp 1701704242
transform 1 0 14260 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[24\].dly_stg
timestamp 1701704242
transform 1 0 14352 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[25\].dly_stg
timestamp 1701704242
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[26\].dly_stg
timestamp 1701704242
transform 1 0 15364 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[27\].dly_stg
timestamp 1701704242
transform -1 0 13432 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[28\].dly_stg
timestamp 1701704242
transform 1 0 14168 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[29\].dly_stg
timestamp 1701704242
transform -1 0 13616 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[30\].dly_stg
timestamp 1701704242
transform -1 0 10580 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[31\].dly_stg
timestamp 1701704242
transform -1 0 7728 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[32\].dly_stg
timestamp 1701704242
transform -1 0 8924 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[33\].dly_stg
timestamp 1701704242
transform -1 0 7452 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[34\].dly_stg
timestamp 1701704242
transform -1 0 6900 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[35\].dly_stg
timestamp 1701704242
transform 1 0 7084 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[36\].dly_stg
timestamp 1701704242
transform -1 0 6808 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[37\].dly_stg
timestamp 1701704242
transform 1 0 6900 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[38\].dly_stg
timestamp 1701704242
transform -1 0 5428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[39\].dly_stg
timestamp 1701704242
transform 1 0 5796 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[40\].dly_stg
timestamp 1701704242
transform -1 0 5704 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[41\].dly_stg
timestamp 1701704242
transform 1 0 4232 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[42\].dly_stg
timestamp 1701704242
transform 1 0 4784 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[43\].dly_stg
timestamp 1701704242
transform -1 0 3772 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[44\].dly_stg
timestamp 1701704242
transform 1 0 3128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[45\].dly_stg
timestamp 1701704242
transform -1 0 2760 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[46\].dly_stg
timestamp 1701704242
transform 1 0 2024 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[47\].dly_stg
timestamp 1701704242
transform -1 0 1472 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[48\].dly_stg
timestamp 1701704242
transform -1 0 1932 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[49\].dly_stg
timestamp 1701704242
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[50\].dly_stg
timestamp 1701704242
transform -1 0 1288 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[51\].dly_stg
timestamp 1701704242
transform -1 0 1748 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[52\].dly_stg
timestamp 1701704242
transform -1 0 2576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[53\].dly_stg
timestamp 1701704242
transform -1 0 2576 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[54\].dly_stg
timestamp 1701704242
transform 1 0 3404 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[55\].dly_stg
timestamp 1701704242
transform -1 0 4140 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[56\].dly_stg
timestamp 1701704242
transform 1 0 5152 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[57\].dly_stg
timestamp 1701704242
transform -1 0 4600 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[58\].dly_stg
timestamp 1701704242
transform 1 0 5980 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[59\].dly_stg
timestamp 1701704242
transform 1 0 5152 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[60\].dly_stg
timestamp 1701704242
transform 1 0 6072 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[61\].dly_stg
timestamp 1701704242
transform 1 0 5796 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[62\].dly_stg
timestamp 1701704242
transform -1 0 6072 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[63\].dly_stg
timestamp 1701704242
transform -1 0 4784 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[64\].dly_stg
timestamp 1701704242
transform -1 0 5796 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[65\].dly_stg
timestamp 1701704242
transform -1 0 4692 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[66\].dly_stg
timestamp 1701704242
transform -1 0 3680 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[67\].dly_stg
timestamp 1701704242
transform -1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[68\].dly_stg
timestamp 1701704242
transform -1 0 4048 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[69\].dly_stg
timestamp 1701704242
transform 1 0 3404 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[70\].dly_stg
timestamp 1701704242
transform -1 0 2576 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[71\].dly_stg
timestamp 1701704242
transform -1 0 2024 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[72\].dly_stg
timestamp 1701704242
transform -1 0 2208 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[73\].dly_stg
timestamp 1701704242
transform 1 0 1656 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[74\].dly_stg
timestamp 1701704242
transform -1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[75\].dly_stg
timestamp 1701704242
transform -1 0 1472 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[76\].dly_stg
timestamp 1701704242
transform 1 0 1840 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[77\].dly_stg
timestamp 1701704242
transform 1 0 1288 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[78\].dly_stg
timestamp 1701704242
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[79\].dly_stg
timestamp 1701704242
transform 1 0 1288 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[80\].dly_stg
timestamp 1701704242
transform 1 0 1564 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[81\].dly_stg
timestamp 1701704242
transform -1 0 2116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[82\].dly_stg
timestamp 1701704242
transform 1 0 1380 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[83\].dly_stg
timestamp 1701704242
transform -1 0 2024 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[84\].dly_stg
timestamp 1701704242
transform 1 0 3036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[85\].dly_stg
timestamp 1701704242
transform -1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[86\].dly_stg
timestamp 1701704242
transform 1 0 3312 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[87\].dly_stg
timestamp 1701704242
transform -1 0 5060 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[88\].dly_stg
timestamp 1701704242
transform 1 0 5152 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[89\].dly_stg
timestamp 1701704242
transform -1 0 6072 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[90\].dly_stg
timestamp 1701704242
transform 1 0 6256 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[91\].dly_stg
timestamp 1701704242
transform -1 0 7360 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[92\].dly_stg
timestamp 1701704242
transform 1 0 7636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[93\].dly_stg
timestamp 1701704242
transform -1 0 8648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[94\].dly_stg
timestamp 1701704242
transform 1 0 8464 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[95\].dly_stg
timestamp 1701704242
transform 1 0 10580 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[96\].dly_stg
timestamp 1701704242
transform 1 0 10948 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[97\].dly_stg
timestamp 1701704242
transform -1 0 12052 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[98\].dly_stg
timestamp 1701704242
transform -1 0 12972 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[99\].dly_stg
timestamp 1701704242
transform -1 0 13800 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[100\].dly_stg
timestamp 1701704242
transform -1 0 13800 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[101\].dly_stg
timestamp 1701704242
transform 1 0 14904 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[102\].dly_stg
timestamp 1701704242
transform 1 0 14444 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[103\].dly_stg
timestamp 1701704242
transform 1 0 16100 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[104\].dly_stg
timestamp 1701704242
transform -1 0 16376 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[105\].dly_stg
timestamp 1701704242
transform -1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[106\].dly_stg
timestamp 1701704242
transform 1 0 15272 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[107\].dly_stg
timestamp 1701704242
transform -1 0 15640 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[108\].dly_stg
timestamp 1701704242
transform -1 0 16928 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[109\].dly_stg
timestamp 1701704242
transform -1 0 16192 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[110\].dly_stg
timestamp 1701704242
transform -1 0 17112 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[111\].dly_stg
timestamp 1701704242
transform -1 0 17940 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[112\].dly_stg
timestamp 1701704242
transform -1 0 16744 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[113\].dly_stg
timestamp 1701704242
transform -1 0 17572 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[114\].dly_stg
timestamp 1701704242
transform 1 0 18676 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[115\].dly_stg
timestamp 1701704242
transform -1 0 17756 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[116\].dly_stg
timestamp 1701704242
transform 1 0 17756 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[117\].dly_stg
timestamp 1701704242
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[118\].dly_stg
timestamp 1701704242
transform 1 0 18768 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[119\].dly_stg
timestamp 1701704242
transform 1 0 18676 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[120\].dly_stg
timestamp 1701704242
transform 1 0 18676 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[121\].dly_stg
timestamp 1701704242
transform 1 0 18860 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[122\].dly_stg
timestamp 1701704242
transform -1 0 18216 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[123\].dly_stg
timestamp 1701704242
transform -1 0 18032 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[124\].dly_stg
timestamp 1701704242
transform -1 0 17756 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[125\].dly_stg
timestamp 1701704242
transform -1 0 18124 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[126\].dly_stg
timestamp 1701704242
transform 1 0 18124 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[127\].dly_stg
timestamp 1701704242
transform 1 0 18676 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  tdc0.g_dly_chain_odd\[128\].dly_stg
timestamp 1701704242
transform 1 0 16744 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_12 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18860 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_13
timestamp 1701704242
transform -1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_14
timestamp 1701704242
transform -1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_15
timestamp 1701704242
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_16
timestamp 1701704242
transform 1 0 18860 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_17
timestamp 1701704242
transform 1 0 18860 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_18
timestamp 1701704242
transform 1 0 18860 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_19
timestamp 1701704242
transform -1 0 1104 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_20
timestamp 1701704242
transform -1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_21
timestamp 1701704242
transform 1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_22
timestamp 1701704242
transform 1 0 18860 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_23
timestamp 1701704242
transform -1 0 2668 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_24
timestamp 1701704242
transform -1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_25
timestamp 1701704242
transform 1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_26
timestamp 1701704242
transform -1 0 1656 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_27
timestamp 1701704242
transform -1 0 1656 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  wire8
timestamp 1701704242
transform 1 0 12144 0 -1 5984
box -38 -48 406 592
<< labels >>
flabel metal4 s 5106 496 5426 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9821 496 10141 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14536 496 14856 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 19251 496 19571 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2749 496 3069 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7464 496 7784 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12179 496 12499 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 16894 496 17214 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 16328 400 16448 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 18 0 74 400 0 FreeSans 224 90 0 0 ena
port 3 nsew signal input
flabel metal2 s 4526 0 4582 400 0 FreeSans 224 90 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 19600 11568 20000 11688 0 FreeSans 480 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal2 s 3882 0 3938 400 0 FreeSans 224 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal2 s 3238 0 3294 400 0 FreeSans 224 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal2 s 12898 0 12954 400 0 FreeSans 224 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal2 s 10322 0 10378 400 0 FreeSans 224 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal2 s 12254 0 12310 400 0 FreeSans 224 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal2 s 11610 0 11666 400 0 FreeSans 224 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal2 s 2594 0 2650 400 0 FreeSans 224 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal2 s 7102 0 7158 400 0 FreeSans 224 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal2 s 6458 0 6514 400 0 FreeSans 224 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal2 s 5814 0 5870 400 0 FreeSans 224 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal2 s 5170 0 5226 400 0 FreeSans 224 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal2 s 9678 0 9734 400 0 FreeSans 224 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal2 s 9034 0 9090 400 0 FreeSans 224 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal2 s 8390 0 8446 400 0 FreeSans 224 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal2 s 7746 0 7802 400 0 FreeSans 224 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 19600 17008 20000 17128 0 FreeSans 480 0 0 0 uio_oe[0]
port 21 nsew signal tristate
flabel metal3 s 0 19728 400 19848 0 FreeSans 480 0 0 0 uio_oe[1]
port 22 nsew signal tristate
flabel metal3 s 0 17008 400 17128 0 FreeSans 480 0 0 0 uio_oe[2]
port 23 nsew signal tristate
flabel metal3 s 19600 8 20000 128 0 FreeSans 480 0 0 0 uio_oe[3]
port 24 nsew signal tristate
flabel metal3 s 19600 18368 20000 18488 0 FreeSans 480 0 0 0 uio_oe[4]
port 25 nsew signal tristate
flabel metal3 s 19600 1368 20000 1488 0 FreeSans 480 0 0 0 uio_oe[5]
port 26 nsew signal tristate
flabel metal3 s 19600 688 20000 808 0 FreeSans 480 0 0 0 uio_oe[6]
port 27 nsew signal tristate
flabel metal2 s 662 0 718 400 0 FreeSans 224 90 0 0 uio_oe[7]
port 28 nsew signal tristate
flabel metal3 s 0 18368 400 18488 0 FreeSans 480 0 0 0 uio_out[0]
port 29 nsew signal tristate
flabel metal3 s 19600 2048 20000 2168 0 FreeSans 480 0 0 0 uio_out[1]
port 30 nsew signal tristate
flabel metal3 s 19600 17688 20000 17808 0 FreeSans 480 0 0 0 uio_out[2]
port 31 nsew signal tristate
flabel metal2 s 1950 0 2006 400 0 FreeSans 224 90 0 0 uio_out[3]
port 32 nsew signal tristate
flabel metal3 s 0 17688 400 17808 0 FreeSans 480 0 0 0 uio_out[4]
port 33 nsew signal tristate
flabel metal3 s 19600 19048 20000 19168 0 FreeSans 480 0 0 0 uio_out[5]
port 34 nsew signal tristate
flabel metal3 s 0 19048 400 19168 0 FreeSans 480 0 0 0 uio_out[6]
port 35 nsew signal tristate
flabel metal2 s 1306 0 1362 400 0 FreeSans 224 90 0 0 uio_out[7]
port 36 nsew signal tristate
flabel metal3 s 19600 12248 20000 12368 0 FreeSans 480 0 0 0 uo_out[0]
port 37 nsew signal tristate
flabel metal3 s 19600 8168 20000 8288 0 FreeSans 480 0 0 0 uo_out[1]
port 38 nsew signal tristate
flabel metal3 s 19600 12928 20000 13048 0 FreeSans 480 0 0 0 uo_out[2]
port 39 nsew signal tristate
flabel metal3 s 19600 10208 20000 10328 0 FreeSans 480 0 0 0 uo_out[3]
port 40 nsew signal tristate
flabel metal3 s 19600 8848 20000 8968 0 FreeSans 480 0 0 0 uo_out[4]
port 41 nsew signal tristate
flabel metal3 s 19600 10888 20000 11008 0 FreeSans 480 0 0 0 uo_out[5]
port 42 nsew signal tristate
flabel metal3 s 19600 9528 20000 9648 0 FreeSans 480 0 0 0 uo_out[6]
port 43 nsew signal tristate
flabel metal2 s 11610 19600 11666 20000 0 FreeSans 224 90 0 0 uo_out[7]
port 44 nsew signal tristate
rlabel via1 10061 19040 10061 19040 0 VGND
rlabel metal1 9982 18496 9982 18496 0 VPWR
rlabel metal1 10534 8330 10534 8330 0 _000_
rlabel metal1 14076 7514 14076 7514 0 _001_
rlabel metal1 10166 8330 10166 8330 0 _002_
rlabel metal1 12282 8432 12282 8432 0 _003_
rlabel metal3 12282 8364 12282 8364 0 _004_
rlabel metal1 14950 8976 14950 8976 0 _005_
rlabel metal2 12558 8092 12558 8092 0 _006_
rlabel metal1 8965 12750 8965 12750 0 _007_
rlabel metal1 14858 9010 14858 9010 0 _008_
rlabel metal2 13846 8126 13846 8126 0 _009_
rlabel metal1 6854 7344 6854 7344 0 _010_
rlabel metal1 14122 8806 14122 8806 0 _011_
rlabel metal1 10672 9010 10672 9010 0 _012_
rlabel metal1 14030 6222 14030 6222 0 _013_
rlabel metal1 14352 9010 14352 9010 0 _014_
rlabel via2 14950 7939 14950 7939 0 _015_
rlabel metal1 9798 10574 9798 10574 0 _016_
rlabel metal2 14122 7174 14122 7174 0 _017_
rlabel metal1 15502 9078 15502 9078 0 _018_
rlabel metal2 9752 5134 9752 5134 0 _019_
rlabel metal1 9062 6120 9062 6120 0 _020_
rlabel metal1 9384 6358 9384 6358 0 _021_
rlabel metal2 10626 12891 10626 12891 0 _022_
rlabel metal1 8878 6834 8878 6834 0 _023_
rlabel metal1 8326 13158 8326 13158 0 _024_
rlabel metal2 9430 7446 9430 7446 0 _025_
rlabel metal2 9614 6358 9614 6358 0 _026_
rlabel metal1 9614 6664 9614 6664 0 _027_
rlabel metal2 8878 8602 8878 8602 0 _028_
rlabel metal1 8234 8330 8234 8330 0 _029_
rlabel metal1 9016 8398 9016 8398 0 _030_
rlabel metal1 9568 8602 9568 8602 0 _031_
rlabel metal2 9752 17068 9752 17068 0 _032_
rlabel metal1 9476 10982 9476 10982 0 _033_
rlabel metal2 9706 10948 9706 10948 0 _034_
rlabel metal2 9522 6171 9522 6171 0 _035_
rlabel metal1 9982 11288 9982 11288 0 _036_
rlabel metal1 11730 10642 11730 10642 0 _037_
rlabel metal2 9982 2397 9982 2397 0 _038_
rlabel metal1 11638 10506 11638 10506 0 _039_
rlabel metal2 11408 15538 11408 15538 0 _040_
rlabel metal1 11868 10778 11868 10778 0 _041_
rlabel metal1 6118 13158 6118 13158 0 _042_
rlabel metal1 11730 9690 11730 9690 0 _043_
rlabel metal1 12098 9894 12098 9894 0 _044_
rlabel metal1 15134 8024 15134 8024 0 _045_
rlabel metal1 12880 9010 12880 9010 0 _046_
rlabel metal1 14398 7854 14398 7854 0 _047_
rlabel metal1 8786 8024 8786 8024 0 _048_
rlabel metal1 13294 7956 13294 7956 0 _049_
rlabel metal2 13110 6222 13110 6222 0 _050_
rlabel metal1 13386 7718 13386 7718 0 _051_
rlabel metal2 13754 10608 13754 10608 0 _052_
rlabel metal2 11408 17204 11408 17204 0 _053_
rlabel metal2 10534 11492 10534 11492 0 _054_
rlabel metal1 10948 5338 10948 5338 0 _055_
rlabel metal1 11638 11798 11638 11798 0 _056_
rlabel metal1 10856 12410 10856 12410 0 _057_
rlabel metal1 10120 12614 10120 12614 0 _058_
rlabel metal1 10994 12818 10994 12818 0 _059_
rlabel via2 10626 2635 10626 2635 0 _060_
rlabel metal1 11362 12614 11362 12614 0 _061_
rlabel metal2 9384 5882 9384 5882 0 _062_
rlabel metal1 16008 6426 16008 6426 0 _063_
rlabel metal1 16238 5882 16238 5882 0 _064_
rlabel metal2 15594 6018 15594 6018 0 _065_
rlabel metal1 16284 6358 16284 6358 0 _066_
rlabel metal2 8050 12585 8050 12585 0 _067_
rlabel metal1 8096 12954 8096 12954 0 _068_
rlabel metal1 8464 12818 8464 12818 0 _069_
rlabel metal1 4600 12614 4600 12614 0 _070_
rlabel metal1 8939 12104 8939 12104 0 _071_
rlabel metal2 12006 11254 12006 11254 0 _072_
rlabel metal1 11592 8806 11592 8806 0 _073_
rlabel metal1 13478 5338 13478 5338 0 _074_
rlabel metal1 11730 8602 11730 8602 0 _075_
rlabel metal2 12558 9350 12558 9350 0 _076_
rlabel metal1 5336 9146 5336 9146 0 _077_
rlabel metal1 10028 9894 10028 9894 0 _078_
rlabel metal2 9614 9588 9614 9588 0 _079_
rlabel metal1 11592 4794 11592 4794 0 _080_
rlabel metal1 12696 9486 12696 9486 0 _081_
rlabel via2 9706 5627 9706 5627 0 _082_
rlabel metal1 14904 5338 14904 5338 0 _083_
rlabel metal1 15824 5202 15824 5202 0 _084_
rlabel metal1 15502 5134 15502 5134 0 _085_
rlabel metal1 14766 5270 14766 5270 0 _086_
rlabel metal2 7130 12585 7130 12585 0 _087_
rlabel metal1 6900 12954 6900 12954 0 _088_
rlabel metal1 12834 13328 12834 13328 0 _089_
rlabel metal1 6164 12682 6164 12682 0 _090_
rlabel metal1 7636 12954 7636 12954 0 _091_
rlabel metal2 9430 6392 9430 6392 0 _092_
rlabel metal2 16422 7990 16422 7990 0 _093_
rlabel metal2 16330 7684 16330 7684 0 _094_
rlabel metal1 16146 7888 16146 7888 0 _095_
rlabel metal2 16606 9044 16606 9044 0 _096_
rlabel metal2 6394 8228 6394 8228 0 _097_
rlabel metal2 6578 14484 6578 14484 0 _098_
rlabel metal1 7360 10642 7360 10642 0 _099_
rlabel metal1 5520 10506 5520 10506 0 _100_
rlabel metal1 6946 10472 6946 10472 0 _101_
rlabel metal3 1395 16388 1395 16388 0 clk
rlabel metal1 13386 14552 13386 14552 0 clknet_0_clk
rlabel metal1 3450 1258 3450 1258 0 clknet_4_0_0_clk
rlabel metal1 17664 1870 17664 1870 0 clknet_4_10_0_clk
rlabel metal1 16514 9554 16514 9554 0 clknet_4_11_0_clk
rlabel metal1 12374 12308 12374 12308 0 clknet_4_12_0_clk
rlabel metal1 14536 17646 14536 17646 0 clknet_4_13_0_clk
rlabel metal1 14950 10098 14950 10098 0 clknet_4_14_0_clk
rlabel metal1 15686 16150 15686 16150 0 clknet_4_15_0_clk
rlabel metal1 1334 8942 1334 8942 0 clknet_4_1_0_clk
rlabel metal2 6578 1904 6578 1904 0 clknet_4_2_0_clk
rlabel metal1 7636 9010 7636 9010 0 clknet_4_3_0_clk
rlabel metal1 1196 13362 1196 13362 0 clknet_4_4_0_clk
rlabel metal1 2024 17646 2024 17646 0 clknet_4_5_0_clk
rlabel metal1 5382 12886 5382 12886 0 clknet_4_6_0_clk
rlabel metal1 8740 14382 8740 14382 0 clknet_4_7_0_clk
rlabel metal1 10902 1938 10902 1938 0 clknet_4_8_0_clk
rlabel metal2 13018 4624 13018 4624 0 clknet_4_9_0_clk
rlabel metal2 18630 12240 18630 12240 0 net1
rlabel metal1 13248 7446 13248 7446 0 net10
rlabel metal1 15134 13804 15134 13804 0 net11
rlabel metal2 19090 16847 19090 16847 0 net12
rlabel metal2 1150 19261 1150 19261 0 net13
rlabel metal3 590 17068 590 17068 0 net14
rlabel metal3 19144 68 19144 68 0 net15
rlabel metal3 19420 18428 19420 18428 0 net16
rlabel metal3 19420 1428 19420 1428 0 net17
rlabel metal3 19420 748 19420 748 0 net18
rlabel metal2 690 568 690 568 0 net19
rlabel metal2 11914 3604 11914 3604 0 net2
rlabel metal3 590 18428 590 18428 0 net20
rlabel metal3 19420 2108 19420 2108 0 net21
rlabel metal3 19420 17748 19420 17748 0 net22
rlabel metal2 1978 636 1978 636 0 net23
rlabel metal3 590 17748 590 17748 0 net24
rlabel via2 18538 18819 18538 18819 0 net25
rlabel metal1 1104 18802 1104 18802 0 net26
rlabel metal2 1334 568 1334 568 0 net27
rlabel metal1 11362 9044 11362 9044 0 net28
rlabel metal1 10074 6834 10074 6834 0 net3
rlabel metal1 11362 5032 11362 5032 0 net4
rlabel metal1 11914 5134 11914 5134 0 net5
rlabel metal1 10350 15912 10350 15912 0 net6
rlabel metal2 10994 6409 10994 6409 0 net7
rlabel metal1 12236 5746 12236 5746 0 net8
rlabel metal2 9430 17544 9430 17544 0 net9
rlabel metal1 15962 12274 15962 12274 0 tdc0.o_result\[0\]
rlabel metal1 14444 3706 14444 3706 0 tdc0.o_result\[100\]
rlabel metal1 18078 1530 18078 1530 0 tdc0.o_result\[101\]
rlabel metal1 11132 3162 11132 3162 0 tdc0.o_result\[102\]
rlabel metal1 18078 2074 18078 2074 0 tdc0.o_result\[103\]
rlabel metal2 16698 4148 16698 4148 0 tdc0.o_result\[104\]
rlabel metal1 13018 3944 13018 3944 0 tdc0.o_result\[105\]
rlabel metal2 14490 6273 14490 6273 0 tdc0.o_result\[106\]
rlabel metal1 16008 4794 16008 4794 0 tdc0.o_result\[107\]
rlabel metal1 8188 4454 8188 4454 0 tdc0.o_result\[108\]
rlabel metal1 10212 4250 10212 4250 0 tdc0.o_result\[109\]
rlabel metal1 14398 5644 14398 5644 0 tdc0.o_result\[10\]
rlabel metal1 17204 3162 17204 3162 0 tdc0.o_result\[110\]
rlabel metal1 9936 4794 9936 4794 0 tdc0.o_result\[111\]
rlabel metal1 17572 3706 17572 3706 0 tdc0.o_result\[112\]
rlabel metal1 13294 4658 13294 4658 0 tdc0.o_result\[113\]
rlabel metal1 17305 4794 17305 4794 0 tdc0.o_result\[114\]
rlabel metal1 16192 7174 16192 7174 0 tdc0.o_result\[115\]
rlabel metal2 9614 6817 9614 6817 0 tdc0.o_result\[116\]
rlabel metal1 18722 8976 18722 8976 0 tdc0.o_result\[117\]
rlabel metal1 15962 7956 15962 7956 0 tdc0.o_result\[118\]
rlabel metal2 18262 8874 18262 8874 0 tdc0.o_result\[119\]
rlabel metal1 14996 7990 14996 7990 0 tdc0.o_result\[11\]
rlabel via2 8694 12699 8694 12699 0 tdc0.o_result\[120\]
rlabel metal1 13590 8568 13590 8568 0 tdc0.o_result\[121\]
rlabel metal1 16928 14518 16928 14518 0 tdc0.o_result\[122\]
rlabel metal2 8694 11985 8694 11985 0 tdc0.o_result\[123\]
rlabel metal1 16192 13838 16192 13838 0 tdc0.o_result\[124\]
rlabel metal1 10580 15946 10580 15946 0 tdc0.o_result\[125\]
rlabel metal1 16422 17680 16422 17680 0 tdc0.o_result\[126\]
rlabel metal1 13202 15980 13202 15980 0 tdc0.o_result\[127\]
rlabel metal1 15042 13974 15042 13974 0 tdc0.o_result\[12\]
rlabel metal1 10764 10642 10764 10642 0 tdc0.o_result\[13\]
rlabel metal1 11178 14246 11178 14246 0 tdc0.o_result\[14\]
rlabel metal2 10534 12937 10534 12937 0 tdc0.o_result\[15\]
rlabel metal1 7866 17136 7866 17136 0 tdc0.o_result\[16\]
rlabel metal2 10350 14960 10350 14960 0 tdc0.o_result\[17\]
rlabel metal1 6394 17782 6394 17782 0 tdc0.o_result\[18\]
rlabel metal1 6394 16728 6394 16728 0 tdc0.o_result\[19\]
rlabel metal1 12834 9486 12834 9486 0 tdc0.o_result\[1\]
rlabel metal2 12926 15198 12926 15198 0 tdc0.o_result\[20\]
rlabel metal1 10166 17782 10166 17782 0 tdc0.o_result\[21\]
rlabel metal1 16652 17714 16652 17714 0 tdc0.o_result\[22\]
rlabel metal2 11270 17782 11270 17782 0 tdc0.o_result\[23\]
rlabel metal1 16146 17578 16146 17578 0 tdc0.o_result\[24\]
rlabel metal2 11546 15878 11546 15878 0 tdc0.o_result\[25\]
rlabel metal1 16284 15334 16284 15334 0 tdc0.o_result\[26\]
rlabel metal2 16330 9809 16330 9809 0 tdc0.o_result\[27\]
rlabel metal1 13800 14790 13800 14790 0 tdc0.o_result\[28\]
rlabel metal2 9890 12041 9890 12041 0 tdc0.o_result\[29\]
rlabel metal1 14674 12818 14674 12818 0 tdc0.o_result\[2\]
rlabel metal1 10534 8942 10534 8942 0 tdc0.o_result\[30\]
rlabel metal1 9706 12784 9706 12784 0 tdc0.o_result\[31\]
rlabel metal1 8510 5814 8510 5814 0 tdc0.o_result\[32\]
rlabel metal1 9338 9010 9338 9010 0 tdc0.o_result\[33\]
rlabel via2 9430 5763 9430 5763 0 tdc0.o_result\[34\]
rlabel metal1 8556 6902 8556 6902 0 tdc0.o_result\[35\]
rlabel metal1 7268 13362 7268 13362 0 tdc0.o_result\[36\]
rlabel metal1 9982 16014 9982 16014 0 tdc0.o_result\[37\]
rlabel metal2 6394 14076 6394 14076 0 tdc0.o_result\[38\]
rlabel metal2 10810 16388 10810 16388 0 tdc0.o_result\[39\]
rlabel metal2 16422 10234 16422 10234 0 tdc0.o_result\[3\]
rlabel metal1 7268 17102 7268 17102 0 tdc0.o_result\[40\]
rlabel metal1 11270 15572 11270 15572 0 tdc0.o_result\[41\]
rlabel metal1 5888 17714 5888 17714 0 tdc0.o_result\[42\]
rlabel viali 6128 16626 6128 16626 0 tdc0.o_result\[43\]
rlabel metal1 6900 15334 6900 15334 0 tdc0.o_result\[44\]
rlabel metal1 10350 17680 10350 17680 0 tdc0.o_result\[45\]
rlabel metal1 4646 9452 4646 9452 0 tdc0.o_result\[46\]
rlabel metal1 3680 17306 3680 17306 0 tdc0.o_result\[47\]
rlabel metal1 2668 12342 2668 12342 0 tdc0.o_result\[48\]
rlabel metal1 4002 14246 4002 14246 0 tdc0.o_result\[49\]
rlabel metal1 14766 9044 14766 9044 0 tdc0.o_result\[4\]
rlabel metal2 3542 12784 3542 12784 0 tdc0.o_result\[50\]
rlabel metal1 2990 10506 2990 10506 0 tdc0.o_result\[51\]
rlabel metal1 7774 13294 7774 13294 0 tdc0.o_result\[52\]
rlabel metal1 10074 10642 10074 10642 0 tdc0.o_result\[53\]
rlabel metal2 6118 13430 6118 13430 0 tdc0.o_result\[54\]
rlabel metal1 10166 11152 10166 11152 0 tdc0.o_result\[55\]
rlabel metal1 8418 12716 8418 12716 0 tdc0.o_result\[56\]
rlabel metal1 8832 12274 8832 12274 0 tdc0.o_result\[57\]
rlabel metal2 7314 6477 7314 6477 0 tdc0.o_result\[58\]
rlabel metal2 7590 11492 7590 11492 0 tdc0.o_result\[59\]
rlabel metal1 11546 11084 11546 11084 0 tdc0.o_result\[5\]
rlabel metal1 12926 9384 12926 9384 0 tdc0.o_result\[60\]
rlabel metal1 9338 11322 9338 11322 0 tdc0.o_result\[61\]
rlabel metal2 11086 9724 11086 9724 0 tdc0.o_result\[62\]
rlabel metal2 9246 12580 9246 12580 0 tdc0.o_result\[63\]
rlabel metal1 6440 7310 6440 7310 0 tdc0.o_result\[64\]
rlabel metal1 8280 8534 8280 8534 0 tdc0.o_result\[65\]
rlabel metal1 5612 6222 5612 6222 0 tdc0.o_result\[66\]
rlabel metal1 5566 4794 5566 4794 0 tdc0.o_result\[67\]
rlabel metal1 7222 5338 7222 5338 0 tdc0.o_result\[68\]
rlabel metal1 9476 5066 9476 5066 0 tdc0.o_result\[69\]
rlabel metal2 12466 9384 12466 9384 0 tdc0.o_result\[6\]
rlabel metal1 5014 8806 5014 8806 0 tdc0.o_result\[70\]
rlabel metal1 10626 5134 10626 5134 0 tdc0.o_result\[71\]
rlabel metal1 2530 11866 2530 11866 0 tdc0.o_result\[72\]
rlabel metal2 2990 8857 2990 8857 0 tdc0.o_result\[73\]
rlabel metal1 3220 12274 3220 12274 0 tdc0.o_result\[74\]
rlabel metal1 2484 9690 2484 9690 0 tdc0.o_result\[75\]
rlabel metal1 9062 6800 9062 6800 0 tdc0.o_result\[76\]
rlabel metal1 6486 9928 6486 9928 0 tdc0.o_result\[77\]
rlabel metal1 7314 4692 7314 4692 0 tdc0.o_result\[78\]
rlabel metal1 3082 5270 3082 5270 0 tdc0.o_result\[79\]
rlabel metal1 12558 11798 12558 11798 0 tdc0.o_result\[7\]
rlabel metal1 4186 3366 4186 3366 0 tdc0.o_result\[80\]
rlabel metal1 3956 3162 3956 3162 0 tdc0.o_result\[81\]
rlabel metal1 3772 1530 3772 1530 0 tdc0.o_result\[82\]
rlabel metal1 4968 3706 4968 3706 0 tdc0.o_result\[83\]
rlabel metal2 4830 1683 4830 1683 0 tdc0.o_result\[84\]
rlabel metal1 6118 1768 6118 1768 0 tdc0.o_result\[85\]
rlabel metal1 7314 3910 7314 3910 0 tdc0.o_result\[86\]
rlabel metal2 7406 2176 7406 2176 0 tdc0.o_result\[87\]
rlabel metal1 8004 4794 8004 4794 0 tdc0.o_result\[88\]
rlabel metal1 8326 2346 8326 2346 0 tdc0.o_result\[89\]
rlabel metal1 14770 5746 14770 5746 0 tdc0.o_result\[8\]
rlabel metal1 8648 3706 8648 3706 0 tdc0.o_result\[90\]
rlabel metal2 8372 6834 8372 6834 0 tdc0.o_result\[91\]
rlabel metal1 8464 3910 8464 3910 0 tdc0.o_result\[92\]
rlabel metal1 9430 2448 9430 2448 0 tdc0.o_result\[93\]
rlabel metal1 10304 9010 10304 9010 0 tdc0.o_result\[94\]
rlabel metal1 10166 2482 10166 2482 0 tdc0.o_result\[95\]
rlabel metal1 14812 2278 14812 2278 0 tdc0.o_result\[96\]
rlabel metal1 12236 2074 12236 2074 0 tdc0.o_result\[97\]
rlabel metal1 14306 2618 14306 2618 0 tdc0.o_result\[98\]
rlabel metal1 14904 1530 14904 1530 0 tdc0.o_result\[99\]
rlabel metal1 11224 9078 11224 9078 0 tdc0.o_result\[9\]
rlabel metal1 13652 1394 13652 1394 0 tdc0.w_dly_sig\[100\]
rlabel metal1 13248 1870 13248 1870 0 tdc0.w_dly_sig\[101\]
rlabel metal1 14766 1190 14766 1190 0 tdc0.w_dly_sig\[102\]
rlabel metal1 13938 2074 13938 2074 0 tdc0.w_dly_sig\[103\]
rlabel metal1 16820 1802 16820 1802 0 tdc0.w_dly_sig\[104\]
rlabel metal1 15911 1802 15911 1802 0 tdc0.w_dly_sig\[105\]
rlabel metal1 16100 2278 16100 2278 0 tdc0.w_dly_sig\[106\]
rlabel metal1 14582 3570 14582 3570 0 tdc0.w_dly_sig\[107\]
rlabel metal1 15456 4046 15456 4046 0 tdc0.w_dly_sig\[108\]
rlabel metal1 14770 3706 14770 3706 0 tdc0.w_dly_sig\[109\]
rlabel metal1 13570 12954 13570 12954 0 tdc0.w_dly_sig\[10\]
rlabel metal1 15134 3978 15134 3978 0 tdc0.w_dly_sig\[110\]
rlabel metal1 17756 2482 17756 2482 0 tdc0.w_dly_sig\[111\]
rlabel metal1 10580 4250 10580 4250 0 tdc0.w_dly_sig\[112\]
rlabel metal1 17756 2618 17756 2618 0 tdc0.w_dly_sig\[113\]
rlabel metal1 17250 4726 17250 4726 0 tdc0.w_dly_sig\[114\]
rlabel metal1 18588 4658 18588 4658 0 tdc0.w_dly_sig\[115\]
rlabel metal1 17392 7310 17392 7310 0 tdc0.w_dly_sig\[116\]
rlabel metal1 18538 6290 18538 6290 0 tdc0.w_dly_sig\[117\]
rlabel metal1 17015 9078 17015 9078 0 tdc0.w_dly_sig\[118\]
rlabel metal1 18354 11662 18354 11662 0 tdc0.w_dly_sig\[119\]
rlabel metal1 13570 13158 13570 13158 0 tdc0.w_dly_sig\[11\]
rlabel metal1 17158 9418 17158 9418 0 tdc0.w_dly_sig\[120\]
rlabel metal1 18860 14042 18860 14042 0 tdc0.w_dly_sig\[121\]
rlabel metal1 18952 15130 18952 15130 0 tdc0.w_dly_sig\[122\]
rlabel metal1 18446 15572 18446 15572 0 tdc0.w_dly_sig\[123\]
rlabel metal1 17664 15334 17664 15334 0 tdc0.w_dly_sig\[124\]
rlabel metal1 17572 16218 17572 16218 0 tdc0.w_dly_sig\[125\]
rlabel metal1 18082 16626 18082 16626 0 tdc0.w_dly_sig\[126\]
rlabel metal1 17066 17034 17066 17034 0 tdc0.w_dly_sig\[127\]
rlabel metal1 18364 17714 18364 17714 0 tdc0.w_dly_sig\[128\]
rlabel metal1 17802 17306 17802 17306 0 tdc0.w_dly_sig\[129\]
rlabel metal1 14025 8398 14025 8398 0 tdc0.w_dly_sig\[12\]
rlabel metal1 13984 13906 13984 13906 0 tdc0.w_dly_sig\[13\]
rlabel metal1 12581 15538 12581 15538 0 tdc0.w_dly_sig\[14\]
rlabel metal1 11592 16014 11592 16014 0 tdc0.w_dly_sig\[15\]
rlabel metal1 11224 16490 11224 16490 0 tdc0.w_dly_sig\[16\]
rlabel metal1 8372 17102 8372 17102 0 tdc0.w_dly_sig\[17\]
rlabel metal1 9660 17102 9660 17102 0 tdc0.w_dly_sig\[18\]
rlabel metal2 8510 17714 8510 17714 0 tdc0.w_dly_sig\[19\]
rlabel metal1 14950 12240 14950 12240 0 tdc0.w_dly_sig\[1\]
rlabel metal2 9614 17680 9614 17680 0 tdc0.w_dly_sig\[20\]
rlabel metal2 12558 18496 12558 18496 0 tdc0.w_dly_sig\[21\]
rlabel metal1 13754 18836 13754 18836 0 tdc0.w_dly_sig\[22\]
rlabel metal1 13708 18938 13708 18938 0 tdc0.w_dly_sig\[23\]
rlabel metal1 14168 17850 14168 17850 0 tdc0.w_dly_sig\[24\]
rlabel metal1 14618 17714 14618 17714 0 tdc0.w_dly_sig\[25\]
rlabel metal2 15042 16575 15042 16575 0 tdc0.w_dly_sig\[26\]
rlabel metal1 14766 16694 14766 16694 0 tdc0.w_dly_sig\[27\]
rlabel metal1 14122 15504 14122 15504 0 tdc0.w_dly_sig\[28\]
rlabel metal1 13110 15504 13110 15504 0 tdc0.w_dly_sig\[29\]
rlabel metal2 17710 11016 17710 11016 0 tdc0.w_dly_sig\[2\]
rlabel metal1 13340 15674 13340 15674 0 tdc0.w_dly_sig\[30\]
rlabel metal2 9154 14042 9154 14042 0 tdc0.w_dly_sig\[31\]
rlabel metal1 8694 14960 8694 14960 0 tdc0.w_dly_sig\[32\]
rlabel metal1 8280 13974 8280 13974 0 tdc0.w_dly_sig\[33\]
rlabel metal1 7866 13872 7866 13872 0 tdc0.w_dly_sig\[34\]
rlabel metal1 6716 14246 6716 14246 0 tdc0.w_dly_sig\[35\]
rlabel metal1 7590 13838 7590 13838 0 tdc0.w_dly_sig\[36\]
rlabel metal1 6578 15538 6578 15538 0 tdc0.w_dly_sig\[37\]
rlabel metal1 8142 15980 8142 15980 0 tdc0.w_dly_sig\[38\]
rlabel metal1 5653 14858 5653 14858 0 tdc0.w_dly_sig\[39\]
rlabel metal1 15880 13362 15880 13362 0 tdc0.w_dly_sig\[3\]
rlabel metal1 8142 16218 8142 16218 0 tdc0.w_dly_sig\[40\]
rlabel metal2 5014 16830 5014 16830 0 tdc0.w_dly_sig\[41\]
rlabel metal2 6854 16184 6854 16184 0 tdc0.w_dly_sig\[42\]
rlabel metal1 4784 17306 4784 17306 0 tdc0.w_dly_sig\[43\]
rlabel metal1 2530 16524 2530 16524 0 tdc0.w_dly_sig\[44\]
rlabel metal1 3496 16762 3496 16762 0 tdc0.w_dly_sig\[45\]
rlabel metal1 1794 17714 1794 17714 0 tdc0.w_dly_sig\[46\]
rlabel metal1 2622 16014 2622 16014 0 tdc0.w_dly_sig\[47\]
rlabel via1 1881 17102 1881 17102 0 tdc0.w_dly_sig\[48\]
rlabel metal1 1794 15606 1794 15606 0 tdc0.w_dly_sig\[49\]
rlabel metal1 15134 11220 15134 11220 0 tdc0.w_dly_sig\[4\]
rlabel metal1 2336 14450 2336 14450 0 tdc0.w_dly_sig\[50\]
rlabel metal1 1656 14450 1656 14450 0 tdc0.w_dly_sig\[51\]
rlabel metal1 1518 14042 1518 14042 0 tdc0.w_dly_sig\[52\]
rlabel metal1 2484 13702 2484 13702 0 tdc0.w_dly_sig\[53\]
rlabel metal1 2484 12614 2484 12614 0 tdc0.w_dly_sig\[54\]
rlabel via1 4549 13362 4549 13362 0 tdc0.w_dly_sig\[55\]
rlabel metal2 4002 11866 4002 11866 0 tdc0.w_dly_sig\[56\]
rlabel metal1 4876 12818 4876 12818 0 tdc0.w_dly_sig\[57\]
rlabel metal1 4738 11662 4738 11662 0 tdc0.w_dly_sig\[58\]
rlabel metal1 5842 9418 5842 9418 0 tdc0.w_dly_sig\[59\]
rlabel metal1 14674 10608 14674 10608 0 tdc0.w_dly_sig\[5\]
rlabel metal1 5474 11186 5474 11186 0 tdc0.w_dly_sig\[60\]
rlabel metal1 6210 9452 6210 9452 0 tdc0.w_dly_sig\[61\]
rlabel metal1 7728 10574 7728 10574 0 tdc0.w_dly_sig\[62\]
rlabel metal1 6578 9690 6578 9690 0 tdc0.w_dly_sig\[63\]
rlabel metal1 7314 10778 7314 10778 0 tdc0.w_dly_sig\[64\]
rlabel metal1 5520 8262 5520 8262 0 tdc0.w_dly_sig\[65\]
rlabel via1 6297 8398 6297 8398 0 tdc0.w_dly_sig\[66\]
rlabel metal2 4922 7548 4922 7548 0 tdc0.w_dly_sig\[67\]
rlabel metal1 4646 5712 4646 5712 0 tdc0.w_dly_sig\[68\]
rlabel metal1 5336 6086 5336 6086 0 tdc0.w_dly_sig\[69\]
rlabel metal1 14214 11628 14214 11628 0 tdc0.w_dly_sig\[6\]
rlabel metal1 4043 5066 4043 5066 0 tdc0.w_dly_sig\[70\]
rlabel metal1 2438 8432 2438 8432 0 tdc0.w_dly_sig\[71\]
rlabel metal1 2438 7990 2438 7990 0 tdc0.w_dly_sig\[72\]
rlabel metal1 1426 11215 1426 11215 0 tdc0.w_dly_sig\[73\]
rlabel metal1 1748 8058 1748 8058 0 tdc0.w_dly_sig\[74\]
rlabel metal2 1334 11832 1334 11832 0 tdc0.w_dly_sig\[75\]
rlabel metal1 1242 8330 1242 8330 0 tdc0.w_dly_sig\[76\]
rlabel metal1 1334 5712 1334 5712 0 tdc0.w_dly_sig\[77\]
rlabel metal1 1518 9146 1518 9146 0 tdc0.w_dly_sig\[78\]
rlabel metal1 1640 4726 1640 4726 0 tdc0.w_dly_sig\[79\]
rlabel metal1 14490 11186 14490 11186 0 tdc0.w_dly_sig\[7\]
rlabel via1 1973 5066 1973 5066 0 tdc0.w_dly_sig\[80\]
rlabel metal1 1748 2550 1748 2550 0 tdc0.w_dly_sig\[81\]
rlabel metal1 1748 2618 1748 2618 0 tdc0.w_dly_sig\[82\]
rlabel metal2 1518 1632 1518 1632 0 tdc0.w_dly_sig\[83\]
rlabel metal1 2806 2550 2806 2550 0 tdc0.w_dly_sig\[84\]
rlabel metal1 3450 2550 3450 2550 0 tdc0.w_dly_sig\[85\]
rlabel metal2 3542 2176 3542 2176 0 tdc0.w_dly_sig\[86\]
rlabel metal1 4232 2618 4232 2618 0 tdc0.w_dly_sig\[87\]
rlabel metal1 5244 2550 5244 2550 0 tdc0.w_dly_sig\[88\]
rlabel metal1 5658 2550 5658 2550 0 tdc0.w_dly_sig\[89\]
rlabel metal1 13294 11730 13294 11730 0 tdc0.w_dly_sig\[8\]
rlabel metal1 5934 2482 5934 2482 0 tdc0.w_dly_sig\[90\]
rlabel metal1 6716 2958 6716 2958 0 tdc0.w_dly_sig\[91\]
rlabel via1 7217 1394 7217 1394 0 tdc0.w_dly_sig\[92\]
rlabel metal1 8372 2482 8372 2482 0 tdc0.w_dly_sig\[93\]
rlabel metal1 8234 1938 8234 1938 0 tdc0.w_dly_sig\[94\]
rlabel metal1 9430 1394 9430 1394 0 tdc0.w_dly_sig\[95\]
rlabel metal1 9138 1802 9138 1802 0 tdc0.w_dly_sig\[96\]
rlabel metal1 11730 2482 11730 2482 0 tdc0.w_dly_sig\[97\]
rlabel metal1 11408 1394 11408 1394 0 tdc0.w_dly_sig\[98\]
rlabel via1 12737 2482 12737 2482 0 tdc0.w_dly_sig\[99\]
rlabel metal1 14858 7276 14858 7276 0 tdc0.w_dly_sig\[9\]
rlabel metal1 18262 13362 18262 13362 0 tdc0.w_dly_sig_n\[0\]
rlabel metal1 14168 1870 14168 1870 0 tdc0.w_dly_sig_n\[100\]
rlabel metal2 13938 1360 13938 1360 0 tdc0.w_dly_sig_n\[101\]
rlabel metal1 14490 1836 14490 1836 0 tdc0.w_dly_sig_n\[102\]
rlabel metal1 15686 1360 15686 1360 0 tdc0.w_dly_sig_n\[103\]
rlabel metal1 16100 1394 16100 1394 0 tdc0.w_dly_sig_n\[104\]
rlabel metal1 16238 2482 16238 2482 0 tdc0.w_dly_sig_n\[105\]
rlabel metal1 16698 2618 16698 2618 0 tdc0.w_dly_sig_n\[106\]
rlabel viali 15594 3569 15594 3569 0 tdc0.w_dly_sig_n\[107\]
rlabel metal2 15778 3264 15778 3264 0 tdc0.w_dly_sig_n\[108\]
rlabel metal1 16330 3434 16330 3434 0 tdc0.w_dly_sig_n\[109\]
rlabel metal1 13800 13362 13800 13362 0 tdc0.w_dly_sig_n\[10\]
rlabel metal1 16974 4080 16974 4080 0 tdc0.w_dly_sig_n\[110\]
rlabel metal1 17250 2618 17250 2618 0 tdc0.w_dly_sig_n\[111\]
rlabel metal1 17296 3978 17296 3978 0 tdc0.w_dly_sig_n\[112\]
rlabel metal1 18308 4114 18308 4114 0 tdc0.w_dly_sig_n\[113\]
rlabel metal1 17848 3978 17848 3978 0 tdc0.w_dly_sig_n\[114\]
rlabel metal1 17710 5780 17710 5780 0 tdc0.w_dly_sig_n\[115\]
rlabel metal1 17848 5882 17848 5882 0 tdc0.w_dly_sig_n\[116\]
rlabel metal1 18354 8432 18354 8432 0 tdc0.w_dly_sig_n\[117\]
rlabel metal1 18768 8262 18768 8262 0 tdc0.w_dly_sig_n\[118\]
rlabel metal1 18538 11628 18538 11628 0 tdc0.w_dly_sig_n\[119\]
rlabel metal1 13202 13294 13202 13294 0 tdc0.w_dly_sig_n\[11\]
rlabel metal1 18860 13838 18860 13838 0 tdc0.w_dly_sig_n\[120\]
rlabel metal2 18446 12308 18446 12308 0 tdc0.w_dly_sig_n\[121\]
rlabel metal1 18722 15572 18722 15572 0 tdc0.w_dly_sig_n\[122\]
rlabel metal1 18170 15538 18170 15538 0 tdc0.w_dly_sig_n\[123\]
rlabel metal1 17756 16014 17756 16014 0 tdc0.w_dly_sig_n\[124\]
rlabel metal1 17756 15878 17756 15878 0 tdc0.w_dly_sig_n\[125\]
rlabel metal1 16698 17034 16698 17034 0 tdc0.w_dly_sig_n\[126\]
rlabel metal1 18032 16422 18032 16422 0 tdc0.w_dly_sig_n\[127\]
rlabel via1 16790 17306 16790 17306 0 tdc0.w_dly_sig_n\[128\]
rlabel metal1 13064 14042 13064 14042 0 tdc0.w_dly_sig_n\[12\]
rlabel metal1 13248 14926 13248 14926 0 tdc0.w_dly_sig_n\[13\]
rlabel metal1 12788 15606 12788 15606 0 tdc0.w_dly_sig_n\[14\]
rlabel metal1 11868 15878 11868 15878 0 tdc0.w_dly_sig_n\[15\]
rlabel metal1 11822 17136 11822 17136 0 tdc0.w_dly_sig_n\[16\]
rlabel metal1 11592 17578 11592 17578 0 tdc0.w_dly_sig_n\[17\]
rlabel metal1 11822 18224 11822 18224 0 tdc0.w_dly_sig_n\[18\]
rlabel metal1 12742 18156 12742 18156 0 tdc0.w_dly_sig_n\[19\]
rlabel metal2 15134 11849 15134 11849 0 tdc0.w_dly_sig_n\[1\]
rlabel metal1 12052 18802 12052 18802 0 tdc0.w_dly_sig_n\[20\]
rlabel metal1 13248 18054 13248 18054 0 tdc0.w_dly_sig_n\[21\]
rlabel metal1 13156 18598 13156 18598 0 tdc0.w_dly_sig_n\[22\]
rlabel metal1 13984 17306 13984 17306 0 tdc0.w_dly_sig_n\[23\]
rlabel metal1 14168 17578 14168 17578 0 tdc0.w_dly_sig_n\[24\]
rlabel metal1 14674 17102 14674 17102 0 tdc0.w_dly_sig_n\[25\]
rlabel metal1 14260 16626 14260 16626 0 tdc0.w_dly_sig_n\[26\]
rlabel metal1 14766 16422 14766 16422 0 tdc0.w_dly_sig_n\[27\]
rlabel metal1 14076 16218 14076 16218 0 tdc0.w_dly_sig_n\[28\]
rlabel metal1 12880 15334 12880 15334 0 tdc0.w_dly_sig_n\[29\]
rlabel metal1 16560 11662 16560 11662 0 tdc0.w_dly_sig_n\[2\]
rlabel metal2 9430 15028 9430 15028 0 tdc0.w_dly_sig_n\[30\]
rlabel metal1 11408 14586 11408 14586 0 tdc0.w_dly_sig_n\[31\]
rlabel metal1 9016 14790 9016 14790 0 tdc0.w_dly_sig_n\[32\]
rlabel metal1 8464 14858 8464 14858 0 tdc0.w_dly_sig_n\[33\]
rlabel metal2 7866 14484 7866 14484 0 tdc0.w_dly_sig_n\[34\]
rlabel metal1 6532 14926 6532 14926 0 tdc0.w_dly_sig_n\[35\]
rlabel metal2 7406 15334 7406 15334 0 tdc0.w_dly_sig_n\[36\]
rlabel metal1 6026 15470 6026 15470 0 tdc0.w_dly_sig_n\[37\]
rlabel metal1 6716 15402 6716 15402 0 tdc0.w_dly_sig_n\[38\]
rlabel metal1 5612 16218 5612 16218 0 tdc0.w_dly_sig_n\[39\]
rlabel metal1 16054 11696 16054 11696 0 tdc0.w_dly_sig_n\[3\]
rlabel metal1 5658 16592 5658 16592 0 tdc0.w_dly_sig_n\[40\]
rlabel metal1 4324 16626 4324 16626 0 tdc0.w_dly_sig_n\[41\]
rlabel metal1 4002 16762 4002 16762 0 tdc0.w_dly_sig_n\[42\]
rlabel metal1 3542 16626 3542 16626 0 tdc0.w_dly_sig_n\[43\]
rlabel metal1 2392 16762 2392 16762 0 tdc0.w_dly_sig_n\[44\]
rlabel metal1 2668 16626 2668 16626 0 tdc0.w_dly_sig_n\[45\]
rlabel metal1 1840 17306 1840 17306 0 tdc0.w_dly_sig_n\[46\]
rlabel metal1 1518 16626 1518 16626 0 tdc0.w_dly_sig_n\[47\]
rlabel metal1 1886 15980 1886 15980 0 tdc0.w_dly_sig_n\[48\]
rlabel metal1 2254 15538 2254 15538 0 tdc0.w_dly_sig_n\[49\]
rlabel metal1 15502 11730 15502 11730 0 tdc0.w_dly_sig_n\[4\]
rlabel metal1 2254 15402 2254 15402 0 tdc0.w_dly_sig_n\[50\]
rlabel metal1 2622 13974 2622 13974 0 tdc0.w_dly_sig_n\[51\]
rlabel metal1 1932 14042 1932 14042 0 tdc0.w_dly_sig_n\[52\]
rlabel metal1 2530 12818 2530 12818 0 tdc0.w_dly_sig_n\[53\]
rlabel metal1 3358 12716 3358 12716 0 tdc0.w_dly_sig_n\[54\]
rlabel metal1 4048 12274 4048 12274 0 tdc0.w_dly_sig_n\[55\]
rlabel metal1 3680 12614 3680 12614 0 tdc0.w_dly_sig_n\[56\]
rlabel metal1 4692 12138 4692 12138 0 tdc0.w_dly_sig_n\[57\]
rlabel metal2 4738 11832 4738 11832 0 tdc0.w_dly_sig_n\[58\]
rlabel metal1 5290 11594 5290 11594 0 tdc0.w_dly_sig_n\[59\]
rlabel metal1 15824 11594 15824 11594 0 tdc0.w_dly_sig_n\[5\]
rlabel metal1 5290 10982 5290 10982 0 tdc0.w_dly_sig_n\[60\]
rlabel metal1 5612 10438 5612 10438 0 tdc0.w_dly_sig_n\[61\]
rlabel metal1 5750 9894 5750 9894 0 tdc0.w_dly_sig_n\[62\]
rlabel via1 4830 9486 4830 9486 0 tdc0.w_dly_sig_n\[63\]
rlabel metal1 5750 8874 5750 8874 0 tdc0.w_dly_sig_n\[64\]
rlabel metal1 4968 8262 4968 8262 0 tdc0.w_dly_sig_n\[65\]
rlabel metal1 4968 7718 4968 7718 0 tdc0.w_dly_sig_n\[66\]
rlabel metal1 3956 7446 3956 7446 0 tdc0.w_dly_sig_n\[67\]
rlabel metal1 3818 6630 3818 6630 0 tdc0.w_dly_sig_n\[68\]
rlabel metal1 3128 6630 3128 6630 0 tdc0.w_dly_sig_n\[69\]
rlabel metal1 14766 11662 14766 11662 0 tdc0.w_dly_sig_n\[6\]
rlabel metal1 2530 7276 2530 7276 0 tdc0.w_dly_sig_n\[70\]
rlabel metal2 2162 7650 2162 7650 0 tdc0.w_dly_sig_n\[71\]
rlabel metal1 2116 7922 2116 7922 0 tdc0.w_dly_sig_n\[72\]
rlabel via1 1610 7922 1610 7922 0 tdc0.w_dly_sig_n\[73\]
rlabel metal2 1242 8160 1242 8160 0 tdc0.w_dly_sig_n\[74\]
rlabel metal2 1058 7956 1058 7956 0 tdc0.w_dly_sig_n\[75\]
rlabel metal1 874 6426 874 6426 0 tdc0.w_dly_sig_n\[76\]
rlabel metal1 1380 5882 1380 5882 0 tdc0.w_dly_sig_n\[77\]
rlabel metal1 1564 4794 1564 4794 0 tdc0.w_dly_sig_n\[78\]
rlabel metal1 1472 3978 1472 3978 0 tdc0.w_dly_sig_n\[79\]
rlabel metal1 14030 11696 14030 11696 0 tdc0.w_dly_sig_n\[7\]
rlabel metal1 1748 2482 1748 2482 0 tdc0.w_dly_sig_n\[80\]
rlabel metal1 2162 2482 2162 2482 0 tdc0.w_dly_sig_n\[81\]
rlabel metal1 1380 2074 1380 2074 0 tdc0.w_dly_sig_n\[82\]
rlabel metal1 2070 1904 2070 1904 0 tdc0.w_dly_sig_n\[83\]
rlabel metal1 2622 1836 2622 1836 0 tdc0.w_dly_sig_n\[84\]
rlabel metal2 3634 1632 3634 1632 0 tdc0.w_dly_sig_n\[85\]
rlabel metal1 3358 1836 3358 1836 0 tdc0.w_dly_sig_n\[86\]
rlabel metal2 5060 1394 5060 1394 0 tdc0.w_dly_sig_n\[87\]
rlabel metal1 5198 2448 5198 2448 0 tdc0.w_dly_sig_n\[88\]
rlabel metal1 5428 1530 5428 1530 0 tdc0.w_dly_sig_n\[89\]
rlabel metal2 14306 12546 14306 12546 0 tdc0.w_dly_sig_n\[8\]
rlabel metal1 6578 1394 6578 1394 0 tdc0.w_dly_sig_n\[90\]
rlabel metal1 7498 1904 7498 1904 0 tdc0.w_dly_sig_n\[91\]
rlabel metal1 7774 1904 7774 1904 0 tdc0.w_dly_sig_n\[92\]
rlabel metal2 8234 2176 8234 2176 0 tdc0.w_dly_sig_n\[93\]
rlabel metal1 8004 1802 8004 1802 0 tdc0.w_dly_sig_n\[94\]
rlabel metal1 9568 1462 9568 1462 0 tdc0.w_dly_sig_n\[95\]
rlabel metal2 10442 1632 10442 1632 0 tdc0.w_dly_sig_n\[96\]
rlabel metal2 11362 2176 11362 2176 0 tdc0.w_dly_sig_n\[97\]
rlabel metal1 12144 1394 12144 1394 0 tdc0.w_dly_sig_n\[98\]
rlabel metal1 12742 1258 12742 1258 0 tdc0.w_dly_sig_n\[99\]
rlabel metal1 13800 12614 13800 12614 0 tdc0.w_dly_sig_n\[9\]
rlabel metal2 19090 11407 19090 11407 0 ui_in[0]
rlabel metal2 12926 534 12926 534 0 ui_in[3]
rlabel metal2 10350 415 10350 415 0 ui_in[4]
rlabel metal2 12282 534 12282 534 0 ui_in[5]
rlabel metal2 11638 415 11638 415 0 ui_in[6]
rlabel via2 17342 12291 17342 12291 0 uo_out[0]
rlabel metal3 13662 8432 13662 8432 0 uo_out[1]
rlabel metal1 16514 12954 16514 12954 0 uo_out[2]
rlabel metal1 17296 10030 17296 10030 0 uo_out[3]
rlabel via2 15962 8925 15962 8925 0 uo_out[4]
rlabel metal1 12788 11118 12788 11118 0 uo_out[5]
rlabel metal1 13708 9146 13708 9146 0 uo_out[6]
rlabel metal2 11684 17340 11684 17340 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
