* PEX produced on Sun Mar 17 01:30:16 PM CET 2024 using /foss/tools/osic-multitool/iic-pex.sh with m=1 and s=1
* NGSPICE file created from tt_um_hpretl_tt06_tdc_v1.ext - technology: sky130A

.subckt tt_um_hpretl_tt06_tdc_v1 clk ena rst_n ui_in[1] ui_in[2] ui_in[5] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[1] uio_oe[2] uio_oe[5] uio_oe[7] uio_out[0] uio_out[3] uio_out[7] uo_out[1]
+ uo_out[2] uo_out[3] uo_out[5] uo_out[6] ui_in[0] ui_in[4] ui_in[6] uio_out[2] uio_out[5]
+ uio_oe[4] uio_oe[0] uo_out[0] uo_out[4] uio_out[4] ui_in[3] uio_out[1] uio_out[6]
+ uo_out[7] uio_oe[6] uio_oe[3] VPWR VGND
X0 a_23315_17833# a_23179_17673# a_22895_17687# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 _051_ a_20359_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2 tdc0.w_dly_sig[61] tdc0.w_dly_sig_n[60] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_25529_2045# a_25191_1831# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5 VPWR tdc0.w_dly_sig_n[177] tdc0.w_dly_sig[179] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 clknet_4_0_0_clk a_6476_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 VPWR _022_ a_13997_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_22261_17833# a_21714_17577# a_21914_17732# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X9 a_11046_5309# a_10607_4943# a_10961_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10 VGND tdc0.w_dly_sig[92] tdc0.w_dly_sig_n[93] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 tdc0.w_dly_sig_n[78] tdc0.w_dly_sig[78] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_19855_7895# _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X13 VGND a_10351_9813# a_10309_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_23053_14557# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X16 VGND a_22971_957# a_23139_859# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_13809_17461# a_13643_17461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR _054_ a_20945_13675# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_21718_5487# a_21279_5493# a_21633_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 VGND tdc0.w_dly_sig[81] tdc0.w_dly_sig_n[82] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VPWR a_9263_14013# a_9431_13915# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X22 tdc0.w_dly_sig[123] tdc0.w_dly_sig_n[121] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 tdc0.o_result[74] a_13019_11739# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR a_8454_7637# a_8381_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X27 a_16210_9839# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X29 a_23457_8207# _010_ a_23385_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 a_10221_14735# a_10055_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X31 a_15236_6575# _031_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X33 _013_ a_15530_6077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X34 VPWR tdc0.w_dly_sig[17] a_29099_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X35 a_13035_5487# a_12171_5493# a_12778_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X36 a_13866_9545# _178_ a_13552_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X37 tdc0.w_dly_sig_n[48] tdc0.w_dly_sig[47] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 a_29541_12559# a_29375_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X40 tdc0.w_dly_sig[13] tdc0.w_dly_sig_n[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X42 tdc0.w_dly_sig_n[75] tdc0.w_dly_sig[75] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X43 VPWR a_11260_5461# clknet_4_2_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X44 VPWR a_11766_18517# a_11693_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X45 VPWR a_12134_15253# a_12061_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X46 net2 a_15575_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X47 a_22178_17277# a_21739_16911# a_22093_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X48 tdc0.w_dly_sig_n[17] tdc0.w_dly_sig[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X49 VGND tdc0.w_dly_sig[13] tdc0.w_dly_sig_n[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X51 _054_ a_17139_8759# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X52 VPWR clknet_4_2_0_clk a_13551_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X53 VPWR a_13955_2223# a_14123_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X54 a_11237_9295# tdc0.w_dly_sig[74] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X55 a_19255_12335# _190_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X56 tdc0.w_dly_sig[184] tdc0.w_dly_sig_n[183] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X57 tdc0.w_dly_sig_n[62] tdc0.w_dly_sig[62] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X58 VGND _058_ a_22445_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X59 tdc0.o_result[165] a_12651_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X60 a_23999_4917# a_24290_5217# a_24241_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X61 VGND a_24490_4917# a_24419_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X62 VPWR tdc0.w_dly_sig_n[60] tdc0.w_dly_sig[62] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X63 a_21886_5461# a_21718_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X64 a_16373_13647# _001_ a_16301_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X65 a_19433_12809# _205_ a_19337_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 VPWR a_20881_11721# uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X67 a_25138_3855# a_24823_4007# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X68 tdc0.o_result[81] a_10903_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X71 VPWR net3 a_15203_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X72 tdc0.w_dly_sig_n[103] tdc0.w_dly_sig[103] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X73 a_13551_11721# _085_ a_13633_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X74 tdc0.w_dly_sig_n[149] tdc0.w_dly_sig[148] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X75 VGND tdc0.w_dly_sig_n[84] tdc0.w_dly_sig[86] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X76 tdc0.o_result[86] a_14675_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X77 VPWR tdc0.w_dly_sig[170] tdc0.w_dly_sig_n[170] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X78 a_30343_11471# a_30123_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X79 tdc0.o_result[68] a_20563_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X80 tdc0.w_dly_sig_n[72] tdc0.w_dly_sig[72] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X81 VGND tdc0.w_dly_sig[2] tdc0.w_dly_sig_n[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X82 tdc0.w_dly_sig[14] tdc0.w_dly_sig_n[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X83 a_17894_8751# _096_ a_17814_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X84 VPWR tdc0.w_dly_sig[101] tdc0.w_dly_sig_n[102] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X85 VGND clknet_4_1_0_clk a_2143_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X86 tdc0.w_dly_sig_n[119] tdc0.w_dly_sig[118] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X87 tdc0.w_dly_sig[193] tdc0.w_dly_sig_n[192] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X88 VGND tdc0.o_result[49] a_24593_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X89 a_29173_4943# a_29007_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X90 VGND _157_ a_12999_8867# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X91 VPWR tdc0.o_result[191] a_20756_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X93 VGND tdc0.w_dly_sig[165] tdc0.w_dly_sig_n[166] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X94 a_11582_7637# a_11414_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X95 VPWR tdc0.w_dly_sig[31] tdc0.w_dly_sig_n[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X96 VGND tdc0.w_dly_sig_n[80] tdc0.w_dly_sig[82] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X97 VPWR tdc0.w_dly_sig_n[133] tdc0.w_dly_sig[135] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X98 VGND tdc0.w_dly_sig_n[43] tdc0.w_dly_sig[45] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X99 a_17481_8457# _101_ a_17409_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X100 a_23189_12335# tdc0.o_result[61] a_22751_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X101 a_12249_9839# tdc0.w_dly_sig[76] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X102 a_29987_11445# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X103 VPWR net1 tdc0.w_dly_sig_n[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X104 a_7734_4399# a_7461_4405# a_7649_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X105 VGND clknet_4_12_0_clk a_22107_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X106 VPWR tdc0.w_dly_sig[181] tdc0.w_dly_sig_n[181] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X107 VGND clknet_4_0_0_clk a_5639_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X108 VGND _155_ a_13722_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X109 a_24915_8983# _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X110 clknet_0_clk a_16210_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X112 a_12521_11837# a_11987_11471# a_12426_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X114 VPWR a_7591_14165# a_7507_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X115 VGND tdc0.w_dly_sig[18] tdc0.w_dly_sig_n[18] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X116 clknet_4_8_0_clk a_21104_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X118 tdc0.w_dly_sig[4] tdc0.w_dly_sig_n[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X119 clknet_4_7_0_clk a_11812_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X120 VPWR a_5199_15253# a_5115_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X121 VPWR tdc0.w_dly_sig_n[120] tdc0.w_dly_sig[122] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X122 VPWR a_6855_13077# a_6771_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X123 a_17665_10927# _094_ a_17415_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X124 tdc0.w_dly_sig[191] tdc0.w_dly_sig_n[189] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X125 tdc0.w_dly_sig_n[76] tdc0.w_dly_sig[75] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X126 a_23634_7637# a_23466_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X127 a_14250_18517# a_14082_18543# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X128 a_23903_2919# a_23999_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X129 a_16451_11265# _034_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X130 a_29998_7663# a_29559_7669# a_29913_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X131 a_27675_12381# a_27455_12393# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X132 a_7553_12021# a_7387_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X133 a_28227_2767# a_28007_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X134 a_27179_3855# a_27043_3829# a_26759_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X136 tdc0.w_dly_sig[154] tdc0.w_dly_sig_n[152] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X137 VPWR a_10506_7119# clknet_4_3_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X139 a_8381_7663# a_7847_7669# a_8286_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X140 a_6998_14191# a_6559_14197# a_6913_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X142 VGND tdc0.w_dly_sig[17] tdc0.w_dly_sig_n[18] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X143 a_14082_18543# a_13809_18549# a_13997_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X144 a_26483_16885# a_26767_16885# a_26702_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X146 tdc0.w_dly_sig_n[172] tdc0.w_dly_sig[171] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X147 VPWR tdc0.w_dly_sig[69] tdc0.w_dly_sig_n[69] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X149 tdc0.w_dly_sig[37] tdc0.w_dly_sig_n[35] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X150 VGND a_7074_15253# a_7032_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X152 a_11172_4943# a_10773_4943# a_11046_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X153 a_14437_8725# _033_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X154 tdc0.o_result[66] a_21759_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X155 VGND a_12254_13103# clknet_4_6_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X156 VGND a_19773_9441# _177_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X157 VGND a_8879_7637# a_8837_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X158 VGND tdc0.w_dly_sig_n[50] tdc0.w_dly_sig[52] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X159 tdc0.o_result[168] a_15595_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X160 VPWR a_10202_3967# a_10129_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X161 VPWR a_8638_3285# a_8565_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X162 tdc0.w_dly_sig[1] tdc0.w_dly_sig_n[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X163 a_21844_5865# a_21445_5493# a_21718_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X164 VPWR clknet_4_13_0_clk a_16587_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X165 VPWR _007_ a_13275_7776# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X166 a_28818_13469# a_28503_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X167 VPWR tdc0.w_dly_sig_n[173] tdc0.w_dly_sig[175] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X168 VGND a_19947_4007# _176_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X170 VGND tdc0.w_dly_sig[88] tdc0.w_dly_sig_n[89] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X171 _093_ a_13551_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X172 VPWR tdc0.w_dly_sig_n[171] tdc0.w_dly_sig[173] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X173 VPWR tdc0.w_dly_sig[173] tdc0.w_dly_sig_n[174] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X174 VPWR a_14887_4631# _162_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X175 VPWR net5 a_16739_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X176 tdc0.w_dly_sig[54] tdc0.w_dly_sig_n[53] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X177 a_24469_12015# tdc0.o_result[5] a_23947_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X178 a_25191_1831# a_25287_1653# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X179 VPWR a_21638_8181# a_21567_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X180 VPWR a_17451_14191# a_17619_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X181 a_3226_14191# a_2787_14197# a_3141_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X183 a_7182_7485# a_6909_7119# a_7097_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X184 a_26575_15511# a_26866_15401# a_26817_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X185 tdc0.w_dly_sig[47] tdc0.w_dly_sig_n[46] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X186 a_10129_4221# a_9595_3855# a_10034_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X187 VPWR a_4555_4373# a_4471_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X188 tdc0.w_dly_sig[179] tdc0.w_dly_sig_n[177] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X190 a_22178_17277# a_21905_16911# a_22093_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X191 a_25755_15797# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X192 a_17703_6895# net5 _064_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X193 a_10459_3133# a_9761_2767# a_10202_2879# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X194 tdc0.w_dly_sig[103] tdc0.w_dly_sig_n[101] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X196 tdc0.w_dly_sig[5] tdc0.w_dly_sig_n[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X197 VPWR tdc0.o_result[158] a_14287_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X198 VGND a_14250_18517# a_14208_18921# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X199 a_11655_2045# a_10791_1679# a_11398_1791# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X200 _161_ a_19150_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X201 a_16692_18921# a_16293_18549# a_16566_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X202 a_8565_15823# a_8399_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X203 tdc0.o_result[31] a_22679_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X204 VGND _166_ a_12434_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X205 VPWR a_29895_4617# a_29902_4521# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X206 a_19395_7895# _011_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X207 VPWR tdc0.w_dly_sig_n[38] tdc0.w_dly_sig[40] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X208 VPWR a_23903_4007# _128_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X209 a_6940_16745# a_6541_16373# a_6814_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X211 VPWR clknet_4_14_0_clk a_29375_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X212 a_26203_11623# a_26299_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X213 a_14507_18543# a_13809_18549# a_14250_18517# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X215 VPWR tdc0.w_dly_sig[35] tdc0.w_dly_sig_n[36] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X216 a_27505_9129# a_26958_8873# a_27158_9028# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X217 tdc0.w_dly_sig_n[11] tdc0.w_dly_sig[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X218 VGND tdc0.w_dly_sig_n[182] tdc0.w_dly_sig[183] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X219 a_15101_16911# tdc0.w_dly_sig[89] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X221 tdc0.w_dly_sig_n[67] tdc0.w_dly_sig[66] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X222 VGND a_7699_15101# a_7867_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X224 VPWR a_12594_11583# a_12521_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X225 a_8197_16373# a_8031_16373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X226 a_1849_11471# a_1683_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X227 a_21327_11159# a_21423_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X228 a_16113_2767# tdc0.w_dly_sig[174] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X229 a_29725_14197# a_29559_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X230 VPWR clknet_0_clk a_6550_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X232 tdc0.w_dly_sig[53] tdc0.w_dly_sig_n[52] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X233 VGND a_16762_15797# a_16691_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X234 net6 a_18151_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X235 VGND a_15333_4737# _039_ VGND sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X236 VPWR a_27503_5705# a_27510_5609# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X237 a_1738_7231# a_1570_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X238 VPWR a_9263_9661# a_9431_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X239 a_22849_3855# _056_ a_22777_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X240 VPWR tdc0.w_dly_sig_n[27] tdc0.w_dly_sig[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X241 a_8872_17833# a_8473_17461# a_8746_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X242 a_15170_2197# a_15002_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X243 tdc0.w_dly_sig_n[19] tdc0.w_dly_sig[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X244 VPWR tdc0.w_dly_sig_n[25] tdc0.w_dly_sig[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X245 VGND clknet_4_1_0_clk a_4167_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X246 tdc0.w_dly_sig[151] tdc0.w_dly_sig_n[149] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X248 a_23999_4917# a_24283_4917# a_24218_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X249 a_9758_9839# a_9319_9845# a_9673_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X250 tdc0.w_dly_sig[91] tdc0.w_dly_sig_n[89] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X251 VGND tdc0.w_dly_sig_n[70] tdc0.w_dly_sig[72] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X252 a_10018_2197# a_9850_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X253 a_13257_2229# a_13091_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X254 a_16635_4007# tdc0.o_result[173] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X256 VPWR clknet_4_0_0_clk a_5639_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X257 VGND a_9834_4373# a_9792_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X258 VGND a_25410_3829# a_25339_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X259 VGND tdc0.w_dly_sig_n[55] tdc0.w_dly_sig[56] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X260 VPWR tdc0.w_dly_sig_n[65] tdc0.w_dly_sig[66] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X261 VPWR _010_ a_19395_6807# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X262 a_18590_2223# a_18317_2229# a_18505_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X263 a_20102_9545# _176_ a_20022_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X264 VPWR tdc0.w_dly_sig_n[172] tdc0.w_dly_sig[174] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X265 a_18003_18365# a_17139_17999# a_17746_18111# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X266 VGND tdc0.w_dly_sig[80] tdc0.w_dly_sig_n[80] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X267 tdc0.w_dly_sig_n[190] tdc0.w_dly_sig[189] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X268 a_7399_6031# a_7270_6305# a_6979_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X269 a_28078_2741# a_27878_3041# a_28227_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X270 a_8565_3311# a_8031_3317# a_8470_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X271 a_5989_4405# a_5823_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X272 a_25707_1679# a_25571_1653# a_25287_1653# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X273 a_2589_7663# tdc0.w_dly_sig[116] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X274 VGND a_16555_15797# a_16562_16097# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X275 a_13797_13647# _001_ a_13725_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X277 a_16350_8751# tdc0.o_result[67] a_16193_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X278 a_17673_18365# a_17139_17999# a_17578_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X279 a_28841_12015# a_28503_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X280 VGND clknet_4_9_0_clk a_21279_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X281 a_11923_6397# a_11141_6031# a_11839_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X282 a_10402_18365# a_10129_17999# a_10317_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X283 VGND a_11214_5055# a_11172_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X284 VGND a_6883_6183# tdc0.o_result[136] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X285 _063_ a_16587_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X287 tdc0.w_dly_sig_n[152] tdc0.w_dly_sig[151] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X288 tdc0.w_dly_sig[102] tdc0.w_dly_sig_n[101] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X289 tdc0.w_dly_sig_n[43] tdc0.w_dly_sig[42] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X290 a_18237_11721# _145_ a_18141_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X291 tdc0.w_dly_sig[156] tdc0.w_dly_sig_n[154] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X292 tdc0.w_dly_sig[133] tdc0.w_dly_sig_n[131] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X294 tdc0.w_dly_sig[82] tdc0.w_dly_sig_n[81] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X295 tdc0.w_dly_sig[80] tdc0.w_dly_sig_n[79] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X296 tdc0.w_dly_sig_n[37] tdc0.w_dly_sig[36] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X297 a_15737_12335# tdc0.o_result[142] a_15299_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X298 VPWR a_22615_4007# _163_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X299 a_17875_3855# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X300 tdc0.w_dly_sig_n[60] tdc0.w_dly_sig[60] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X301 VGND tdc0.w_dly_sig[39] tdc0.w_dly_sig_n[39] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X302 clknet_4_10_0_clk a_25428_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X303 VPWR a_13019_16091# a_12935_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X304 tdc0.w_dly_sig_n[112] tdc0.w_dly_sig[111] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X305 a_19586_18517# a_19418_18543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X307 tdc0.w_dly_sig_n[118] tdc0.w_dly_sig[117] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X308 VGND clknet_4_7_0_clk a_14655_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X309 a_28818_12381# a_28503_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X311 VPWR a_13203_5461# a_13119_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X312 a_30194_11204# a_29994_11049# a_30343_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X313 tdc0.w_dly_sig_n[137] tdc0.w_dly_sig[136] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X314 a_14533_7119# _022_ a_14461_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X315 VGND _076_ a_11865_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X317 a_25019_3529# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X318 a_2953_14197# a_2787_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X320 VGND _004_ a_23844_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X321 VGND tdc0.w_dly_sig_n[158] tdc0.w_dly_sig[160] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X322 a_19825_6397# a_19487_6183# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X323 VPWR clknet_0_clk a_25410_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X324 VGND _026_ a_11313_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X325 VPWR net26 a_27505_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X326 VPWR clk a_16210_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X327 VGND a_24653_9545# uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X328 VPWR clknet_4_15_0_clk a_29559_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X329 a_12171_4512# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X330 a_16543_17063# a_16639_16885# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X331 a_25931_9269# a_26222_9569# a_26173_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X333 clknet_4_4_0_clk a_6550_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X334 a_13081_4943# tdc0.o_result[164] a_12999_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X335 tdc0.w_dly_sig_n[141] tdc0.w_dly_sig[140] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X336 tdc0.w_dly_sig[143] tdc0.w_dly_sig_n[142] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X337 VPWR tdc0.w_dly_sig[25] tdc0.w_dly_sig_n[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X338 a_26351_9295# a_26222_9569# a_25931_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X339 VPWR a_26974_16885# a_26903_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X340 VPWR a_19890_13103# clknet_4_13_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X341 VPWR tdc0.w_dly_sig_n[23] tdc0.w_dly_sig[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X342 VPWR tdc0.w_dly_sig[21] tdc0.w_dly_sig_n[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X343 VPWR _012_ a_15575_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X344 VPWR tdc0.w_dly_sig[119] tdc0.w_dly_sig_n[120] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X345 a_19557_3677# _056_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X346 _075_ a_14182_10159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X347 a_21787_2455# a_21883_2455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X348 VGND a_14250_17429# a_14208_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X349 a_26309_15823# a_25762_16097# a_25962_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X350 VPWR a_26203_11623# tdc0.o_result[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X352 VGND a_6430_4373# a_6388_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X353 VGND tdc0.w_dly_sig[25] a_23825_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X354 a_8929_2601# a_7939_2229# a_8803_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X355 a_25962_12533# a_25762_12833# a_26111_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X356 VPWR a_23662_11204# a_23591_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X357 VPWR tdc0.w_dly_sig[13] tdc0.w_dly_sig_n[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X358 tdc0.w_dly_sig_n[87] tdc0.w_dly_sig[86] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X359 tdc0.w_dly_sig[21] tdc0.w_dly_sig_n[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X360 a_12448_7663# tdc0.o_result[115] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X361 a_14741_9545# _084_ a_14645_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X362 tdc0.o_result[92] a_15595_18267# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X363 a_17567_9447# _018_ a_17741_9323# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X364 VGND tdc0.w_dly_sig_n[20] tdc0.w_dly_sig[22] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X365 VPWR tdc0.w_dly_sig_n[52] tdc0.w_dly_sig[54] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X366 VGND tdc0.w_dly_sig[19] tdc0.w_dly_sig_n[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X367 tdc0.w_dly_sig[192] tdc0.w_dly_sig_n[190] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X368 a_11260_5461# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X369 VGND tdc0.w_dly_sig[67] tdc0.w_dly_sig_n[67] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X370 a_7090_10749# a_6817_10383# a_7005_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X371 tdc0.w_dly_sig_n[34] tdc0.w_dly_sig[33] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X372 VPWR _026_ a_11435_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X373 tdc0.w_dly_sig_n[83] tdc0.w_dly_sig[82] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X374 a_9834_4373# a_9666_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X375 tdc0.w_dly_sig_n[65] tdc0.w_dly_sig[64] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X376 VGND a_23386_17732# a_23315_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X378 VPWR a_7902_4373# a_7829_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X379 a_4774_15253# a_4606_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X380 VGND clknet_4_5_0_clk a_6467_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X382 a_22633_4917# tdc0.o_result[180] a_22886_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X383 a_5031_15279# a_4333_15285# a_4774_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X384 a_21879_12711# a_21975_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X385 tdc0.w_dly_sig[126] tdc0.w_dly_sig_n[125] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X386 a_5123_12015# a_4425_12021# a_4866_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X387 VGND tdc0.w_dly_sig_n[3] tdc0.w_dly_sig[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X388 VPWR a_11679_8983# _027_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X389 VGND tdc0.w_dly_sig[5] tdc0.w_dly_sig_n[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X391 a_13273_13423# _039_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X394 VGND a_6855_13077# a_6813_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X395 _012_ a_19807_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X396 a_22086_4399# a_21813_4405# a_22001_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X397 VPWR tdc0.w_dly_sig[48] tdc0.w_dly_sig_n[49] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X398 VPWR a_18489_9839# uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X399 a_19211_7271# a_19307_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X400 a_16733_4917# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.229 ps=1.75 w=0.42 l=0.15
X401 VPWR tdc0.w_dly_sig[14] tdc0.w_dly_sig_n[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X402 a_7829_4399# a_7295_4405# a_7734_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X404 a_28425_2767# a_27871_2741# a_28078_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X405 VPWR a_17159_859# a_17075_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X406 VPWR a_14255_6835# _035_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X407 VPWR a_17746_18111# a_17673_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X408 uo_out[2] a_17937_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X409 tdc0.o_result[94] a_10995_18267# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X410 a_20966_1791# a_20798_2045# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X411 VGND _020_ a_15012_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X412 tdc0.w_dly_sig[84] tdc0.w_dly_sig_n[83] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X413 _102_ a_15391_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X414 a_18785_14735# tdc0.o_result[121] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X415 VGND tdc0.w_dly_sig[177] tdc0.w_dly_sig_n[177] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X416 a_23300_5807# tdc0.o_result[183] a_23110_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X417 VPWR a_7074_15253# a_7001_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X418 VGND tdc0.w_dly_sig_n[159] tdc0.w_dly_sig[160] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X419 a_16025_9545# _113_ a_15943_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X420 VPWR tdc0.w_dly_sig_n[91] tdc0.w_dly_sig[93] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X421 tdc0.w_dly_sig_n[100] tdc0.w_dly_sig[99] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X422 a_20499_5719# _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X424 VGND a_16205_10901# _085_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X425 VGND a_22852_7093# clknet_4_9_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X426 tdc0.w_dly_sig[77] tdc0.w_dly_sig_n[76] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X427 a_23598_9839# _127_ a_23518_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X428 a_7258_10495# a_7090_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X429 VPWR a_22530_15253# a_22457_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X430 VGND a_21104_6005# clknet_4_8_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X431 VGND tdc0.w_dly_sig_n[27] tdc0.w_dly_sig[28] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X432 VPWR a_21313_13441# _004_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X433 a_18703_11471# tdc0.o_result[4] a_19225_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X434 VPWR tdc0.w_dly_sig[129] tdc0.w_dly_sig_n[129] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X435 VGND a_26939_10071# tdc0.o_result[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X436 a_29274_16644# a_29074_16489# a_29423_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X437 tdc0.o_result[179] a_23139_859# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X438 VGND a_9263_9661# a_9431_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X439 VPWR a_10275_2223# a_10443_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X440 a_10275_2223# a_9577_2229# a_10018_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X441 a_19583_6005# a_19867_6005# a_19802_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X443 a_25402_14013# a_25155_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X444 a_5859_16189# a_4995_15823# a_5602_15935# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X445 VGND a_5602_15935# a_5560_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X446 VPWR a_1922_10901# a_1849_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X448 a_22143_5487# a_21279_5493# a_21886_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X449 a_13622_16367# a_13349_16373# a_13537_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X450 VGND a_3302_15253# a_3260_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X451 VPWR _054_ a_23855_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X452 VGND tdc0.w_dly_sig_n[167] tdc0.w_dly_sig[168] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X453 a_24919_3829# a_25203_3829# a_25138_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X454 a_26951_8969# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X455 VPWR a_7350_7231# a_7277_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X456 a_19982_9071# tdc0.o_result[137] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X457 VPWR tdc0.o_result[36] a_23240_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X458 VPWR tdc0.w_dly_sig[157] tdc0.w_dly_sig_n[158] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X459 a_2217_12925# a_1683_12559# a_2122_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X460 VPWR tdc0.w_dly_sig[160] tdc0.w_dly_sig_n[161] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X461 VGND a_27319_12233# a_27326_12137# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X462 tdc0.w_dly_sig[114] tdc0.w_dly_sig_n[113] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X463 VGND a_7994_11989# a_7952_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X464 clknet_0_clk a_16210_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X465 a_21665_17455# a_21327_17687# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X466 VGND a_12283_3035# a_12241_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X467 VPWR net2 a_16495_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X468 a_23179_17673# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X469 a_2631_11837# a_1849_11471# a_2547_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X470 a_14533_6031# _060_ a_14461_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X471 a_9899_7485# a_9117_7119# a_9815_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X472 tdc0.w_dly_sig_n[125] tdc0.w_dly_sig[125] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X474 tdc0.o_result[137] a_12007_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X475 a_4061_16911# tdc0.w_dly_sig[101] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X476 VGND clknet_0_clk a_11812_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X477 clknet_4_12_0_clk a_21380_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X478 VPWR tdc0.w_dly_sig[115] tdc0.w_dly_sig_n[116] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X480 VPWR a_11823_1947# a_11739_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X481 a_15657_13647# tdc0.o_result[111] a_15575_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X482 VPWR tdc0.w_dly_sig[137] a_7817_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X483 VGND tdc0.w_dly_sig[112] tdc0.w_dly_sig_n[112] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X484 VPWR tdc0.w_dly_sig[182] tdc0.w_dly_sig_n[182] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X485 VPWR tdc0.w_dly_sig_n[160] tdc0.w_dly_sig[162] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X486 a_26939_10071# a_27035_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X487 VPWR _047_ a_13633_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X488 a_23124_4943# _031_ a_22633_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X490 tdc0.w_dly_sig[10] tdc0.w_dly_sig_n[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X491 clknet_4_5_0_clk a_7378_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X492 a_12341_11471# tdc0.w_dly_sig[75] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X493 VPWR a_14983_7093# _007_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X494 tdc0.o_result[155] a_4923_3035# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X495 VGND _022_ a_16373_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X496 VGND a_9723_8751# a_9891_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X497 a_30239_12925# a_29541_12559# a_29982_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X498 VPWR _043_ a_12999_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X499 VGND tdc0.w_dly_sig[186] tdc0.w_dly_sig_n[186] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X501 VPWR clknet_4_13_0_clk a_19347_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X502 VPWR tdc0.w_dly_sig[78] tdc0.w_dly_sig_n[79] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X504 tdc0.w_dly_sig[157] tdc0.w_dly_sig_n[155] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X505 VGND tdc0.w_dly_sig[178] tdc0.w_dly_sig_n[179] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X506 a_12153_15823# a_11987_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X507 tdc0.w_dly_sig[190] tdc0.w_dly_sig_n[188] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X508 a_12153_14735# a_11987_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X509 a_18130_591# a_17953_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X510 tdc0.o_result[79] a_8051_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X511 a_4755_3133# a_4057_2767# a_4498_2879# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X512 a_24837_18921# a_24283_18761# a_24490_18820# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X513 a_26571_8359# a_26667_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X514 VPWR tdc0.w_dly_sig_n[17] tdc0.w_dly_sig[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X515 VPWR a_26215_9269# a_26222_9569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X516 tdc0.w_dly_sig_n[113] tdc0.w_dly_sig[112] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X517 _003_ a_18703_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X518 VPWR _055_ a_18785_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X519 a_27215_15645# a_26995_15657# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X520 VPWR a_20395_14191# a_20563_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X521 VPWR tdc0.w_dly_sig[192] tdc0.w_dly_sig_n[192] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X522 a_19970_14191# a_19531_14197# a_19885_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X523 VGND tdc0.w_dly_sig[59] tdc0.w_dly_sig_n[59] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X524 VGND a_10478_12671# a_10436_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X525 tdc0.w_dly_sig[105] tdc0.w_dly_sig_n[104] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X526 VPWR a_3175_6549# a_3091_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X528 tdc0.o_result[30] a_23507_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X529 a_11605_2767# tdc0.w_dly_sig[168] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X530 VGND tdc0.w_dly_sig[1] tdc0.w_dly_sig_n[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X531 a_22303_2601# a_22174_2345# a_21883_2455# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X532 VGND a_24639_3543# tdc0.o_result[186] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X533 a_21591_15101# a_20893_14735# a_21334_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X534 a_5077_10633# tdc0.o_result[150] a_4995_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X535 a_25573_13647# a_25019_13621# a_25226_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X536 VGND a_26387_17063# tdc0.o_result[50] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X537 _174_ a_15299_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X538 VGND _007_ a_15419_4737# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X539 a_9263_16189# a_8399_15823# a_9006_15935# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X540 VGND a_9006_15935# a_8964_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X541 tdc0.w_dly_sig[88] tdc0.w_dly_sig_n[87] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X542 VPWR a_21327_3543# _082_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X543 VGND a_24059_7637# a_24017_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X544 a_19097_3677# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X545 a_22277_2767# tdc0.w_dly_sig[185] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X546 VPWR tdc0.w_dly_sig[65] tdc0.w_dly_sig_n[66] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X547 a_6813_13481# a_5823_13109# a_6687_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X548 tdc0.w_dly_sig_n[161] tdc0.w_dly_sig[160] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X549 VGND _073_ a_14182_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X550 VGND tdc0.w_dly_sig_n[98] tdc0.w_dly_sig[100] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X551 a_15059_10927# a_14361_10933# a_14802_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X552 VPWR a_21104_6005# clknet_4_8_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X554 VGND tdc0.w_dly_sig_n[153] tdc0.w_dly_sig[155] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X555 tdc0.w_dly_sig[110] tdc0.w_dly_sig_n[109] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X556 a_27518_7663# a_27271_8041# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X557 a_22914_8751# a_22475_8757# a_22829_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X558 VGND tdc0.w_dly_sig[6] tdc0.w_dly_sig_n[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X559 VGND tdc0.w_dly_sig_n[184] tdc0.w_dly_sig[185] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X560 a_27087_9129# a_26958_8873# a_26667_8983# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X561 VPWR tdc0.w_dly_sig[169] tdc0.w_dly_sig_n[169] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X562 a_9581_4399# tdc0.w_dly_sig[142] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X564 tdc0.w_dly_sig_n[90] tdc0.w_dly_sig[90] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X565 a_10405_14013# a_9871_13647# a_10310_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X566 a_27455_12393# a_27326_12137# a_27035_12247# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X567 tdc0.w_dly_sig_n[101] tdc0.w_dly_sig[100] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X568 VPWR tdc0.w_dly_sig_n[45] tdc0.w_dly_sig[47] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X569 a_25226_13621# a_25019_13621# a_25402_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X570 VGND tdc0.w_dly_sig[127] tdc0.w_dly_sig_n[127] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X573 tdc0.w_dly_sig_n[30] tdc0.w_dly_sig[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X574 a_4606_15279# a_4333_15285# a_4521_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X576 a_4882_8573# a_4443_8207# a_4797_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X577 VGND tdc0.w_dly_sig_n[16] tdc0.w_dly_sig[17] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X578 VGND a_8711_7663# a_8879_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X579 VGND tdc0.w_dly_sig[113] tdc0.w_dly_sig_n[113] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X580 a_19145_18549# a_18979_18549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X581 VGND tdc0.w_dly_sig[106] tdc0.w_dly_sig_n[106] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X582 VPWR a_6476_7637# clknet_4_1_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X583 tdc0.w_dly_sig[116] tdc0.w_dly_sig_n[114] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X584 a_24419_15823# a_24290_16097# a_23999_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X585 a_10478_13759# a_10310_14013# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X586 VGND _053_ a_16587_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X587 VPWR a_29423_5719# tdc0.o_result[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X588 VPWR tdc0.w_dly_sig_n[28] tdc0.w_dly_sig[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X589 tdc0.o_result[159] a_7867_3035# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X590 VPWR _026_ a_16350_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X591 VGND clknet_4_5_0_clk a_6559_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X592 a_25155_13647# a_25019_13621# a_24735_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X593 a_10919_15101# a_10221_14735# a_10662_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X594 VPWR _012_ a_23351_14423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X596 tdc0.w_dly_sig_n[82] tdc0.w_dly_sig[81] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X598 VPWR a_12851_11837# a_13019_11739# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X599 VGND tdc0.w_dly_sig[150] tdc0.w_dly_sig_n[151] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X600 VPWR tdc0.w_dly_sig[122] tdc0.w_dly_sig_n[122] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X601 a_17685_12809# _072_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X602 a_15002_2223# a_14563_2229# a_14917_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X603 a_29607_11159# a_29703_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X605 VPWR tdc0.w_dly_sig_n[106] tdc0.w_dly_sig[108] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X606 a_12254_13103# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X607 VPWR tdc0.w_dly_sig_n[99] tdc0.w_dly_sig[101] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X608 a_14717_10383# _058_ a_14645_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X609 a_10735_12925# a_9871_12559# a_10478_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X610 a_3229_15279# a_2695_15285# a_3134_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X611 a_20003_6031# a_19867_6005# a_19583_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X612 VGND a_18059_7663# _001_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X613 tdc0.w_dly_sig[101] tdc0.w_dly_sig_n[100] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X614 a_20395_14191# a_19531_14197# a_20138_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X615 VGND clknet_4_14_0_clk a_29375_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X616 a_16301_6575# net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X617 _195_ a_14931_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X618 a_14250_15253# a_14082_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X620 a_12426_16189# a_11987_15823# a_12341_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X622 VGND _190_ a_19255_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X623 a_25191_1831# a_25287_1653# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X625 tdc0.w_dly_sig_n[177] tdc0.w_dly_sig[176] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X626 VGND _031_ a_24580_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X627 a_20065_14191# a_19531_14197# a_19970_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X628 a_17695_6575# net6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X629 VPWR tdc0.w_dly_sig[20] a_27137_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X630 uo_out[0] a_20881_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X631 VPWR tdc0.w_dly_sig[86] tdc0.w_dly_sig_n[86] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X632 tdc0.w_dly_sig_n[46] tdc0.w_dly_sig[45] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X633 a_20039_13799# _003_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X635 VPWR tdc0.w_dly_sig[118] tdc0.w_dly_sig_n[118] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X636 tdc0.w_dly_sig_n[22] tdc0.w_dly_sig[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X637 a_23193_7669# a_23027_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X638 VPWR tdc0.w_dly_sig[26] tdc0.w_dly_sig_n[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X639 tdc0.w_dly_sig[86] tdc0.w_dly_sig_n[84] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X642 VPWR a_26859_15497# a_26866_15401# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X643 tdc0.w_dly_sig_n[102] tdc0.w_dly_sig[101] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X644 VPWR tdc0.w_dly_sig[10] tdc0.w_dly_sig_n[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X645 VPWR a_11582_14165# a_11509_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X646 VGND tdc0.w_dly_sig_n[153] tdc0.w_dly_sig[154] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X647 tdc0.w_dly_sig_n[78] tdc0.w_dly_sig[77] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X648 a_11414_6575# a_10975_6581# a_11329_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X649 tdc0.w_dly_sig[39] tdc0.w_dly_sig_n[38] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X651 a_15101_7637# _011_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X652 a_12885_10217# a_11895_9845# a_12759_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X653 VGND a_10827_18365# a_10995_18267# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X654 a_12153_14735# a_11987_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X655 a_16566_957# a_16293_591# a_16481_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X656 clknet_0_clk a_16210_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X657 VGND a_3394_14165# a_3352_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X658 a_15013_3855# tdc0.o_result[143] a_14931_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X659 tdc0.w_dly_sig_n[138] tdc0.w_dly_sig[138] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X660 VGND a_25111_11445# a_25118_11745# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X661 a_6177_4399# tdc0.w_dly_sig[152] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X662 tdc0.o_result[147] a_4279_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X663 tdc0.o_result[149] a_2163_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X664 clknet_4_8_0_clk a_21104_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X665 VPWR tdc0.w_dly_sig[90] tdc0.w_dly_sig_n[91] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X666 tdc0.w_dly_sig[82] tdc0.w_dly_sig_n[80] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X667 a_4698_12015# a_4259_12021# a_4613_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X668 VGND tdc0.w_dly_sig_n[102] tdc0.w_dly_sig[103] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X669 a_15370_12925# a_14931_12559# a_15285_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X670 a_12772_9545# _087_ a_12670_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X671 a_11509_6397# a_10975_6031# a_11414_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X672 VPWR _011_ a_20039_13799# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X674 VPWR a_22254_4373# a_22181_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X675 a_10310_12925# a_10037_12559# a_10225_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X676 VPWR tdc0.w_dly_sig_n[164] tdc0.w_dly_sig[165] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X677 tdc0.w_dly_sig[56] tdc0.w_dly_sig_n[54] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X679 a_9021_3689# a_8031_3317# a_8895_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X680 VPWR _112_ a_17967_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X681 VPWR a_9006_15935# a_8933_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X682 a_6587_4221# a_5805_3855# a_6503_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X683 tdc0.w_dly_sig_n[74] tdc0.w_dly_sig[74] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X684 VPWR a_10478_13759# a_10405_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X685 tdc0.w_dly_sig_n[136] tdc0.w_dly_sig[136] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X686 VGND tdc0.w_dly_sig_n[123] tdc0.w_dly_sig[125] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X687 VGND tdc0.w_dly_sig[8] tdc0.w_dly_sig_n[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X688 a_20074_11204# a_19874_11049# a_20223_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X689 a_5307_6397# a_4609_6031# a_5050_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X690 tdc0.w_dly_sig_n[98] tdc0.w_dly_sig[97] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X691 a_29939_5865# a_29810_5609# a_29519_5719# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X692 VGND a_14805_6549# _080_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X693 VGND tdc0.w_dly_sig_n[118] tdc0.w_dly_sig[120] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X694 _050_ a_16916_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X695 a_25046_7119# a_24731_7271# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X696 VPWR a_15227_10901# a_15143_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X697 a_16481_591# tdc0.w_dly_sig[171] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X698 VGND a_16219_1143# net3 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X699 a_11853_9089# _026_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X702 VGND a_15595_18267# a_15553_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X703 VGND clknet_4_4_0_clk a_7387_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X704 a_19289_13441# _011_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X705 VGND clknet_4_0_0_clk a_5823_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X706 VGND tdc0.w_dly_sig[114] tdc0.w_dly_sig_n[114] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X707 VPWR tdc0.w_dly_sig[48] a_27413_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X709 a_5802_3133# a_5529_2767# a_5717_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X710 a_19867_11145# clknet_4_13_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X711 VGND a_18003_18365# a_18171_18267# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X713 VGND _063_ a_20359_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X714 VGND a_8895_3311# a_9063_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X715 VGND _034_ a_13797_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X716 VPWR a_17619_2197# a_17535_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X717 a_1485_7119# tdc0.w_dly_sig[114] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X718 a_5008_8207# a_4609_8207# a_4882_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X719 VGND a_25962_15797# a_25891_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X720 a_25046_11471# a_24731_11623# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X721 VGND net3 _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X722 a_11325_18549# a_11159_18549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X723 VGND tdc0.w_dly_sig[93] tdc0.w_dly_sig_n[94] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X724 a_30124_3689# a_29725_3317# a_29998_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X726 a_24659_12015# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X727 a_15262_15935# a_15094_16189# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X728 a_20053_3677# _038_ a_19981_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X729 a_30370_11837# a_30123_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X730 a_15170_2197# a_15002_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X731 VPWR tdc0.w_dly_sig[2] tdc0.w_dly_sig_n[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X732 VGND a_9926_9813# a_9884_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X734 VPWR a_22311_5461# a_22227_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X735 VPWR tdc0.o_result[54] a_20204_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X736 VPWR tdc0.w_dly_sig_n[66] tdc0.w_dly_sig[67] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X737 tdc0.o_result[93] a_12191_18517# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X738 a_24419_2767# a_24283_2741# a_23999_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X739 a_21975_12533# a_22259_12533# a_22194_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X740 tdc0.w_dly_sig_n[169] tdc0.w_dly_sig[169] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X741 VGND _168_ a_12434_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X742 VPWR tdc0.w_dly_sig_n[74] tdc0.w_dly_sig[76] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X743 tdc0.w_dly_sig_n[18] tdc0.w_dly_sig[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X744 VGND tdc0.w_dly_sig_n[141] tdc0.w_dly_sig[142] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X745 VGND _120_ a_14274_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X746 tdc0.w_dly_sig_n[8] tdc0.w_dly_sig[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X747 _009_ net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X748 tdc0.o_result[93] a_12191_18517# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X749 VPWR tdc0.w_dly_sig[80] tdc0.w_dly_sig_n[81] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X750 VPWR a_25502_8181# a_25431_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X751 a_15564_8207# tdc0.o_result[50] a_14989_8353# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X752 a_29909_12925# a_29375_12559# a_29814_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X753 a_10528_11471# a_10129_11471# a_10402_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X754 tdc0.w_dly_sig_n[58] tdc0.w_dly_sig[57] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X755 VGND a_21380_14165# clknet_4_12_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X756 a_19826_5193# _136_ a_19746_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X757 VGND a_4739_7637# a_4697_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X758 tdc0.w_dly_sig_n[101] tdc0.w_dly_sig[101] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X759 a_18046_4719# tdc0.o_result[148] a_17965_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X760 a_17415_11247# tdc0.o_result[2] a_17937_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X761 a_7645_11721# tdc0.o_result[114] a_7561_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X762 VPWR a_20138_14165# a_20065_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X763 VGND a_25019_3529# a_25026_3433# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X764 a_11609_3855# tdc0.o_result[159] a_11527_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X765 VPWR tdc0.w_dly_sig_n[37] tdc0.w_dly_sig[38] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X766 tdc0.w_dly_sig[174] tdc0.w_dly_sig_n[173] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X767 VPWR _039_ a_13552_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X768 VGND tdc0.w_dly_sig_n[175] tdc0.w_dly_sig[177] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X769 VPWR tdc0.w_dly_sig_n[11] tdc0.w_dly_sig[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X770 VGND a_25755_15797# a_25762_16097# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X771 VGND a_18758_2197# a_18716_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X772 a_27277_12015# a_26939_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X773 a_7442_14847# a_7274_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X774 a_6369_12335# tdc0.o_result[119] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X775 a_29725_7669# a_29559_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X776 tdc0.o_result[130] a_9431_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X778 VGND tdc0.w_dly_sig_n[17] tdc0.w_dly_sig[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X779 _166_ a_12539_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X780 VGND a_24363_4007# _108_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X781 a_17685_12809# _055_ a_17887_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X784 a_22273_13109# a_22107_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X785 a_23339_8751# a_22641_8757# a_23082_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X786 a_22898_10495# a_22730_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X787 a_11046_5309# a_10773_4943# a_10961_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X788 VPWR clknet_4_1_0_clk a_8859_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X789 a_16481_18543# tdc0.w_dly_sig[57] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X790 a_22181_4399# a_21647_4405# a_22086_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X791 VPWR _117_ a_15365_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X792 a_11540_6953# a_11141_6581# a_11414_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X793 VPWR tdc0.w_dly_sig_n[49] tdc0.w_dly_sig[50] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X794 VGND tdc0.w_dly_sig_n[76] tdc0.w_dly_sig[78] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R0 VGND uio_out[1] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X795 VPWR a_17467_10357# _034_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X796 VGND _183_ a_20417_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X798 tdc0.w_dly_sig[155] tdc0.w_dly_sig_n[154] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X799 a_23733_17833# a_23179_17673# a_23386_17732# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X800 a_3141_3311# tdc0.w_dly_sig[155] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X803 tdc0.o_result[81] a_10903_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X804 a_20614_3133# a_20341_2767# a_20529_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X806 clknet_4_1_0_clk a_6476_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X808 VGND a_21327_11159# tdc0.o_result[34] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X810 tdc0.w_dly_sig[141] tdc0.w_dly_sig_n[140] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X811 VPWR tdc0.w_dly_sig_n[19] tdc0.w_dly_sig[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X812 a_17695_6575# _001_ _064_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X813 a_10551_17277# a_9687_16911# a_10294_17023# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X814 VGND a_10294_17023# a_10252_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X815 a_7461_4405# a_7295_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X816 a_24666_16189# a_24419_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X818 VGND tdc0.w_dly_sig_n[107] tdc0.w_dly_sig[109] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X819 tdc0.o_result[133] a_5199_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X820 tdc0.o_result[61] a_22771_17179# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X821 VPWR tdc0.w_dly_sig_n[108] tdc0.w_dly_sig[109] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X822 _017_ a_19289_13441# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X823 a_11839_7663# a_11141_7669# a_11582_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X824 tdc0.w_dly_sig_n[110] tdc0.w_dly_sig[110] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X825 a_12864_7663# _123_ a_12762_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X826 a_12107_18543# a_11325_18549# a_12023_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X827 tdc0.w_dly_sig[72] tdc0.w_dly_sig_n[70] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X828 VGND clknet_4_1_0_clk a_4259_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X829 tdc0.w_dly_sig_n[108] tdc0.w_dly_sig[108] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X830 VGND tdc0.w_dly_sig_n[67] tdc0.w_dly_sig[68] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X831 tdc0.o_result[155] a_4923_3035# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X832 a_16495_12559# _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X833 a_7258_10495# a_7090_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X834 VGND tdc0.w_dly_sig_n[122] tdc0.w_dly_sig[123] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X835 tdc0.w_dly_sig_n[166] tdc0.w_dly_sig[165] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X836 tdc0.w_dly_sig[66] tdc0.w_dly_sig_n[65] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X837 tdc0.w_dly_sig[172] tdc0.w_dly_sig_n[170] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X838 a_27689_8041# a_27142_7785# a_27342_7940# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X839 tdc0.w_dly_sig[104] tdc0.w_dly_sig_n[103] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X840 _058_ a_18703_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X841 VGND tdc0.w_dly_sig[139] tdc0.w_dly_sig_n[140] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X842 tdc0.o_result[67] a_15687_16091# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X843 a_2037_12559# tdc0.w_dly_sig[108] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X844 VPWR a_1811_6397# a_1979_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X845 tdc0.w_dly_sig[60] tdc0.w_dly_sig_n[58] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X846 a_3873_7669# a_3707_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X847 tdc0.w_dly_sig_n[121] tdc0.w_dly_sig[120] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X849 VPWR tdc0.w_dly_sig[54] tdc0.w_dly_sig_n[55] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X850 VGND tdc0.w_dly_sig_n[2] tdc0.w_dly_sig[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X851 VPWR tdc0.w_dly_sig_n[166] tdc0.w_dly_sig[168] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X853 tdc0.o_result[77] a_11455_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X854 tdc0.w_dly_sig_n[49] tdc0.w_dly_sig[48] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X855 a_30194_11445# a_29987_11445# a_30370_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X856 VGND a_16645_11989# _062_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X858 tdc0.w_dly_sig[165] tdc0.w_dly_sig_n[164] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X859 VGND a_4387_4399# a_4555_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X860 VGND a_17937_10927# uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X861 VGND tdc0.w_dly_sig_n[73] tdc0.w_dly_sig[74] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X862 a_23339_8751# a_22475_8757# a_23082_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X863 tdc0.o_result[44] a_30591_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X864 VGND tdc0.w_dly_sig[22] tdc0.w_dly_sig_n[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X865 VGND a_19807_12559# _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X866 a_6687_4399# a_5823_4405# a_6430_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X867 _013_ net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X869 tdc0.w_dly_sig_n[99] tdc0.w_dly_sig[99] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X870 a_24283_15797# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X871 a_30123_11471# a_29987_11445# a_29703_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X872 VGND a_23075_4007# _052_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X873 VGND clknet_4_10_0_clk a_29651_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X874 a_17026_14191# a_16587_14197# a_16941_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X875 VPWR tdc0.w_dly_sig[179] tdc0.w_dly_sig_n[179] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X876 VPWR tdc0.w_dly_sig[50] tdc0.w_dly_sig_n[50] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X877 VPWR tdc0.w_dly_sig[162] tdc0.w_dly_sig_n[163] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X878 tdc0.w_dly_sig_n[121] tdc0.w_dly_sig[121] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X879 VGND tdc0.w_dly_sig_n[165] tdc0.w_dly_sig[167] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X880 a_21104_6005# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X881 a_14983_7093# _006_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X882 VPWR a_11839_6575# a_12007_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X883 tdc0.w_dly_sig_n[128] tdc0.w_dly_sig[128] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X884 a_20172_9071# tdc0.o_result[9] a_19982_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X885 a_4977_6397# a_4443_6031# a_4882_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X886 a_11831_9661# a_11049_9295# a_11747_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X887 a_26479_15511# a_26575_15511# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X888 VGND _068_ a_20981_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X889 a_6906_15279# a_6467_15285# a_6821_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X890 _119_ a_13735_14304# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X891 a_26886_9117# a_26571_8983# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X892 _130_ a_15115_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X893 uo_out[7] a_20697_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X894 VGND net2 _000_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X895 VGND clknet_4_5_0_clk a_2787_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X896 a_16869_3855# _038_ a_16797_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X897 a_30711_6794# tdc0.w_dly_sig[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X898 a_12977_11471# a_11987_11471# a_12851_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X899 a_22615_4007# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X900 clknet_4_2_0_clk a_11260_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X902 a_18045_6031# net5 a_17691_6281# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X903 VGND tdc0.w_dly_sig[17] a_29099_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X904 VGND tdc0.w_dly_sig_n[123] tdc0.w_dly_sig[124] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X905 VPWR a_14675_18517# a_14591_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X906 tdc0.w_dly_sig_n[51] tdc0.w_dly_sig[51] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X907 VGND tdc0.w_dly_sig[68] tdc0.w_dly_sig_n[68] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X908 a_15427_2223# a_14729_2229# a_15170_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X909 VPWR a_15427_2223# a_15595_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X910 VGND _165_ a_12999_8867# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X911 tdc0.w_dly_sig_n[62] tdc0.w_dly_sig[61] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X912 a_8293_2223# tdc0.w_dly_sig[162] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X913 VGND a_16623_3133# a_16791_3035# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X914 VPWR tdc0.w_dly_sig[120] tdc0.w_dly_sig_n[120] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X915 clknet_4_7_0_clk a_11812_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X916 VGND a_25962_4917# a_25891_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X917 VPWR tdc0.w_dly_sig_n[108] tdc0.w_dly_sig[110] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X918 a_6813_5865# a_5823_5493# a_6687_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X919 a_17313_8457# _109_ a_17231_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X920 VGND a_16991_18543# a_17159_18517# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X921 a_20348_9295# tdc0.o_result[54] a_19773_9441# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X922 VGND a_25410_13103# clknet_4_15_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X923 tdc0.o_result[159] a_7867_3035# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X924 tdc0.w_dly_sig[168] tdc0.w_dly_sig_n[166] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X925 a_2405_4399# tdc0.w_dly_sig[153] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X926 VPWR a_7378_13103# clknet_4_5_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X928 tdc0.w_dly_sig[148] tdc0.w_dly_sig_n[147] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X929 VGND tdc0.w_dly_sig[95] tdc0.w_dly_sig_n[95] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X930 VGND tdc0.w_dly_sig[141] tdc0.w_dly_sig_n[142] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X932 a_19777_12015# _064_ a_19255_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X933 tdc0.o_result[175] a_19183_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X934 tdc0.w_dly_sig[54] tdc0.w_dly_sig_n[52] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X935 a_25690_12559# a_25375_12711# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X936 VPWR a_27158_8181# a_27087_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X937 _075_ a_14182_10159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X939 a_24490_15797# a_24283_15797# a_24666_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X940 tdc0.o_result[103] a_6027_16091# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X942 a_19970_14191# a_19697_14197# a_19885_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X943 VGND a_22898_10495# a_22856_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X944 VPWR tdc0.w_dly_sig[143] tdc0.w_dly_sig_n[144] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X945 tdc0.w_dly_sig_n[25] tdc0.w_dly_sig[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X946 tdc0.w_dly_sig_n[27] tdc0.w_dly_sig[26] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X947 a_17773_6031# _030_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X950 a_22001_4399# tdc0.w_dly_sig[32] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X951 a_16569_17461# a_16403_17461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X952 clknet_4_14_0_clk a_26882_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X953 VPWR a_16635_4007# _168_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X954 _110_ a_17231_8457# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X955 a_15186_17277# a_14747_16911# a_15101_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X957 a_24419_15823# a_24283_15797# a_23999_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X958 a_27242_15279# a_26995_15657# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X959 tdc0.w_dly_sig[4] tdc0.w_dly_sig_n[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X960 VGND clknet_4_4_0_clk a_6651_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X961 tdc0.w_dly_sig_n[5] tdc0.w_dly_sig[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X963 _191_ a_8491_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X964 VGND tdc0.w_dly_sig_n[152] tdc0.w_dly_sig[153] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X965 a_13633_11721# tdc0.o_result[106] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X966 VPWR a_16210_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X967 VGND a_9171_17455# a_9339_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X969 VPWR tdc0.w_dly_sig_n[151] tdc0.w_dly_sig[153] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R1 VGND uio_out[4] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X970 a_19487_11159# a_19583_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X971 VPWR tdc0.w_dly_sig_n[180] tdc0.w_dly_sig[182] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X972 a_28599_13335# a_28883_13321# a_28818_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X973 tdc0.w_dly_sig_n[34] tdc0.w_dly_sig[34] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X974 a_8243_4399# a_7461_4405# a_8159_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X975 VGND _177_ a_19163_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X977 VPWR tdc0.w_dly_sig_n[72] tdc0.w_dly_sig[73] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X978 a_5050_8319# a_4882_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X980 a_3049_15279# tdc0.w_dly_sig[105] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X981 a_22488_15657# a_22089_15285# a_22362_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X982 VPWR a_5970_2879# a_5897_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X983 VGND _047_ a_13724_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X984 a_2290_13077# a_2122_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X985 _098_ a_14103_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X986 VGND tdc0.w_dly_sig_n[30] tdc0.w_dly_sig[32] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X987 VPWR a_3099_7663# a_3267_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X988 VGND a_8454_7637# a_8412_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X989 VPWR tdc0.w_dly_sig_n[133] tdc0.w_dly_sig[134] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X990 VGND tdc0.w_dly_sig[132] tdc0.w_dly_sig_n[133] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X991 VPWR tdc0.w_dly_sig[36] tdc0.w_dly_sig_n[36] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X992 VGND a_13035_5487# a_13203_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X993 tdc0.w_dly_sig_n[19] tdc0.w_dly_sig[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X994 a_29239_13469# a_29019_13481# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X995 VGND a_13955_2223# a_14123_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X996 VGND _007_ a_13061_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X997 a_29955_5309# a_29173_4943# a_29871_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X998 a_18785_14985# tdc0.o_result[57] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1000 VPWR tdc0.w_dly_sig_n[0] tdc0.w_dly_sig[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1001 VGND ui_in[0] a_30347_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1002 tdc0.w_dly_sig_n[117] tdc0.w_dly_sig[116] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1003 VPWR tdc0.w_dly_sig_n[10] tdc0.w_dly_sig[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1004 VPWR a_18059_7663# _001_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1005 VPWR a_26790_11445# a_26719_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1006 VGND a_12927_9813# a_12885_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1007 tdc0.w_dly_sig[176] tdc0.w_dly_sig_n[174] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1008 VPWR a_18151_1135# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1009 tdc0.w_dly_sig_n[145] tdc0.w_dly_sig[144] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1011 tdc0.w_dly_sig[63] tdc0.w_dly_sig_n[61] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1012 a_16753_14197# a_16587_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1013 a_13997_15279# tdc0.w_dly_sig[87] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1014 tdc0.w_dly_sig[187] tdc0.w_dly_sig_n[186] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1015 VPWR tdc0.o_result[85] a_12999_12128# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1016 VGND a_23903_18775# tdc0.o_result[53] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1017 a_17703_6895# net5 _064_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1018 tdc0.w_dly_sig[47] tdc0.w_dly_sig_n[45] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1019 tdc0.w_dly_sig_n[128] tdc0.w_dly_sig[127] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1020 a_2290_12671# a_2122_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1021 VPWR tdc0.w_dly_sig[76] tdc0.w_dly_sig_n[77] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1022 _193_ a_23110_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X1023 a_12241_1513# a_11251_1141# a_12115_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1024 tdc0.w_dly_sig_n[57] tdc0.w_dly_sig[56] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1025 a_23114_17821# a_22799_17687# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1026 a_15427_2223# a_14563_2229# a_15170_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1027 a_18154_5847# net2 a_18073_5847# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0536 ps=0.675 w=0.42 l=0.15
X1028 _170_ a_12999_8867# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X1029 VPWR tdc0.w_dly_sig[188] tdc0.w_dly_sig_n[188] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1030 VGND _069_ a_20900_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1031 VGND _054_ a_14717_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1033 a_27123_16911# a_26903_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1034 tdc0.w_dly_sig_n[130] tdc0.w_dly_sig[130] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1035 a_4038_11583# a_3870_11837# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1037 _161_ a_19150_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X1038 a_20605_10217# a_20051_10057# a_20258_10116# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1039 a_3505_10933# a_3339_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1040 a_14039_2223# a_13257_2229# a_13955_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1042 a_27689_8041# a_27135_7881# a_27342_7940# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1043 clknet_4_5_0_clk a_7378_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1044 VGND tdc0.w_dly_sig_n[110] tdc0.w_dly_sig[112] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1045 a_2547_11837# a_1683_11471# a_2290_11583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1046 tdc0.o_result[120] a_5935_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1048 VPWR tdc0.w_dly_sig_n[142] tdc0.w_dly_sig[144] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1050 VGND tdc0.w_dly_sig_n[128] tdc0.w_dly_sig[129] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1051 a_9171_17455# a_8307_17461# a_8914_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1052 tdc0.w_dly_sig_n[163] tdc0.w_dly_sig[162] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1053 VPWR a_10995_18267# a_10911_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1054 VGND tdc0.w_dly_sig[156] tdc0.w_dly_sig_n[156] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1056 VGND a_5935_9563# a_5893_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1057 tdc0.o_result[79] a_8051_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1058 a_19777_12015# tdc0.o_result[6] a_19255_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X1059 a_16198_3133# a_15925_2767# a_16113_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1061 a_29729_9839# tdc0.w_dly_sig[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1062 VGND a_19855_8359# _159_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1063 a_18505_2223# tdc0.w_dly_sig[176] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1064 VPWR tdc0.o_result[172] a_17875_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1065 tdc0.o_result[151] a_6855_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1066 VGND tdc0.w_dly_sig[151] tdc0.w_dly_sig_n[152] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1067 VPWR a_11214_5055# a_11141_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1068 a_12325_4765# _026_ a_12253_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1069 a_12061_9845# a_11895_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1070 a_14131_12353# _001_ a_14045_12353# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1071 tdc0.w_dly_sig_n[79] tdc0.w_dly_sig[78] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1072 VPWR clknet_4_7_0_clk a_11987_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1073 VGND tdc0.w_dly_sig_n[11] tdc0.w_dly_sig[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1074 a_18348_16745# a_17949_16373# a_18222_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1076 VPWR tdc0.w_dly_sig_n[155] tdc0.w_dly_sig[157] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1077 VGND tdc0.w_dly_sig[175] tdc0.w_dly_sig_n[175] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1078 VGND clknet_4_6_0_clk a_11987_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1079 a_29913_3311# tdc0.w_dly_sig[191] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1080 VPWR a_20782_2879# a_20709_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1081 _071_ a_20543_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X1082 a_27066_15556# a_26859_15497# a_27242_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1083 a_14839_13897# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X1084 VPWR a_15609_4971# _008_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X1085 a_9807_8751# a_9025_8757# a_9723_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1086 VGND tdc0.w_dly_sig_n[29] tdc0.w_dly_sig[31] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1087 VPWR tdc0.w_dly_sig[51] a_27321_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1088 tdc0.w_dly_sig_n[86] tdc0.w_dly_sig[86] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1089 a_24827_7093# a_25111_7093# a_25046_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1090 VGND tdc0.w_dly_sig[132] tdc0.w_dly_sig_n[132] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1091 VPWR a_11030_8319# a_10957_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1092 a_22971_16189# a_22107_15823# a_22714_15935# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1093 VGND a_22714_15935# a_22672_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1094 tdc0.w_dly_sig_n[21] tdc0.w_dly_sig[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1095 _210_ a_19255_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1096 VPWR a_17231_4399# _043_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1097 tdc0.w_dly_sig[139] tdc0.w_dly_sig_n[137] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1098 a_15328_9839# _004_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1099 VGND a_19777_12015# uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1100 a_30370_10927# a_30123_11305# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1101 VGND a_21523_13799# _068_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1102 a_23390_11293# a_23075_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1103 VPWR a_23323_10651# a_23239_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1105 tdc0.w_dly_sig[136] tdc0.w_dly_sig_n[134] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1106 a_18953_11721# _134_ a_18703_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1107 VPWR tdc0.w_dly_sig_n[135] tdc0.w_dly_sig[137] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1109 tdc0.o_result[117] a_4739_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1110 a_7549_14569# a_6559_14197# a_7423_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1111 VGND tdc0.w_dly_sig[166] tdc0.w_dly_sig_n[167] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1112 VGND a_16739_7895# _021_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1113 tdc0.w_dly_sig_n[2] tdc0.w_dly_sig[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1114 a_27319_10057# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1115 a_15186_17277# a_14913_16911# a_15101_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1116 VGND a_10202_2879# a_10160_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1117 a_17137_3855# _039_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X1118 tdc0.w_dly_sig_n[116] tdc0.w_dly_sig[115] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1119 VPWR tdc0.w_dly_sig_n[48] tdc0.w_dly_sig[49] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1120 VGND tdc0.w_dly_sig[28] tdc0.w_dly_sig_n[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1121 VGND a_19395_3543# _204_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1122 a_22641_16189# a_22107_15823# a_22546_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1123 tdc0.w_dly_sig_n[38] tdc0.w_dly_sig[37] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1125 tdc0.w_dly_sig[10] tdc0.w_dly_sig_n[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1126 tdc0.w_dly_sig[145] tdc0.w_dly_sig_n[144] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1127 VPWR _030_ a_18659_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1128 VGND clknet_4_4_0_clk a_4259_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1129 a_18758_2197# a_18590_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1130 a_25471_4917# a_25755_4917# a_25690_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1131 VPWR tdc0.w_dly_sig[138] tdc0.w_dly_sig_n[138] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1132 a_2122_11837# a_1849_11471# a_2037_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1133 tdc0.w_dly_sig[186] tdc0.w_dly_sig_n[185] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1134 VPWR tdc0.w_dly_sig[89] tdc0.w_dly_sig_n[90] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1135 a_12693_6941# _060_ a_12621_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1136 VPWR _022_ a_14045_12353# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1137 a_24283_4917# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1139 _094_ a_16679_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X1140 VPWR tdc0.o_result[163] a_12539_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1141 a_5123_12015# a_4259_12021# a_4866_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1142 a_13641_6031# _039_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X1143 a_19418_18543# a_19145_18549# a_19333_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1144 a_17559_12711# _111_ a_17887_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1146 VPWR tdc0.w_dly_sig[175] tdc0.w_dly_sig_n[176] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1147 a_18545_9117# _019_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1148 VGND tdc0.w_dly_sig[106] tdc0.w_dly_sig_n[107] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1149 VGND tdc0.w_dly_sig[162] tdc0.w_dly_sig_n[162] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1150 VPWR clknet_4_7_0_clk a_13643_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1151 a_14802_10901# a_14634_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1152 tdc0.o_result[63] a_22955_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1153 VGND a_7378_13103# clknet_4_5_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R2 tt_um_hpretl_tt06_tdc_v1_21.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1154 tdc0.o_result[110] a_2347_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1155 VPWR a_7683_10651# a_7599_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1156 VGND tdc0.w_dly_sig_n[190] tdc0.w_dly_sig[192] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1157 VPWR a_23507_8725# a_23423_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1158 VPWR tdc0.w_dly_sig_n[57] tdc0.w_dly_sig[59] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1159 VPWR a_16734_703# a_16661_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1161 VGND tdc0.w_dly_sig[103] tdc0.w_dly_sig_n[103] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1162 tdc0.w_dly_sig_n[82] tdc0.w_dly_sig[82] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1163 VGND a_4866_11989# a_4824_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1164 a_4330_3133# a_3891_2767# a_4245_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1165 tdc0.o_result[12] a_30039_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1166 a_2731_9839# a_2033_9845# a_2474_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1167 VPWR a_6855_4373# a_6771_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1168 VGND tdc0.w_dly_sig_n[31] tdc0.w_dly_sig[32] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1169 a_21905_16911# a_21739_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1170 tdc0.w_dly_sig[182] tdc0.w_dly_sig_n[180] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1171 a_29239_12381# a_29019_12393# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1172 VGND tdc0.w_dly_sig[117] tdc0.w_dly_sig_n[118] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1173 tdc0.w_dly_sig_n[149] tdc0.w_dly_sig[149] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1174 a_14634_10927# a_14361_10933# a_14549_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1175 a_15115_9545# _121_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1176 a_19567_957# a_18869_591# a_19310_703# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1177 a_16205_10901# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X1178 a_18046_4719# _144_ a_18292_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X1179 VPWR clknet_4_4_0_clk a_1683_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1181 a_4797_8207# tdc0.w_dly_sig[133] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1182 a_15023_10383# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1183 a_10773_4943# a_10607_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1184 a_16573_14735# tdc0.w_dly_sig[70] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1185 tdc0.w_dly_sig_n[154] tdc0.w_dly_sig[154] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1186 VPWR tdc0.w_dly_sig_n[13] tdc0.w_dly_sig[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1187 a_19855_7895# tdc0.o_result[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1188 a_18893_8029# _030_ a_18821_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1189 a_24021_14985# tdc0.o_result[63] a_23937_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1190 VGND tdc0.w_dly_sig_n[77] tdc0.w_dly_sig[78] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1191 tdc0.w_dly_sig_n[122] tdc0.w_dly_sig[122] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1192 VGND a_29607_11159# tdc0.o_result[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1193 VPWR a_25428_7637# clknet_4_10_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1194 a_16691_15823# a_16555_15797# a_16271_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1195 tdc0.w_dly_sig[101] tdc0.w_dly_sig_n[99] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1196 tdc0.w_dly_sig[108] tdc0.w_dly_sig_n[106] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1197 a_10202_3967# a_10034_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1198 a_2290_11583# a_2122_11837# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1199 a_7124_14569# a_6725_14197# a_6998_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1200 VPWR tdc0.w_dly_sig[2] a_26769_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1201 uo_out[5] a_24469_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1202 a_16121_10383# tdc0.o_result[92] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X1203 a_19353_5853# _010_ a_19281_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1204 VGND _174_ a_19255_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1205 a_11141_5309# a_10607_4943# a_11046_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1206 VGND a_30683_6299# a_30641_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1207 VPWR a_29423_6196# net28 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1208 tdc0.w_dly_sig[28] tdc0.w_dly_sig_n[27] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1209 VGND clknet_4_4_0_clk a_1683_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1210 VPWR tdc0.w_dly_sig_n[1] tdc0.w_dly_sig[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1211 tdc0.w_dly_sig[137] tdc0.w_dly_sig_n[135] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1212 VGND tdc0.w_dly_sig[91] tdc0.w_dly_sig_n[91] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1213 a_12621_3677# tdc0.o_result[163] a_12539_3424# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1214 _041_ a_13735_4512# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1217 a_10570_18111# a_10402_18365# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1218 tdc0.w_dly_sig_n[122] tdc0.w_dly_sig[121] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1219 a_16210_9839# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1221 a_18087_18365# a_17305_17999# a_18003_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1222 clknet_4_12_0_clk a_21380_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1223 a_21327_3543# tdc0.o_result[177] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1224 VPWR _011_ a_15023_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1225 a_18046_4719# _143_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X1226 VGND a_18737_6059# _031_ VGND sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X1227 tdc0.w_dly_sig_n[12] tdc0.w_dly_sig[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1228 VPWR ui_in[4] a_16219_1143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1229 a_8753_13647# tdc0.w_dly_sig[125] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1230 a_19089_3133# a_18751_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1231 a_4146_17277# a_3707_16911# a_4061_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1233 tdc0.w_dly_sig_n[171] tdc0.w_dly_sig[170] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1234 _153_ a_13082_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X1235 VGND a_26571_8983# tdc0.o_result[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1236 a_20395_14191# a_19697_14197# a_20138_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1237 a_7826_12015# a_7387_12021# a_7741_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1238 VPWR tdc0.w_dly_sig[85] tdc0.w_dly_sig_n[85] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1239 VGND _023_ a_8745_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1240 tdc0.o_result[89] a_14215_16341# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1241 VPWR a_12254_13103# clknet_4_6_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1242 a_17565_8725# _033_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X1243 VPWR clknet_4_0_0_clk a_7295_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1245 a_30194_11204# a_29987_11145# a_30370_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1247 VPWR _012_ a_19899_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X1248 VPWR tdc0.w_dly_sig_n[53] tdc0.w_dly_sig[55] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1249 a_8573_11247# tdc0.o_result[135] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1250 VGND a_7902_4373# a_7860_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1251 VGND tdc0.w_dly_sig[96] tdc0.w_dly_sig_n[97] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1252 VPWR tdc0.w_dly_sig[50] tdc0.w_dly_sig_n[51] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1253 VPWR clknet_4_6_0_clk a_11987_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1254 VGND tdc0.w_dly_sig_n[130] tdc0.w_dly_sig[131] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1255 tdc0.o_result[60] a_18815_16341# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1256 a_14937_3677# _038_ a_14865_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1257 a_5549_11247# _027_ a_5115_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1258 a_24183_15511# _066_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X1259 a_2263_10927# a_1481_10933# a_2179_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1260 VGND _033_ a_16737_9441# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X1261 tdc0.w_dly_sig_n[91] tdc0.w_dly_sig[90] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1262 VPWR a_22714_15935# a_22641_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1263 tdc0.w_dly_sig[42] tdc0.w_dly_sig_n[40] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1264 VGND tdc0.w_dly_sig_n[142] tdc0.w_dly_sig[143] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1265 tdc0.w_dly_sig[103] tdc0.w_dly_sig_n[102] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1266 a_30123_11305# a_29987_11145# a_29703_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1267 tdc0.w_dly_sig[127] tdc0.w_dly_sig_n[125] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1268 a_6273_12015# _191_ a_6191_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1269 _181_ a_13722_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X1270 a_7274_3133# a_6835_2767# a_7189_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1271 VPWR a_16547_4373# _056_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1272 VGND _055_ a_23189_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X1273 a_20992_4719# tdc0.o_result[46] a_20417_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X1274 VGND a_1811_6397# a_1979_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1275 a_6629_3855# a_5639_3855# a_6503_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1276 a_30423_15279# a_29559_15285# a_30166_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1277 tdc0.w_dly_sig_n[109] tdc0.w_dly_sig[109] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1279 tdc0.w_dly_sig_n[147] tdc0.w_dly_sig[147] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1280 VPWR a_21914_17732# a_21843_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1281 tdc0.o_result[77] a_11455_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1282 VGND tdc0.w_dly_sig[55] a_22261_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1283 VGND tdc0.w_dly_sig[65] a_17109_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1284 VGND _133_ a_15943_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1285 tdc0.w_dly_sig[168] tdc0.w_dly_sig_n[167] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1286 a_22790_5193# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X1287 a_21334_14847# a_21166_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1288 a_26886_8207# a_26571_8359# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1289 VPWR tdc0.w_dly_sig_n[176] tdc0.w_dly_sig[177] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1290 a_21327_3543# tdc0.o_result[177] a_21561_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1291 a_29541_9845# a_29375_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1292 VPWR a_16623_3133# a_16791_3035# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1293 VGND tdc0.w_dly_sig[146] tdc0.w_dly_sig_n[146] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1295 VGND a_19798_7093# a_19727_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1297 tdc0.w_dly_sig_n[189] tdc0.w_dly_sig[188] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1298 tdc0.w_dly_sig_n[92] tdc0.w_dly_sig[91] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1299 a_30093_15279# a_29559_15285# a_29998_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1301 VGND tdc0.w_dly_sig[40] a_25573_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1302 VGND a_4555_4373# a_4513_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1303 a_2221_9839# tdc0.w_dly_sig[113] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1304 VPWR a_9006_9407# a_8933_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1305 VGND tdc0.w_dly_sig_n[131] tdc0.w_dly_sig[132] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1306 tdc0.w_dly_sig[35] tdc0.w_dly_sig_n[33] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1307 tdc0.w_dly_sig_n[100] tdc0.w_dly_sig[100] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1309 a_7825_14735# a_6835_14735# a_7699_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1310 tdc0.w_dly_sig_n[5] tdc0.w_dly_sig[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1311 a_24131_9545# _071_ a_24381_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1312 VPWR _035_ a_14839_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X1313 VGND _003_ a_19375_13441# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1314 tdc0.w_dly_sig_n[160] tdc0.w_dly_sig[159] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1315 a_15134_6575# _078_ a_15054_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X1317 a_15925_2767# a_15759_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1318 a_17218_3855# _104_ a_17464_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X1319 a_22093_16911# tdc0.w_dly_sig[62] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1320 a_7917_11471# tdc0.o_result[98] a_7479_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1321 a_4456_2767# a_4057_2767# a_4330_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1322 VGND tdc0.w_dly_sig[108] tdc0.w_dly_sig_n[109] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1323 VGND a_14045_12353# _072_ VGND sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X1324 VPWR tdc0.w_dly_sig_n[119] tdc0.w_dly_sig[121] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1325 VPWR tdc0.w_dly_sig_n[192] tdc0.w_dly_sig[193] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1327 VGND a_17010_17429# a_16968_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1329 VGND _082_ a_14897_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X1330 VGND tdc0.w_dly_sig[164] tdc0.w_dly_sig_n[165] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1332 VPWR tdc0.w_dly_sig[71] tdc0.w_dly_sig_n[71] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1333 a_8201_7663# tdc0.w_dly_sig[132] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1334 tdc0.w_dly_sig[155] tdc0.w_dly_sig_n[153] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1335 VPWR tdc0.w_dly_sig[53] tdc0.w_dly_sig_n[54] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1336 VGND tdc0.w_dly_sig[47] tdc0.w_dly_sig_n[47] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1338 a_30005_6031# net25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1339 VGND a_11839_6397# a_12007_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1340 tdc0.w_dly_sig_n[46] tdc0.w_dly_sig[46] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1341 tdc0.w_dly_sig[185] tdc0.w_dly_sig_n[183] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1342 a_2674_7663# a_2235_7669# a_2589_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1343 tdc0.w_dly_sig_n[116] tdc0.w_dly_sig[116] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R3 tt_um_hpretl_tt06_tdc_v1_17.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1344 VPWR a_15595_2197# a_15511_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1345 VGND a_2163_7387# a_2121_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1346 VGND a_22799_17687# tdc0.o_result[52] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1347 a_8470_16367# a_8031_16373# a_8385_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1348 a_29998_14191# a_29559_14197# a_29913_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1349 a_29853_4399# a_29515_4631# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1351 a_6909_16367# a_6375_16373# a_6814_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1352 tdc0.w_dly_sig_n[69] tdc0.w_dly_sig[68] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1353 VGND tdc0.w_dly_sig_n[187] tdc0.w_dly_sig[189] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1354 VPWR a_25410_13103# clknet_4_15_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1355 tdc0.w_dly_sig[118] tdc0.w_dly_sig_n[117] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1356 VPWR a_14989_8353# _101_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X1358 tdc0.w_dly_sig[38] tdc0.w_dly_sig_n[37] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1360 a_25375_8983# tdc0.o_result[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1361 a_12249_9839# tdc0.w_dly_sig[76] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1362 VPWR tdc0.w_dly_sig_n[173] tdc0.w_dly_sig[174] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1363 tdc0.w_dly_sig_n[131] tdc0.w_dly_sig[130] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1364 VGND tdc0.w_dly_sig[69] tdc0.w_dly_sig_n[70] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1365 a_23891_7663# a_23193_7669# a_23634_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1366 a_22895_17687# a_23179_17673# a_23114_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1367 tdc0.w_dly_sig[9] tdc0.w_dly_sig_n[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1368 a_10436_13647# a_10037_13647# a_10310_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1369 VPWR a_16366_2879# a_16293_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1371 VGND tdc0.w_dly_sig_n[139] tdc0.w_dly_sig[140] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1372 VPWR a_16645_11989# _062_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X1373 VPWR tdc0.w_dly_sig_n[148] tdc0.w_dly_sig[150] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1374 VPWR a_4463_11739# a_4379_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1376 tdc0.w_dly_sig[177] tdc0.w_dly_sig_n[176] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1377 _004_ a_21313_13441# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X1378 VGND tdc0.w_dly_sig_n[105] tdc0.w_dly_sig[107] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1379 VGND a_17194_14165# a_17152_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1380 a_4146_17277# a_3873_16911# a_4061_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1381 tdc0.o_result[65] a_20379_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1382 VPWR tdc0.w_dly_sig[14] tdc0.w_dly_sig_n[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1383 VGND tdc0.w_dly_sig[155] tdc0.w_dly_sig_n[156] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1384 VGND clknet_4_13_0_clk a_22107_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1386 a_19513_15285# a_19347_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1387 a_4054_4221# a_3781_3855# a_3969_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1388 a_25318_11445# a_25118_11745# a_25467_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1390 tdc0.o_result[65] a_20379_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1391 VGND _040_ a_13889_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1392 VPWR tdc0.w_dly_sig_n[41] tdc0.w_dly_sig[42] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1394 tdc0.w_dly_sig[50] tdc0.w_dly_sig_n[49] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1395 tdc0.w_dly_sig_n[111] tdc0.w_dly_sig[110] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1396 VPWR clknet_4_0_0_clk a_7939_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1397 a_26939_10071# a_27035_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1398 VPWR tdc0.w_dly_sig[58] tdc0.w_dly_sig_n[58] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1399 a_27127_13335# a_27418_13225# a_27369_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1400 _151_ a_17691_14985# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1401 _034_ a_17467_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1403 VPWR tdc0.w_dly_sig_n[107] tdc0.w_dly_sig[108] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1404 _085_ a_16205_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.38 ps=2.76 w=1 l=0.15
X1405 VPWR a_10183_9839# a_10351_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1406 VGND clknet_0_clk a_26882_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1407 a_5066_15101# a_4627_14735# a_4981_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1408 a_25506_1679# a_25191_1831# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1410 a_22633_4917# _031_ a_22790_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1411 a_7400_2767# a_7001_2767# a_7274_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1412 tdc0.w_dly_sig[137] tdc0.w_dly_sig_n[136] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1413 a_22871_3133# a_22089_2767# a_22787_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1414 VGND tdc0.w_dly_sig[60] tdc0.w_dly_sig_n[60] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1415 a_25069_7485# a_24731_7271# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1416 VPWR tdc0.w_dly_sig_n[55] tdc0.w_dly_sig[57] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1417 VPWR a_19119_5719# _078_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1418 VGND tdc0.w_dly_sig[133] tdc0.w_dly_sig_n[133] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1419 VGND tdc0.w_dly_sig_n[182] tdc0.w_dly_sig[184] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1420 a_11517_7119# tdc0.o_result[131] a_11435_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1421 VPWR a_30166_15253# a_30093_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1422 VGND _150_ a_18703_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X1423 VGND _045_ a_13722_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X1424 a_5989_10927# tdc0.o_result[116] a_5905_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1425 VGND a_10275_2223# a_10443_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1426 VGND tdc0.w_dly_sig_n[20] tdc0.w_dly_sig[21] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1427 VPWR a_17691_7119# _010_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1428 tdc0.w_dly_sig[87] tdc0.w_dly_sig_n[86] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1429 VPWR tdc0.w_dly_sig[44] tdc0.w_dly_sig_n[44] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1430 tdc0.w_dly_sig[154] tdc0.w_dly_sig_n[153] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1432 tdc0.o_result[87] a_13019_16091# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1433 VPWR a_16355_7969# a_16179_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1434 a_30423_14191# a_29559_14197# a_30166_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1435 _164_ a_12723_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1436 VPWR tdc0.o_result[72] a_16495_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1437 VGND a_22143_5487# a_22311_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1438 tdc0.w_dly_sig[117] tdc0.w_dly_sig_n[116] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1439 tdc0.w_dly_sig[123] tdc0.w_dly_sig_n[122] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1440 VGND tdc0.w_dly_sig[181] tdc0.w_dly_sig_n[182] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1441 a_17279_16911# a_17059_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1442 VPWR a_2715_13915# a_2631_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1443 VGND a_17159_859# a_17117_591# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1444 tdc0.w_dly_sig_n[24] tdc0.w_dly_sig[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1445 VPWR tdc0.w_dly_sig[25] tdc0.w_dly_sig_n[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1446 a_16916_4373# _042_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1447 tdc0.w_dly_sig_n[150] tdc0.w_dly_sig[149] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1448 a_17691_6281# _000_ a_17773_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1450 VGND a_13203_5461# a_13161_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1451 VGND a_15519_16189# a_15687_16091# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1453 VGND a_29803_5705# a_29810_5609# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1454 a_25755_12533# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1455 a_22167_2441# clknet_4_8_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1456 _008_ a_15609_4971# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X1457 tdc0.w_dly_sig[3] tdc0.w_dly_sig_n[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1458 VGND tdc0.w_dly_sig_n[33] tdc0.w_dly_sig[34] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1461 a_30093_14191# a_29559_14197# a_29998_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1462 VGND _035_ a_14257_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1463 VGND a_4498_2879# a_4456_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1464 tdc0.w_dly_sig[18] tdc0.w_dly_sig_n[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1465 VPWR _007_ a_15609_4971# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1467 VGND a_27250_3829# a_27179_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1468 VGND tdc0.w_dly_sig[49] tdc0.w_dly_sig_n[50] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1469 tdc0.w_dly_sig[34] tdc0.w_dly_sig_n[32] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1470 tdc0.w_dly_sig[74] tdc0.w_dly_sig_n[73] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1471 a_15925_2767# a_15759_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1472 VGND a_14583_3035# a_14541_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1473 a_13354_13423# tdc0.o_result[140] a_13273_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X1474 tdc0.w_dly_sig_n[186] tdc0.w_dly_sig[185] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1475 a_10359_2223# a_9577_2229# a_10275_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1476 VPWR tdc0.w_dly_sig[114] tdc0.w_dly_sig_n[115] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1477 tdc0.w_dly_sig_n[93] tdc0.w_dly_sig[93] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1478 VPWR clknet_4_10_0_clk a_29007_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1479 a_29703_11445# a_29994_11745# a_29945_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1480 a_14868_8751# _020_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1481 a_20295_15279# a_19513_15285# a_20211_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1482 a_2800_8041# a_2401_7669# a_2674_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1483 a_10129_11471# a_9963_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1485 a_12805_6031# tdc0.o_result[149] a_12723_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1486 clknet_4_1_0_clk a_6476_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1487 VGND a_20499_13799# _207_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1488 a_16293_3133# a_15759_2767# a_16198_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1490 VGND _039_ a_15737_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X1491 clknet_4_2_0_clk a_11260_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1492 VGND _127_ a_23269_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X1493 VGND a_7591_14165# a_7549_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1494 VPWR a_27031_13335# tdc0.o_result[40] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1495 a_11690_1135# a_11417_1141# a_11605_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1496 VPWR tdc0.w_dly_sig_n[13] tdc0.w_dly_sig[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1497 VPWR tdc0.o_result[133] a_13275_7776# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1498 tdc0.w_dly_sig[51] tdc0.w_dly_sig_n[49] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1499 VGND tdc0.w_dly_sig[43] tdc0.w_dly_sig_n[44] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1500 _028_ a_8399_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1501 VPWR a_20697_12809# uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1502 VGND _012_ a_17808_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X1503 tdc0.w_dly_sig_n[139] tdc0.w_dly_sig[139] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1504 VGND clknet_4_2_0_clk a_9227_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1505 VGND tdc0.w_dly_sig_n[8] tdc0.w_dly_sig[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1507 a_30166_8725# a_29998_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1508 a_30549_9129# a_29559_8757# a_30423_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1510 VGND _088_ a_12526_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X1511 VGND _065_ a_18140_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1512 tdc0.w_dly_sig_n[32] tdc0.w_dly_sig[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1513 a_17967_10159# _112_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1514 clknet_4_7_0_clk a_11812_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1515 VGND a_7591_3285# a_7549_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1516 VPWR a_2290_13759# a_2217_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1517 VPWR net3 a_17383_5095# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1518 VPWR tdc0.o_result[24] a_17168_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X1519 a_12521_16189# a_11987_15823# a_12426_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1521 VGND a_6476_6549# clknet_4_0_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1522 a_19267_2767# a_19131_2741# a_18847_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1523 VPWR a_30407_12827# a_30323_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1524 tdc0.w_dly_sig_n[99] tdc0.w_dly_sig[98] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1525 VPWR clknet_0_clk a_7378_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1526 tdc0.w_dly_sig_n[120] tdc0.w_dly_sig[120] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1527 a_14173_16745# a_13183_16373# a_14047_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1530 VGND _076_ a_13153_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1531 a_13905_2767# tdc0.w_dly_sig[172] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1532 tdc0.w_dly_sig[110] tdc0.w_dly_sig_n[108] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1533 a_23206_6941# a_22891_6807# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1534 a_2769_7663# a_2235_7669# a_2674_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1535 a_25161_4221# a_24823_4007# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1536 tdc0.w_dly_sig[175] tdc0.w_dly_sig_n[174] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1537 tdc0.w_dly_sig_n[140] tdc0.w_dly_sig[140] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1538 a_7607_7485# a_6909_7119# a_7350_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1539 a_10409_14735# tdc0.w_dly_sig[84] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1540 tdc0.w_dly_sig_n[148] tdc0.w_dly_sig[148] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1541 tdc0.w_dly_sig[24] tdc0.w_dly_sig_n[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1542 VPWR tdc0.w_dly_sig_n[24] tdc0.w_dly_sig[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1543 a_10317_17999# tdc0.w_dly_sig[95] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1544 a_10459_4221# a_9595_3855# a_10202_3967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1545 a_19255_12335# _064_ a_19777_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1546 a_16761_10927# _093_ a_16679_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1547 VPWR tdc0.w_dly_sig[22] tdc0.w_dly_sig_n[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1548 VGND tdc0.w_dly_sig_n[71] tdc0.w_dly_sig[72] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1550 VGND a_5859_16189# a_6027_16091# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1551 tdc0.w_dly_sig_n[105] tdc0.w_dly_sig[104] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1552 tdc0.o_result[174] a_19735_859# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1553 VGND _207_ a_19221_13793# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X1554 VPWR tdc0.w_dly_sig[73] tdc0.w_dly_sig_n[73] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1555 a_26138_5309# a_25891_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1556 VPWR a_16210_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1557 tdc0.w_dly_sig_n[20] tdc0.w_dly_sig[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1558 a_21843_11305# a_21714_11049# a_21423_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1559 VGND a_21104_6005# clknet_4_8_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1560 a_7001_15279# a_6467_15285# a_6906_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1561 a_27043_4617# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1562 a_24915_8983# tdc0.o_result[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1564 a_7649_4399# tdc0.w_dly_sig[144] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1565 a_24186_16341# a_24018_16367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1566 VPWR tdc0.w_dly_sig_n[65] tdc0.w_dly_sig[67] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1567 a_5257_9295# tdc0.w_dly_sig[121] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1568 a_19986_10205# a_19671_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1569 a_3099_7663# a_2401_7669# a_2842_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1570 a_24837_15823# a_24283_15797# a_24490_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1571 a_21147_8181# a_21438_8481# a_21389_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1572 a_20421_11305# a_19874_11049# a_20074_11204# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1573 VPWR tdc0.w_dly_sig[116] tdc0.w_dly_sig_n[116] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1574 VGND tdc0.w_dly_sig[123] tdc0.w_dly_sig_n[124] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1576 a_12999_4943# _024_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1577 a_25537_9117# _012_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1578 a_18679_9839# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1579 a_20945_13675# _003_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1580 a_24293_14735# tdc0.o_result[47] a_23855_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1582 VPWR a_30166_14165# a_30093_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1583 a_20175_12559# _210_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1584 VGND a_19487_11159# tdc0.o_result[32] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1585 tdc0.w_dly_sig[152] tdc0.w_dly_sig_n[151] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1586 a_11711_13216# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1587 a_22346_17023# a_22178_17277# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1588 VPWR tdc0.w_dly_sig_n[162] tdc0.w_dly_sig[163] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1589 tdc0.w_dly_sig[14] tdc0.w_dly_sig_n[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1590 tdc0.w_dly_sig_n[132] tdc0.w_dly_sig[131] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1591 VGND clknet_4_4_0_clk a_1683_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1592 a_22730_10749# a_22457_10383# a_22645_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1593 a_21787_2455# a_21883_2455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1594 a_24131_9295# tdc0.o_result[1] a_24653_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X1595 tdc0.w_dly_sig[73] tdc0.w_dly_sig_n[72] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1596 VPWR tdc0.w_dly_sig_n[134] tdc0.w_dly_sig[136] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1597 a_16635_4007# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X1598 VGND a_10506_7119# clknet_4_3_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1599 VGND a_21638_8181# a_21567_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1600 a_23947_12335# _152_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1601 a_30507_3311# a_29725_3317# a_30423_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1602 VPWR a_11812_13621# clknet_4_7_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1603 a_17026_14191# a_16753_14197# a_16941_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1604 tdc0.w_dly_sig[129] tdc0.w_dly_sig_n[127] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1605 _038_ a_16733_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.176 ps=1.84 w=0.65 l=0.15
X1606 tdc0.w_dly_sig_n[136] tdc0.w_dly_sig[135] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1607 _036_ a_16679_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1608 VPWR clknet_4_4_0_clk a_7019_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1609 a_16857_11247# tdc0.o_result[146] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X1610 VPWR tdc0.o_result[153] a_11251_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1611 a_3781_3855# a_3615_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1612 a_17096_13103# _049_ a_16994_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X1613 VPWR net6 a_16401_6691# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X1614 a_10478_12671# a_10310_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1616 a_6311_3133# a_5529_2767# a_6227_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1617 VPWR a_26422_9269# a_26351_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1618 tdc0.w_dly_sig[62] tdc0.w_dly_sig_n[60] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1619 VPWR _076_ a_11711_13216# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1620 _143_ a_12171_4512# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1621 VPWR a_14250_17429# a_14177_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1622 a_25111_11445# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1624 tdc0.w_dly_sig_n[134] tdc0.w_dly_sig[134] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1625 tdc0.w_dly_sig[24] tdc0.w_dly_sig_n[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1628 VGND clknet_4_13_0_clk a_16587_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1629 VGND a_10735_12925# a_10903_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1630 VGND a_8251_12015# a_8419_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1631 VPWR _030_ a_19579_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1632 VGND a_16210_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1633 tdc0.w_dly_sig[71] tdc0.w_dly_sig_n[70] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1634 a_21707_11145# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1635 VPWR _085_ a_16109_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1636 _156_ a_12999_12128# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1637 tdc0.w_dly_sig_n[17] tdc0.w_dly_sig[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1638 a_23271_6793# clknet_4_9_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1639 tdc0.w_dly_sig_n[103] tdc0.w_dly_sig[102] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1640 a_21071_11721# tdc0.o_result[0] a_20881_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X1642 tdc0.w_dly_sig_n[192] tdc0.w_dly_sig[191] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1643 tdc0.o_result[51] a_24611_16341# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1644 VPWR a_12594_15935# a_12521_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1645 a_20017_4737# _043_ a_19931_4737# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1646 tdc0.w_dly_sig_n[143] tdc0.w_dly_sig[143] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1647 VGND a_5050_6143# a_5008_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1648 a_15943_10383# _020_ a_16121_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X1649 VPWR tdc0.w_dly_sig[105] tdc0.w_dly_sig_n[105] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1650 tdc0.w_dly_sig[121] tdc0.w_dly_sig_n[120] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1651 clknet_4_11_0_clk a_26514_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1653 a_7189_2767# tdc0.w_dly_sig[160] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1655 _139_ a_12723_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1656 tdc0.o_result[51] a_24611_16341# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1657 a_26759_3829# a_27043_3829# a_26978_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1658 VGND a_3175_6549# a_3133_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1659 tdc0.w_dly_sig_n[96] tdc0.w_dly_sig[96] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1660 VGND tdc0.w_dly_sig[97] tdc0.w_dly_sig_n[98] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1661 a_5157_15657# a_4167_15285# a_5031_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1662 a_15293_9545# _125_ a_15197_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1663 a_13866_12809# _198_ a_13552_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X1664 tdc0.w_dly_sig[167] tdc0.w_dly_sig_n[165] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1665 tdc0.w_dly_sig_n[0] net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1666 a_5249_12393# a_4259_12021# a_5123_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1667 VPWR a_8803_2223# a_8971_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1668 VPWR a_30102_4676# a_30031_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1669 VPWR a_12007_7637# a_11923_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1670 a_30123_11305# a_29994_11049# a_29703_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1671 VPWR tdc0.w_dly_sig[167] tdc0.w_dly_sig_n[168] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1672 _026_ a_15351_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1673 a_30166_8725# a_29998_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1674 VGND a_29987_11445# a_29994_11745# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1675 tdc0.w_dly_sig_n[1] net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1676 _025_ a_14011_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X1677 a_30549_8041# a_29559_7669# a_30423_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1678 a_16974_12015# _059_ a_16894_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X1679 VGND tdc0.w_dly_sig[44] tdc0.w_dly_sig_n[45] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1681 _122_ a_12539_6688# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1682 VPWR a_11858_2879# a_11785_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1683 VPWR a_4222_3967# a_4149_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1684 VPWR a_20881_11721# uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1685 VGND tdc0.w_dly_sig[186] a_25757_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1687 VGND a_6671_4123# a_6629_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1688 a_11333_4765# tdc0.o_result[153] a_11251_4512# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1689 VPWR a_26514_6575# clknet_4_11_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1690 VPWR a_2915_4399# a_3083_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
R4 tt_um_hpretl_tt06_tdc_v1_7.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1693 a_1570_5487# a_1297_5493# a_1485_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1694 VGND tdc0.w_dly_sig[117] tdc0.w_dly_sig_n[117] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1695 a_20017_8029# _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1696 VPWR tdc0.w_dly_sig_n[160] tdc0.w_dly_sig[161] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1697 VPWR tdc0.w_dly_sig[58] tdc0.w_dly_sig_n[59] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1699 a_10037_13647# a_9871_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1700 a_25891_15823# a_25755_15797# a_25471_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1702 a_26667_8181# a_26951_8181# a_26886_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1703 VPWR a_19843_18543# a_20011_18517# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1704 _033_ a_17691_6281# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.965 w=0.65 l=0.15
X1705 VPWR a_23891_7663# a_24059_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1706 VPWR a_8879_7637# a_8795_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1707 a_24436_8751# _031_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1708 a_12341_11471# tdc0.w_dly_sig[75] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1709 a_26767_16885# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1711 tdc0.w_dly_sig[187] tdc0.w_dly_sig_n[185] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1714 VGND a_19843_18543# a_20011_18517# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1715 a_25247_7119# a_25111_7093# a_24827_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1716 VPWR a_29607_11623# tdc0.o_result[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1717 a_4314_7637# a_4146_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1718 VPWR a_6476_7637# clknet_4_1_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1719 VGND a_27503_5705# a_27510_5609# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1720 a_8251_12015# a_7387_12021# a_7994_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1721 a_18703_11721# _132_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1722 a_4521_15279# tdc0.w_dly_sig[103] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1723 VPWR _003_ a_24731_14423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1724 a_14868_8751# _115_ a_14766_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X1725 VPWR a_22971_957# a_23139_859# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1727 VPWR tdc0.o_result[131] a_11435_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1728 a_5989_13109# a_5823_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1729 a_21123_3133# a_20341_2767# a_21039_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1730 VGND _097_ a_17231_8457# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1731 tdc0.w_dly_sig_n[77] tdc0.w_dly_sig[77] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R5 tt_um_hpretl_tt06_tdc_v1_22.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1732 VPWR tdc0.w_dly_sig_n[69] tdc0.w_dly_sig[70] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1733 VPWR tdc0.w_dly_sig_n[191] tdc0.w_dly_sig[193] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1734 a_17312_9295# tdc0.o_result[24] a_16737_9441# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X1736 VPWR a_3302_15253# a_3229_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1737 a_26725_17277# a_26387_17063# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1738 VPWR a_25226_13621# a_25155_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1739 tdc0.w_dly_sig_n[90] tdc0.w_dly_sig[89] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1740 VGND tdc0.w_dly_sig[39] tdc0.w_dly_sig_n[40] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1741 a_20315_7895# tdc0.o_result[21] a_20549_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1742 VPWR tdc0.w_dly_sig_n[188] tdc0.w_dly_sig[189] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1743 tdc0.o_result[110] a_2347_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1744 VGND a_18059_7663# _001_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1745 VPWR tdc0.w_dly_sig_n[110] tdc0.w_dly_sig[111] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1746 net4 a_17634_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1748 a_22273_591# a_22107_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1749 VGND a_17130_16885# a_17059_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1750 a_16381_9295# tdc0.o_result[75] a_15943_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1751 VPWR a_22787_15279# a_22955_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1752 VPWR tdc0.w_dly_sig[54] tdc0.w_dly_sig_n[54] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1753 VGND tdc0.w_dly_sig_n[85] tdc0.w_dly_sig[87] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1754 a_10953_17999# a_9963_17999# a_10827_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1755 VGND tdc0.w_dly_sig_n[72] tdc0.w_dly_sig[74] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1756 tdc0.w_dly_sig_n[110] tdc0.w_dly_sig[109] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1757 VGND tdc0.w_dly_sig_n[89] tdc0.w_dly_sig[90] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1758 VGND clknet_4_4_0_clk a_1683_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1759 VPWR tdc0.w_dly_sig_n[25] tdc0.w_dly_sig[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1760 clknet_4_0_0_clk a_6476_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1761 VPWR a_16193_8725# _113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X1762 VGND a_22787_15279# a_22955_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1763 VPWR a_21431_8181# a_21438_8481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1764 VGND tdc0.w_dly_sig[105] tdc0.w_dly_sig_n[106] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1765 VGND _076_ a_13153_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1766 a_29703_11445# a_29987_11445# a_29922_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1767 uo_out[6] a_19777_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1768 VPWR a_2179_10927# a_2347_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1769 a_25226_3588# a_25026_3433# a_25375_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1770 tdc0.w_dly_sig[59] tdc0.w_dly_sig_n[57] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1771 VGND tdc0.w_dly_sig_n[44] tdc0.w_dly_sig[46] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1772 tdc0.w_dly_sig[115] tdc0.w_dly_sig_n[114] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1773 a_26387_17063# a_26483_16885# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1774 tdc0.w_dly_sig[22] tdc0.w_dly_sig_n[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1775 tdc0.w_dly_sig_n[138] tdc0.w_dly_sig[137] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1776 tdc0.w_dly_sig[94] tdc0.w_dly_sig_n[92] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1777 VPWR a_25428_7637# clknet_4_10_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1779 a_25954_2045# a_25707_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1780 a_25502_8181# a_25295_8181# a_25678_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1781 a_4245_2767# tdc0.w_dly_sig[156] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1782 a_3781_3855# a_3615_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1783 VGND tdc0.w_dly_sig[49] a_26309_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1784 tdc0.w_dly_sig_n[185] tdc0.w_dly_sig[185] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1785 VGND net6 _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1786 a_12153_11471# a_11987_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1787 tdc0.w_dly_sig[32] tdc0.w_dly_sig_n[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1788 VPWR a_6476_6549# clknet_4_0_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1789 VPWR _002_ a_15837_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1790 VGND tdc0.w_dly_sig_n[63] tdc0.w_dly_sig[64] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1791 tdc0.w_dly_sig_n[133] tdc0.w_dly_sig[132] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1792 tdc0.o_result[88] a_15779_17179# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1793 tdc0.o_result[164] a_11823_1947# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1794 a_30090_6397# a_29651_6031# a_30005_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1795 a_25077_9117# _012_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1796 VPWR tdc0.w_dly_sig_n[113] tdc0.w_dly_sig[115] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1797 a_14250_15253# a_14082_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1798 VGND tdc0.w_dly_sig[112] tdc0.w_dly_sig_n[113] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1799 a_19652_13897# _206_ a_19550_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X1800 VGND a_9815_7485# a_9983_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1801 a_19855_8359# _054_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X1802 clknet_0_clk a_16210_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1803 a_8378_2223# a_8105_2229# a_8293_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1804 VGND a_19855_7895# _115_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1806 a_16271_15797# a_16562_16097# a_16513_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1807 VPWR tdc0.o_result[99] a_17685_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1808 clknet_4_8_0_clk a_21104_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1810 a_27254_12381# a_26939_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1811 VGND a_26203_11623# tdc0.o_result[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1812 a_11785_3133# a_11251_2767# a_11690_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1813 VGND a_6550_12559# clknet_4_4_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1814 clknet_4_12_0_clk a_21380_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1815 VGND _011_ a_19807_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1816 VPWR a_30423_8751# a_30591_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1818 a_8565_9295# a_8399_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1819 VGND clknet_4_15_0_clk a_29559_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1820 a_24005_8725# _186_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X1821 tdc0.o_result[114] a_5291_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1822 a_14082_15279# a_13809_15285# a_13997_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1823 VGND a_17691_7119# _010_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1824 a_22457_3133# a_21923_2767# a_22362_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1825 VPWR net5 a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1826 VPWR tdc0.w_dly_sig_n[39] tdc0.w_dly_sig[41] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1827 a_25287_1653# a_25571_1653# a_25506_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1829 a_21717_14735# a_20727_14735# a_21591_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1831 a_3904_11305# a_3505_10933# a_3778_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1832 a_30711_6794# tdc0.w_dly_sig[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1833 VGND tdc0.w_dly_sig_n[126] tdc0.w_dly_sig[127] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1834 VGND clknet_4_0_0_clk a_3891_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1836 VGND a_18489_9839# uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1837 VPWR a_2715_13077# a_2631_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1838 a_13272_4719# tdc0.o_result[165] a_13082_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X1839 a_2248_12559# a_1849_12559# a_2122_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1840 a_14634_10927# a_14195_10933# a_14549_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1841 tdc0.w_dly_sig[59] tdc0.w_dly_sig_n[58] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1842 a_11597_4943# a_10607_4943# a_11471_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1843 a_30599_6397# a_29817_6031# a_30515_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1844 a_8933_16189# a_8399_15823# a_8838_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1845 tdc0.w_dly_sig_n[85] tdc0.w_dly_sig[85] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1846 a_21879_12711# a_21975_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1847 a_11329_14191# tdc0.w_dly_sig[85] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1848 a_9765_2223# tdc0.w_dly_sig[164] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1849 a_23975_7663# a_23193_7669# a_23891_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1850 VGND tdc0.w_dly_sig[81] tdc0.w_dly_sig_n[81] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1851 VGND _085_ a_16381_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X1852 VPWR a_6550_12559# clknet_4_4_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1853 VGND tdc0.w_dly_sig[158] tdc0.w_dly_sig_n[158] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1854 VPWR a_10627_4123# a_10543_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1855 a_12907_7119# _024_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1856 VGND tdc0.w_dly_sig[27] tdc0.w_dly_sig_n[27] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1857 VGND a_8638_16341# a_8596_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1859 a_5031_7485# a_4333_7119# a_4774_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1860 VPWR a_18647_16367# a_18815_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1861 a_5529_2767# a_5363_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1862 VGND a_19567_957# a_19735_859# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1864 tdc0.w_dly_sig_n[97] tdc0.w_dly_sig[96] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1866 a_13735_4512# _007_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1867 a_26309_4943# a_25762_5217# a_25962_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1868 VGND tdc0.w_dly_sig[83] tdc0.w_dly_sig_n[84] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1870 tdc0.w_dly_sig_n[51] tdc0.w_dly_sig[50] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1871 a_3877_4399# tdc0.w_dly_sig[149] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1872 VGND a_18647_16367# a_18815_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1873 a_3870_11837# a_3597_11471# a_3785_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1874 VGND tdc0.w_dly_sig[79] tdc0.w_dly_sig_n[79] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1875 a_2179_10927# a_1315_10933# a_1922_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1876 VPWR a_17194_2197# a_17121_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1877 a_25755_12533# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1878 a_27001_4399# a_26663_4631# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1879 VPWR tdc0.w_dly_sig_n[5] tdc0.w_dly_sig[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1880 VPWR tdc0.w_dly_sig[43] a_29437_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1881 a_29703_11159# a_29994_11049# a_29945_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1882 a_11141_6031# a_10975_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1883 a_7607_7485# a_6743_7119# a_7350_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1884 VPWR tdc0.w_dly_sig[168] tdc0.w_dly_sig_n[169] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1885 a_19058_4719# tdc0.o_result[151] a_18977_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X1886 tdc0.w_dly_sig[109] tdc0.w_dly_sig_n[108] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1887 a_7263_6005# clknet_4_3_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1889 VPWR a_1738_7231# a_1665_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1890 a_27123_5719# a_27219_5719# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1891 tdc0.w_dly_sig_n[20] tdc0.w_dly_sig[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1892 tdc0.w_dly_sig[140] tdc0.w_dly_sig_n[138] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1893 a_7967_10927# a_7185_10933# a_7883_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1894 tdc0.w_dly_sig[112] tdc0.w_dly_sig_n[111] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1895 tdc0.w_dly_sig[160] tdc0.w_dly_sig_n[158] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1896 VGND a_22311_5461# a_22269_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1897 VPWR a_27066_15556# a_26995_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1898 _134_ a_15943_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X1899 VPWR tdc0.w_dly_sig[157] tdc0.w_dly_sig_n[157] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1900 VGND _014_ a_15564_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1901 a_19890_13103# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1902 a_29621_16745# a_29074_16489# a_29274_16644# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1903 a_4333_15285# a_4167_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1904 clknet_4_9_0_clk a_22852_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1906 VPWR a_22891_6807# tdc0.o_result[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1907 VGND a_11839_6575# a_12007_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1908 VGND a_7683_10651# a_7641_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1909 a_8105_2229# a_7939_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1910 tdc0.w_dly_sig[31] tdc0.w_dly_sig_n[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1911 tdc0.w_dly_sig_n[132] tdc0.w_dly_sig[132] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1912 _047_ a_15101_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.38 ps=2.76 w=1 l=0.15
X1913 VPWR _038_ a_14703_3543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1914 VPWR net2 a_15023_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X1915 a_25111_7093# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1916 a_14507_15279# a_13809_15285# a_14250_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1917 a_23281_10383# a_22291_10383# a_23155_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1918 VPWR tdc0.w_dly_sig_n[115] tdc0.w_dly_sig[117] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1919 a_20359_11471# _016_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1920 a_19549_7485# a_19211_7271# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1921 a_14461_8207# tdc0.o_result[130] a_14379_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1922 VGND tdc0.w_dly_sig[173] tdc0.w_dly_sig_n[173] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1923 tdc0.w_dly_sig[2] tdc0.w_dly_sig_n[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1925 a_8481_10633# tdc0.o_result[128] a_8399_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1926 VPWR a_2290_13077# a_2217_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1928 a_25573_3689# a_25019_3529# a_25226_3588# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1929 tdc0.w_dly_sig_n[18] tdc0.w_dly_sig[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1931 a_4995_10633# _008_ a_5077_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1932 a_18305_10383# _001_ a_18233_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
R6 VPWR tt_um_hpretl_tt06_tdc_v1_8.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1933 VPWR a_4571_7663# a_4739_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1934 a_2037_13647# tdc0.w_dly_sig[107] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1935 VGND a_19225_11721# uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1937 a_12341_15823# tdc0.w_dly_sig[88] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1938 _184_ a_19899_3424# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1939 a_19142_957# a_18703_591# a_19057_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1941 a_4981_14735# tdc0.w_dly_sig[122] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1942 VGND a_15427_2223# a_15595_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1943 VGND clknet_4_9_0_clk a_21647_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1944 _053_ a_16850_13423# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X1945 tdc0.w_dly_sig_n[71] tdc0.w_dly_sig[71] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1946 VGND tdc0.w_dly_sig[125] tdc0.w_dly_sig_n[126] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1947 a_30423_8751# a_29559_8757# a_30166_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1949 VPWR a_15779_17179# a_15695_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1950 tdc0.w_dly_sig_n[47] tdc0.w_dly_sig[47] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1951 VGND _002_ a_18703_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X1952 VGND a_6476_7637# clknet_4_1_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1953 a_29725_8757# a_29559_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1954 a_17695_6575# _010_ _064_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1955 a_14805_6549# _079_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X1956 VPWR tdc0.w_dly_sig_n[47] tdc0.w_dly_sig[49] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1957 VGND tdc0.w_dly_sig_n[15] tdc0.w_dly_sig[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1958 VGND tdc0.w_dly_sig_n[75] tdc0.w_dly_sig[77] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1959 net6 a_18151_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1960 VGND tdc0.w_dly_sig[9] a_30541_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1962 a_30216_6031# a_29817_6031# a_30090_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1963 _178_ a_12907_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1964 tdc0.w_dly_sig[85] tdc0.w_dly_sig_n[84] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1965 a_29725_15285# a_29559_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1966 VGND tdc0.w_dly_sig[158] tdc0.w_dly_sig_n[159] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1967 tdc0.o_result[175] a_19183_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1968 a_23903_5095# a_23999_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1969 a_13153_4943# _024_ a_13081_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1970 VPWR tdc0.w_dly_sig_n[96] tdc0.w_dly_sig[97] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1971 a_27043_3829# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1972 a_16658_15101# a_16219_14735# a_16573_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1973 a_19015_2223# a_18151_2229# a_18758_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1974 a_23179_17673# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1975 tdc0.w_dly_sig_n[169] tdc0.w_dly_sig[168] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1976 a_19237_957# a_18703_591# a_19142_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1977 VPWR tdc0.w_dly_sig_n[117] tdc0.w_dly_sig[118] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1978 tdc0.w_dly_sig_n[171] tdc0.w_dly_sig[171] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1979 VGND _185_ a_19163_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1980 a_29203_16745# a_29067_16585# a_28783_16599# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1981 VPWR a_2547_14013# a_2715_13915# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1982 a_17695_6575# _010_ _064_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1983 tdc0.w_dly_sig_n[70] tdc0.w_dly_sig[69] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1984 a_29998_3311# a_29725_3317# a_29913_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1986 a_15611_17277# a_14913_16911# a_15354_17023# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1988 VPWR tdc0.w_dly_sig_n[170] tdc0.w_dly_sig[171] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1989 VPWR _085_ a_12356_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X1990 a_29541_9845# a_29375_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1991 a_29913_7663# tdc0.w_dly_sig[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1992 VGND tdc0.w_dly_sig[142] tdc0.w_dly_sig_n[143] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1993 tdc0.w_dly_sig_n[177] tdc0.w_dly_sig[177] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1994 tdc0.w_dly_sig_n[49] tdc0.w_dly_sig[49] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1995 a_17121_2223# a_16587_2229# a_17026_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1996 tdc0.o_result[11] a_30407_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1997 VPWR tdc0.o_result[83] a_14103_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1998 tdc0.w_dly_sig[160] tdc0.w_dly_sig_n[159] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1999 tdc0.w_dly_sig[107] tdc0.w_dly_sig_n[105] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2000 VPWR clknet_4_0_0_clk a_3891_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2001 a_7032_15657# a_6633_15285# a_6906_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2002 VPWR a_20211_15279# a_20379_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2003 VGND clknet_0_clk a_19890_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2004 VPWR tdc0.w_dly_sig_n[105] tdc0.w_dly_sig[106] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2005 VPWR a_27043_4617# a_27050_4521# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2006 VGND clknet_4_13_0_clk a_19347_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2008 a_2248_11471# a_1849_11471# a_2122_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2010 tdc0.w_dly_sig_n[13] tdc0.w_dly_sig[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2011 tdc0.o_result[143] a_8327_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2012 tdc0.w_dly_sig_n[162] tdc0.w_dly_sig[162] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2013 a_1665_7485# a_1131_7119# a_1570_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2014 a_29437_13481# a_28883_13321# a_29090_13380# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2015 tdc0.o_result[164] a_11823_1947# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2016 a_8838_14013# a_8399_13647# a_8753_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2017 VGND tdc0.w_dly_sig[79] tdc0.w_dly_sig_n[80] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2018 a_4609_6031# a_4443_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2020 VPWR a_10827_18365# a_10995_18267# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2021 VGND a_3099_7663# a_3267_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2022 tdc0.w_dly_sig[108] tdc0.w_dly_sig_n[107] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2023 a_1811_6397# a_947_6031# a_1554_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2024 VGND a_19395_7895# _158_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2026 tdc0.w_dly_sig_n[53] tdc0.w_dly_sig[53] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2027 tdc0.w_dly_sig[100] tdc0.w_dly_sig_n[99] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2028 a_5529_2767# a_5363_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2029 VGND tdc0.w_dly_sig[176] tdc0.w_dly_sig_n[177] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2030 _023_ a_13997_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.38 ps=2.76 w=1 l=0.15
X2031 a_2401_7669# a_2235_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2032 VPWR a_23139_13077# a_23055_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2033 VPWR a_4203_10927# a_4371_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2034 VPWR tdc0.w_dly_sig[159] tdc0.w_dly_sig_n[160] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2035 a_25559_3855# a_25339_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2036 a_23513_14557# _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X2037 a_22913_2767# a_21923_2767# a_22787_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2039 a_26909_8573# a_26571_8359# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2040 a_25663_14709# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2041 clknet_4_11_0_clk a_26514_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2042 VGND _200_ a_13722_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X2043 tdc0.o_result[85] a_12559_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2044 a_11655_2045# a_10957_1679# a_11398_1791# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2045 VGND clknet_4_0_0_clk a_4443_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2046 VPWR tdc0.w_dly_sig[59] tdc0.w_dly_sig_n[60] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2047 tdc0.w_dly_sig_n[155] tdc0.w_dly_sig[154] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2048 VGND _010_ a_18479_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2049 a_23455_11145# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2050 a_18737_6059# _030_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X2051 VPWR a_19225_11721# uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2052 VPWR tdc0.w_dly_sig[15] tdc0.w_dly_sig_n[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2053 tdc0.o_result[85] a_12559_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2054 VGND tdc0.w_dly_sig_n[71] tdc0.w_dly_sig[73] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2055 VPWR a_26882_12559# clknet_4_14_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2056 a_20421_6031# a_19874_6305# a_20074_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2057 VPWR a_21051_8359# tdc0.o_result[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2058 tdc0.w_dly_sig_n[44] tdc0.w_dly_sig[44] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2059 VGND a_18843_13335# _140_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2060 VPWR a_12851_16189# a_13019_16091# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2061 a_23466_7663# a_23027_7669# a_23381_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2064 a_30343_7284# tdc0.w_dly_sig[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2065 VGND a_5199_15253# a_5157_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2066 tdc0.w_dly_sig_n[112] tdc0.w_dly_sig[112] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2067 VPWR tdc0.w_dly_sig_n[83] tdc0.w_dly_sig[85] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2068 clknet_4_15_0_clk a_25410_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2069 _087_ a_11159_8864# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2070 a_20341_2767# a_20175_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2071 VGND a_10903_13915# a_10861_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2072 VGND a_5291_11989# a_5249_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2073 tdc0.w_dly_sig[149] tdc0.w_dly_sig_n[148] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2074 tdc0.o_result[100] a_4739_17179# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2075 VPWR a_25755_12533# a_25762_12833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2076 a_15285_12559# tdc0.w_dly_sig[73] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2077 a_25755_4917# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2078 clknet_4_2_0_clk a_11260_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2079 a_11873_9295# a_10883_9295# a_11747_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2080 VPWR a_18003_18365# a_18171_18267# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2081 VPWR a_23179_17673# a_23186_17577# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2082 a_14151_10535# tdc0.o_result[89] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2083 VPWR tdc0.w_dly_sig_n[51] tdc0.w_dly_sig[52] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2084 a_29725_3317# a_29559_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2085 _018_ a_17503_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X2086 a_29922_11293# a_29607_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2087 tdc0.w_dly_sig[171] tdc0.w_dly_sig_n[170] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2088 a_11839_6397# a_10975_6031# a_11582_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2089 tdc0.w_dly_sig_n[50] tdc0.w_dly_sig[49] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2090 VGND tdc0.w_dly_sig[40] tdc0.w_dly_sig_n[41] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2091 a_14255_6835# _013_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X2092 VPWR tdc0.w_dly_sig[131] tdc0.w_dly_sig_n[132] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2093 VPWR tdc0.w_dly_sig_n[88] tdc0.w_dly_sig[90] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2094 VPWR tdc0.w_dly_sig[144] tdc0.w_dly_sig_n[145] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2095 VPWR tdc0.w_dly_sig[11] tdc0.w_dly_sig_n[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2097 VGND a_6430_13077# a_6388_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2098 _121_ a_14274_13423# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X2099 VGND a_29515_4631# tdc0.o_result[191] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2100 a_23055_16189# a_22273_15823# a_22971_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2101 VGND a_23155_10749# a_23323_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2102 tdc0.w_dly_sig_n[88] tdc0.w_dly_sig[87] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2103 VGND tdc0.w_dly_sig[94] tdc0.w_dly_sig_n[94] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2105 VGND a_30258_6143# a_30216_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2106 tdc0.w_dly_sig_n[36] tdc0.w_dly_sig[35] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2108 VPWR a_8546_2197# a_8473_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2109 VGND a_15227_10901# a_15185_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2110 VGND a_22891_14423# _147_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2111 a_18703_11721# _134_ a_18953_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2112 a_16753_2229# a_16587_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2113 VPWR a_20325_5089# _197_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X2115 VGND a_29423_6196# net28 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2116 VPWR a_20417_4373# _185_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X2117 a_16842_17455# a_16403_17461# a_16757_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2118 a_6687_13103# a_5989_13109# a_6430_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2119 VGND tdc0.w_dly_sig_n[78] tdc0.w_dly_sig[79] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2120 VGND tdc0.o_result[28] a_23124_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X2121 clknet_4_10_0_clk a_25428_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2122 VPWR tdc0.w_dly_sig[115] tdc0.w_dly_sig_n[115] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2123 a_4203_10927# a_3339_10933# a_3946_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2124 tdc0.w_dly_sig_n[44] tdc0.w_dly_sig[43] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2125 VPWR a_12759_9839# a_12927_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2126 VPWR a_2658_4373# a_2585_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2127 a_10037_13647# a_9871_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2128 VGND tdc0.w_dly_sig[172] tdc0.w_dly_sig_n[173] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2129 uo_out[1] a_24653_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2130 a_7166_14165# a_6998_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2131 tdc0.w_dly_sig[9] tdc0.w_dly_sig_n[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2132 a_27043_3829# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2133 a_12337_5493# a_12171_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2134 a_12475_15279# a_11693_15285# a_12391_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2135 a_5602_15935# a_5434_16189# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2136 tdc0.o_result[117] a_4739_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2137 VGND _112_ a_17967_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2138 VGND a_2715_13077# a_2673_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2139 a_26309_12559# a_25762_12833# a_25962_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2140 a_27035_12247# a_27319_12233# a_27254_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2141 _005_ a_15203_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2142 VPWR _018_ a_18703_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2143 VPWR _064_ a_21071_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2144 VGND a_21914_11204# a_21843_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2145 a_16293_591# a_16127_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2146 VGND a_1995_7485# a_2163_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2147 a_9263_8573# a_8565_8207# a_9006_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2148 VGND tdc0.w_dly_sig_n[59] tdc0.w_dly_sig[60] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2149 a_4521_7119# tdc0.w_dly_sig[134] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2150 tdc0.w_dly_sig_n[16] tdc0.w_dly_sig[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2151 VGND tdc0.w_dly_sig[37] tdc0.w_dly_sig_n[37] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2153 a_4571_7663# a_3707_7669# a_4314_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2154 VPWR tdc0.o_result[124] a_12723_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2155 VGND a_7515_10749# a_7683_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2156 VPWR a_14703_3543# _073_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2157 VGND a_12594_14847# a_12552_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2158 VGND clknet_4_8_0_clk a_18151_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2160 a_14913_16911# a_14747_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2161 a_19796_13647# tdc0.o_result[39] a_19221_13793# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X2162 VPWR _023_ a_12448_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X2163 a_26667_8983# a_26958_8873# a_26909_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2165 tdc0.w_dly_sig_n[113] tdc0.w_dly_sig[113] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2166 tdc0.w_dly_sig[98] tdc0.w_dly_sig_n[97] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2167 VGND clknet_0_clk a_21104_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2168 VGND tdc0.w_dly_sig_n[132] tdc0.w_dly_sig[134] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2169 VGND a_26859_15497# a_26866_15401# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2170 VGND clknet_4_12_0_clk a_21739_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2172 VGND tdc0.w_dly_sig_n[41] tdc0.w_dly_sig[43] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2173 _192_ a_6191_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2174 tdc0.w_dly_sig_n[6] tdc0.w_dly_sig[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2175 a_25410_3829# a_25210_4129# a_25559_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2176 a_17187_13799# tdc0.o_result[64] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2177 VGND _051_ a_23457_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2178 a_19225_11721# tdc0.o_result[4] a_18703_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X2179 _121_ a_14274_13423# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X2180 a_4421_11471# a_3431_11471# a_4295_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2181 VPWR a_7775_7387# a_7691_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2183 _107_ a_21923_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2184 VPWR a_18059_7663# _001_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2185 a_23937_14985# _055_ a_24021_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2186 clknet_4_1_0_clk a_6476_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2187 a_19169_3677# _060_ a_19097_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2188 _076_ a_14064_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2189 a_5031_7485# a_4167_7119# a_4774_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2190 VGND tdc0.w_dly_sig[64] tdc0.w_dly_sig_n[64] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2191 a_22971_957# a_22273_591# a_22714_703# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2193 a_2306_9839# a_2033_9845# a_2221_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2194 tdc0.w_dly_sig[16] tdc0.w_dly_sig_n[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2195 VGND a_21431_8181# a_21438_8481# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2196 a_23269_9813# _126_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X2197 a_25663_14709# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2198 a_12723_6031# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2199 VPWR tdc0.w_dly_sig_n[130] tdc0.w_dly_sig[132] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2200 a_25011_8181# a_25302_8481# a_25253_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2201 a_13997_17455# tdc0.w_dly_sig[91] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2202 VGND a_17194_2197# a_17152_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2203 VPWR tdc0.w_dly_sig_n[144] tdc0.w_dly_sig[145] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2204 a_23592_8041# a_23193_7669# a_23466_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2205 a_24131_9545# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2206 VGND a_27066_15556# a_26995_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2207 VGND tdc0.w_dly_sig[145] tdc0.w_dly_sig_n[146] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2208 VGND tdc0.w_dly_sig_n[147] tdc0.w_dly_sig[149] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2209 VGND a_25318_11445# a_25247_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2210 tdc0.w_dly_sig_n[178] tdc0.w_dly_sig[177] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2211 a_19487_6183# a_19583_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2212 VPWR ui_in[3] a_15575_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2213 VGND _210_ a_20175_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2214 VPWR a_4739_17179# a_4655_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2215 VGND tdc0.w_dly_sig_n[183] tdc0.w_dly_sig[184] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2216 VPWR a_11812_13621# clknet_4_7_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2217 VGND tdc0.w_dly_sig[171] tdc0.w_dly_sig_n[172] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2218 a_19727_7119# a_19591_7093# a_19307_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2219 VPWR tdc0.w_dly_sig[7] tdc0.w_dly_sig_n[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2220 a_16645_11989# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X2221 tdc0.w_dly_sig_n[71] tdc0.w_dly_sig[70] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2222 a_12594_15935# a_12426_16189# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2224 a_14208_17833# a_13809_17461# a_14082_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2225 tdc0.o_result[69] a_17251_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2226 a_14116_2767# a_13717_2767# a_13990_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2227 a_20341_2767# a_20175_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2228 VPWR tdc0.o_result[130] a_14379_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2229 VGND tdc0.w_dly_sig[102] tdc0.w_dly_sig_n[102] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2230 tdc0.o_result[166] a_12283_1109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2231 a_16761_10927# _008_ a_16845_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2232 VPWR a_17507_1143# net5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2233 a_29331_7284# tdc0.w_dly_sig[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2235 a_8473_2223# a_7939_2229# a_8378_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2236 a_11287_8573# a_10589_8207# a_11030_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2237 VGND a_19586_18517# a_19544_18921# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2238 a_22530_2879# a_22362_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2240 a_17923_5719# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.142 ps=1.34 w=0.42 l=0.15
X2241 a_7182_7485# a_6743_7119# a_7097_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2242 tdc0.w_dly_sig[116] tdc0.w_dly_sig_n[115] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2243 a_5066_15101# a_4793_14735# a_4981_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2244 a_23420_5807# _060_ a_23300_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X2245 a_1811_6397# a_1113_6031# a_1554_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2246 a_18980_8457# tdc0.o_result[101] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X2247 a_12759_9839# a_12061_9845# a_12502_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2248 a_2497_6575# tdc0.w_dly_sig[151] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2249 tdc0.w_dly_sig[57] tdc0.w_dly_sig_n[56] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2250 a_7378_13103# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2251 VPWR a_30591_8725# a_30507_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2252 VGND a_16210_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2253 a_11325_18549# a_11159_18549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2254 a_9761_3855# a_9595_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2255 a_12334_9839# a_11895_9845# a_12249_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2256 a_17876_4399# tdc0.o_result[148] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X2257 a_2585_4399# a_2051_4405# a_2490_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2258 tdc0.w_dly_sig_n[23] tdc0.w_dly_sig[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2259 VGND a_22971_16189# a_23139_16091# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2260 VGND _042_ a_17231_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2261 VPWR clknet_0_clk a_22852_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2262 a_19843_18543# a_19145_18549# a_19586_18517# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2263 VGND a_30194_11204# a_30123_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2264 a_24653_9545# tdc0.o_result[1] a_24131_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X2265 a_13537_16367# tdc0.w_dly_sig[90] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2266 a_20325_5089# _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X2267 VGND _037_ a_16587_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X2268 a_11527_3855# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2269 a_12843_9839# a_12061_9845# a_12759_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2270 VGND tdc0.w_dly_sig_n[125] tdc0.w_dly_sig[127] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2271 VGND tdc0.w_dly_sig_n[74] tdc0.w_dly_sig[75] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2273 a_15538_12671# a_15370_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2274 VGND tdc0.w_dly_sig[28] tdc0.w_dly_sig_n[28] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2275 tdc0.o_result[124] a_9431_13915# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2276 a_23237_3855# _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X2277 VGND a_11639_5211# a_11597_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2278 tdc0.w_dly_sig[146] tdc0.w_dly_sig_n[145] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2279 _172_ a_5639_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X2280 a_26995_15657# a_26866_15401# a_26575_15511# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2281 _059_ a_16495_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2282 tdc0.w_dly_sig[1] tdc0.w_dly_sig_n[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2283 VGND _068_ a_18037_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2284 a_15163_3543# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2285 a_11490_9407# a_11322_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2286 VGND tdc0.w_dly_sig[187] tdc0.w_dly_sig_n[188] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2287 tdc0.w_dly_sig[79] tdc0.w_dly_sig_n[77] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2288 _006_ net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2290 VPWR tdc0.w_dly_sig[47] tdc0.w_dly_sig_n[48] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2291 VGND tdc0.w_dly_sig[75] tdc0.w_dly_sig_n[75] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2292 a_26019_14735# a_25799_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2293 VPWR a_10091_4399# a_10259_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2294 a_7626_10901# a_7458_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2295 VGND _018_ a_18703_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2296 a_28595_7284# tdc0.w_dly_sig[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2297 a_8745_10383# tdc0.o_result[112] a_8399_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2298 a_18059_11721# _141_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2299 a_20525_1679# a_20359_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2300 _024_ net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2301 a_15101_16911# tdc0.w_dly_sig[89] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2302 a_24309_15599# _017_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X2303 a_14195_3424# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2304 a_5115_11159# tdc0.o_result[108] a_5261_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X2306 VGND _035_ a_15232_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X2307 a_2673_13481# a_1683_13109# a_2547_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2308 _042_ a_16401_6691# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2309 VPWR a_10662_14847# a_10589_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2310 tdc0.w_dly_sig_n[45] tdc0.w_dly_sig[44] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2311 tdc0.w_dly_sig_n[182] tdc0.w_dly_sig[181] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2312 tdc0.w_dly_sig_n[93] tdc0.w_dly_sig[92] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2314 a_29019_13481# a_28890_13225# a_28599_13335# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2315 VPWR tdc0.o_result[87] a_12999_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2316 VPWR tdc0.w_dly_sig_n[141] tdc0.w_dly_sig[143] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2317 VPWR tdc0.w_dly_sig_n[143] tdc0.w_dly_sig[145] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2318 uo_out[0] a_20881_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2319 tdc0.w_dly_sig_n[179] tdc0.w_dly_sig[178] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2320 a_16991_957# a_16127_591# a_16734_703# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2321 VGND a_18151_1135# net6 VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2323 tdc0.w_dly_sig_n[167] tdc0.w_dly_sig[167] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2324 tdc0.w_dly_sig_n[170] tdc0.w_dly_sig[170] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2325 tdc0.w_dly_sig_n[162] tdc0.w_dly_sig[161] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2326 a_12815_2767# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2327 clknet_4_6_0_clk a_12254_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2328 a_27675_10205# a_27455_10217# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2329 a_9006_13759# a_8838_14013# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2330 a_18383_8983# _019_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2331 VPWR _022_ a_16219_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2332 a_25471_15797# a_25762_16097# a_25713_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2333 a_19058_4719# _204_ a_19304_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X2335 a_25757_3855# a_25203_3829# a_25410_3829# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2336 _180_ a_13367_9952# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2337 VPWR tdc0.w_dly_sig_n[179] tdc0.w_dly_sig[181] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2338 VGND tdc0.w_dly_sig_n[26] tdc0.w_dly_sig[27] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2339 VGND tdc0.w_dly_sig_n[24] tdc0.w_dly_sig[26] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2340 a_27219_5719# a_27510_5609# a_27461_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2341 VGND tdc0.w_dly_sig_n[134] tdc0.w_dly_sig[135] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2342 VGND tdc0.w_dly_sig_n[151] tdc0.w_dly_sig[152] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2343 a_25111_7093# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2344 a_12199_3133# a_11417_2767# a_12115_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2345 tdc0.w_dly_sig_n[187] tdc0.w_dly_sig[187] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2347 VPWR a_23082_8725# a_23009_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2348 a_16193_8725# _068_ a_16350_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2349 VGND tdc0.w_dly_sig[118] tdc0.w_dly_sig_n[119] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2350 a_16991_18543# a_16127_18549# a_16734_18517# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2351 tdc0.w_dly_sig[50] tdc0.w_dly_sig_n[48] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2352 a_13552_9545# tdc0.o_result[126] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X2353 a_6725_3317# a_6559_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2354 a_22021_3677# _060_ a_21949_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2355 a_24009_13647# _003_ a_23937_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2356 VGND a_6855_4373# a_6813_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2357 a_10402_18365# a_9963_17999# a_10317_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2359 VGND tdc0.w_dly_sig_n[73] tdc0.w_dly_sig[75] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2361 VPWR clknet_4_7_0_clk a_11159_18549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2362 VPWR _064_ a_24659_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2363 a_17691_6281# _000_ a_17773_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2365 a_16661_18543# a_16127_18549# a_16566_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2366 VPWR tdc0.w_dly_sig_n[32] tdc0.w_dly_sig[34] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2367 a_2309_6581# a_2143_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2370 tdc0.w_dly_sig[67] tdc0.w_dly_sig_n[66] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2371 VGND a_14011_5487# _025_ VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2372 a_12989_7119# tdc0.o_result[134] a_12907_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2373 VPWR a_12023_18543# a_12191_18517# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2374 VPWR tdc0.w_dly_sig_n[135] tdc0.w_dly_sig[136] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2375 a_20003_11305# a_19874_11049# a_19583_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2376 a_19058_4719# _203_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X2377 VGND a_2179_10927# a_2347_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2378 VPWR tdc0.w_dly_sig_n[2] tdc0.w_dly_sig[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2379 VGND a_4295_11837# a_4463_11739# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2380 VGND tdc0.w_dly_sig[50] a_24837_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2381 a_20315_7895# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2382 a_17415_10927# _094_ a_17665_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2383 VGND a_12023_18543# a_12191_18517# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2384 VGND tdc0.w_dly_sig[29] tdc0.w_dly_sig_n[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2385 VPWR _017_ a_24021_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X2386 VGND a_14158_2879# a_14116_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2387 VPWR _047_ a_5077_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2388 a_24065_3855# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X2389 a_24113_14191# tdc0.o_result[45] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2390 a_26583_11445# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2391 a_17233_6281# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2392 VGND a_11087_15003# a_11045_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2393 a_16205_10901# _012_ a_16451_11265# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2394 VGND tdc0.w_dly_sig[22] a_25665_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2395 VPWR clknet_4_7_0_clk a_13183_16373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2396 tdc0.w_dly_sig[74] tdc0.w_dly_sig_n[72] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2397 tdc0.w_dly_sig[173] tdc0.w_dly_sig_n[172] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2398 VPWR tdc0.w_dly_sig[20] tdc0.w_dly_sig_n[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2399 a_16210_9839# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2400 tdc0.w_dly_sig[90] tdc0.w_dly_sig_n[89] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2401 VPWR a_25295_8181# a_25302_8481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2402 a_29909_9839# a_29375_9845# a_29814_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2403 _208_ a_18703_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2404 VPWR a_27411_13321# a_27418_13225# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2405 a_7308_7119# a_6909_7119# a_7182_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2406 tdc0.w_dly_sig_n[106] tdc0.w_dly_sig[105] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2407 VGND _018_ a_18305_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2408 VPWR a_5199_7387# a_5115_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2409 tdc0.w_dly_sig[147] tdc0.w_dly_sig_n[146] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2410 VGND _043_ a_14257_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2411 a_11582_6143# a_11414_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2412 a_3969_3855# tdc0.w_dly_sig[154] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2413 a_22751_12015# _004_ a_22929_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X2414 a_9006_9407# a_8838_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2415 VGND tdc0.w_dly_sig_n[35] tdc0.w_dly_sig[37] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2417 tdc0.w_dly_sig[170] tdc0.w_dly_sig_n[169] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2418 a_8841_17455# a_8307_17461# a_8746_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2420 tdc0.w_dly_sig[30] tdc0.w_dly_sig_n[28] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2421 a_21914_17732# a_21714_17577# a_22063_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2422 VGND tdc0.w_dly_sig_n[143] tdc0.w_dly_sig[144] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2423 VGND a_13019_16091# a_12977_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2424 a_9761_3855# a_9595_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2425 tdc0.w_dly_sig[8] tdc0.w_dly_sig_n[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2426 a_22304_16911# a_21905_16911# a_22178_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2427 VPWR a_17323_6575# _030_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2428 a_9006_9407# a_8838_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2429 VPWR clknet_4_6_0_clk a_11987_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2430 VGND tdc0.w_dly_sig[190] tdc0.w_dly_sig_n[190] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2431 tdc0.w_dly_sig[94] tdc0.w_dly_sig_n[93] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2433 VPWR a_22679_4373# a_22595_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2434 _194_ a_23855_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2435 a_24653_9545# _064_ a_24131_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2436 clknet_4_12_0_clk a_21380_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X2437 VPWR clknet_4_6_0_clk a_14931_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2438 a_16350_8751# tdc0.o_result[155] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2439 a_3873_16911# a_3707_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2440 tdc0.w_dly_sig[181] tdc0.w_dly_sig_n[179] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2441 a_6262_5487# a_5989_5493# a_6177_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2442 VGND tdc0.w_dly_sig_n[129] tdc0.w_dly_sig[130] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2443 tdc0.w_dly_sig[104] tdc0.w_dly_sig_n[102] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2444 tdc0.w_dly_sig[164] tdc0.w_dly_sig_n[162] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2445 tdc0.o_result[149] a_2163_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2446 tdc0.w_dly_sig[173] tdc0.w_dly_sig_n[171] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2447 tdc0.o_result[147] a_4279_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2448 a_19583_6005# a_19874_6305# a_19825_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2449 VGND a_7166_3285# a_7124_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2450 VPWR a_11260_5461# clknet_4_2_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2452 a_4130_4373# a_3962_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2453 a_11049_9295# a_10883_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2454 a_22615_4007# tdc0.o_result[189] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2455 a_8385_16367# tdc0.w_dly_sig[98] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2456 VPWR a_30347_10357# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2457 VGND tdc0.w_dly_sig[110] tdc0.w_dly_sig_n[110] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2459 VGND tdc0.w_dly_sig[24] tdc0.w_dly_sig_n[25] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2460 VGND a_27158_8181# a_27087_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2461 tdc0.o_result[132] a_5475_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2462 a_14101_10159# _072_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X2463 tdc0.w_dly_sig[49] tdc0.w_dly_sig_n[47] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2464 a_4866_8725# a_4698_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2465 VGND tdc0.w_dly_sig_n[46] tdc0.w_dly_sig[47] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2466 a_30194_11445# a_29994_11745# a_30343_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2467 VPWR a_10735_12925# a_10903_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2468 VGND a_25962_12533# a_25891_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2469 a_14549_10927# tdc0.w_dly_sig[77] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
R7 tt_um_hpretl_tt06_tdc_v1_13.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2470 tdc0.w_dly_sig_n[95] tdc0.w_dly_sig[94] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2471 tdc0.o_result[101] a_7499_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2472 a_17557_4971# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2473 tdc0.w_dly_sig[69] tdc0.w_dly_sig_n[68] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2474 tdc0.w_dly_sig[41] tdc0.w_dly_sig_n[39] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2475 VGND a_22714_13077# a_22672_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2476 VGND _090_ a_24131_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2477 tdc0.w_dly_sig[127] tdc0.w_dly_sig_n[126] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2478 uo_out[3] a_18489_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2480 VPWR tdc0.w_dly_sig_n[3] tdc0.w_dly_sig[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2482 tdc0.o_result[101] a_7499_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2483 tdc0.w_dly_sig[20] tdc0.w_dly_sig_n[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2484 VGND a_19310_703# a_19268_591# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2485 a_4839_3133# a_4057_2767# a_4755_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2486 a_21633_5487# tdc0.w_dly_sig[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2487 VGND a_2842_7637# a_2800_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2488 a_19786_15279# a_19513_15285# a_19701_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2489 VPWR clknet_4_1_0_clk a_5823_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2490 _090_ a_14563_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X2491 tdc0.w_dly_sig[62] tdc0.w_dly_sig_n[61] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2493 a_17415_11247# _110_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2495 a_13790_16341# a_13622_16367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2496 VPWR clknet_4_5_0_clk a_8399_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2497 tdc0.w_dly_sig_n[81] tdc0.w_dly_sig[81] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2498 a_16366_2879# a_16198_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2499 VGND tdc0.w_dly_sig_n[121] tdc0.w_dly_sig[122] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2500 VPWR tdc0.w_dly_sig[135] tdc0.w_dly_sig_n[135] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2501 VGND a_23507_8725# a_23465_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2502 VGND a_5291_8725# a_5249_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2503 tdc0.w_dly_sig_n[69] tdc0.w_dly_sig[69] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2504 a_22971_13103# a_22273_13109# a_22714_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2505 a_22217_12925# a_21879_12711# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2506 a_9263_8573# a_8399_8207# a_9006_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2507 a_10267_9839# a_9485_9845# a_10183_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2509 VGND a_1922_10901# a_1880_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2510 a_23303_8207# _010_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2511 a_5851_9661# a_5069_9295# a_5767_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2512 VPWR tdc0.w_dly_sig[154] tdc0.w_dly_sig_n[154] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2513 tdc0.w_dly_sig[115] tdc0.w_dly_sig_n[113] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2514 VGND a_26882_12559# clknet_4_14_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X2515 a_4793_12015# a_4259_12021# a_4698_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2516 a_30010_5764# a_29810_5609# a_30159_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2517 VGND a_16547_7093# _022_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2519 tdc0.o_result[104] a_3727_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2520 a_23097_13481# a_22107_13109# a_22971_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2521 a_23585_14557# _012_ a_23513_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2522 net1 a_30347_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2523 tdc0.w_dly_sig[148] tdc0.w_dly_sig_n[146] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2524 VPWR a_16734_18517# a_16661_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2525 VGND a_25755_12533# a_25762_12833# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2526 VPWR a_2474_9813# a_2401_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2527 a_2857_10217# a_1867_9845# a_2731_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2528 VPWR clknet_4_1_0_clk a_6743_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2529 VGND tdc0.w_dly_sig[66] tdc0.w_dly_sig_n[67] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2530 clknet_4_9_0_clk a_22852_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2531 a_22714_13077# a_22546_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2532 clknet_4_9_0_clk a_22852_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X2533 tdc0.o_result[104] a_3727_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2534 a_9949_2767# tdc0.w_dly_sig[163] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2535 tdc0.o_result[138] a_10627_4123# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2536 VGND _124_ a_12618_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X2537 VGND a_20782_2879# a_20740_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2538 clknet_4_8_0_clk a_21104_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2539 a_29871_5309# a_29173_4943# a_29614_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2540 VPWR net5 a_17503_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2541 VGND tdc0.w_dly_sig[86] tdc0.w_dly_sig_n[87] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2542 VGND a_30423_14191# a_30591_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2543 VGND a_6503_4221# a_6671_4123# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2544 a_16923_16885# clknet_4_12_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2545 VPWR tdc0.w_dly_sig_n[184] tdc0.w_dly_sig[186] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2546 VPWR tdc0.w_dly_sig[98] tdc0.w_dly_sig_n[98] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2547 a_12426_11837# a_11987_11471# a_12341_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2548 a_8285_4777# a_7295_4405# a_8159_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2549 a_30507_7663# a_29725_7669# a_30423_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2550 tdc0.w_dly_sig_n[29] tdc0.w_dly_sig[28] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2551 a_10091_4399# a_9227_4405# a_9834_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2553 a_6998_3311# a_6559_3317# a_6913_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2554 a_17937_10927# tdc0.o_result[2] a_17415_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X2555 VGND tdc0.w_dly_sig_n[89] tdc0.w_dly_sig[91] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2556 VPWR clknet_4_5_0_clk a_4167_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2557 a_22546_13103# a_22273_13109# a_22461_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2559 a_26951_8181# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2560 a_23913_8353# _106_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X2561 a_18127_10927# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2562 a_20981_9295# tdc0.o_result[65] a_20543_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2563 VPWR tdc0.w_dly_sig[149] tdc0.w_dly_sig_n[150] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2564 VPWR tdc0.w_dly_sig_n[144] tdc0.w_dly_sig[146] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2565 a_14633_18921# a_13643_18549# a_14507_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2566 VGND tdc0.w_dly_sig[64] tdc0.w_dly_sig_n[65] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2567 tdc0.w_dly_sig_n[184] tdc0.w_dly_sig[183] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2568 VGND tdc0.w_dly_sig[147] tdc0.w_dly_sig_n[148] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2569 tdc0.w_dly_sig[166] tdc0.w_dly_sig_n[164] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2571 a_2079_7485# a_1297_7119# a_1995_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2572 VGND a_2715_12827# a_2673_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2573 VPWR a_8914_17429# a_8841_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2574 a_25226_3588# a_25019_3529# a_25402_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2575 VGND _040_ a_20359_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2576 clknet_4_3_0_clk a_10506_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2578 VPWR tdc0.w_dly_sig_n[16] tdc0.w_dly_sig[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2579 VGND a_7350_7231# a_7308_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2580 tdc0.o_result[84] a_12007_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2581 a_18913_4943# _011_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X2582 a_11965_6953# a_10975_6581# a_11839_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2583 tdc0.w_dly_sig_n[55] tdc0.w_dly_sig[55] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2584 VGND tdc0.w_dly_sig[146] tdc0.w_dly_sig_n[147] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2585 a_26951_8969# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2586 a_7415_15279# a_6633_15285# a_7331_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2587 VGND _072_ a_7917_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X2588 a_19786_15279# a_19347_15285# a_19701_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2589 a_3352_14569# a_2953_14197# a_3226_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2590 VGND tdc0.w_dly_sig_n[154] tdc0.w_dly_sig[155] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2591 VGND tdc0.w_dly_sig[189] a_27597_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2594 tdc0.w_dly_sig[71] tdc0.w_dly_sig_n[69] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2595 a_10225_12559# tdc0.w_dly_sig[82] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2596 VPWR a_6883_6183# tdc0.o_result[136] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2597 a_11287_8573# a_10423_8207# a_11030_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2598 a_17201_3677# _038_ a_17129_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2599 a_22871_15279# a_22089_15285# a_22787_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2600 VPWR tdc0.w_dly_sig[42] tdc0.w_dly_sig_n[43] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2601 a_19583_11159# a_19874_11049# a_19825_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2602 _114_ a_15943_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X2603 tdc0.w_dly_sig_n[130] tdc0.w_dly_sig[129] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2604 a_4061_16911# tdc0.w_dly_sig[101] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2605 a_23110_5807# tdc0.o_result[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X2606 a_9305_7119# tdc0.w_dly_sig[135] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2607 tdc0.w_dly_sig[52] tdc0.w_dly_sig_n[51] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2608 tdc0.w_dly_sig[78] tdc0.w_dly_sig_n[76] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2609 a_7783_3133# a_7001_2767# a_7699_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2610 VGND tdc0.w_dly_sig[181] a_24745_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2611 a_30010_5764# a_29803_5705# a_30186_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2612 tdc0.w_dly_sig_n[23] tdc0.w_dly_sig[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2613 VPWR tdc0.w_dly_sig_n[118] tdc0.w_dly_sig[120] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2615 VPWR clknet_4_2_0_clk a_11251_1141# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2616 VPWR tdc0.w_dly_sig_n[81] tdc0.w_dly_sig[82] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2617 VGND tdc0.w_dly_sig[36] tdc0.w_dly_sig_n[37] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2618 a_22641_8757# a_22475_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2619 VGND tdc0.w_dly_sig[164] tdc0.w_dly_sig_n[164] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2620 tdc0.w_dly_sig[142] tdc0.w_dly_sig_n[140] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2621 tdc0.w_dly_sig_n[143] tdc0.w_dly_sig[142] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2622 VGND a_12007_6549# a_11965_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2623 VGND a_3651_3311# a_3819_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2624 VGND tdc0.w_dly_sig_n[82] tdc0.w_dly_sig[84] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2625 VPWR tdc0.w_dly_sig_n[136] tdc0.w_dly_sig[138] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2626 _188_ a_23303_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2627 tdc0.w_dly_sig[56] tdc0.w_dly_sig_n[55] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2628 tdc0.w_dly_sig_n[153] tdc0.w_dly_sig[153] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2629 a_21445_5493# a_21279_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2631 a_4130_4373# a_3962_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2632 tdc0.w_dly_sig_n[80] tdc0.w_dly_sig[80] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2633 a_19310_703# a_19142_957# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2634 tdc0.w_dly_sig[117] tdc0.w_dly_sig_n[115] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2635 a_22063_11293# a_21843_11305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2636 VGND a_25226_3588# a_25155_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2637 VGND clknet_4_0_0_clk a_2787_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2639 VGND tdc0.w_dly_sig_n[86] tdc0.w_dly_sig[87] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2640 tdc0.w_dly_sig[177] tdc0.w_dly_sig_n[175] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2641 a_15023_5309# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2642 a_2217_4405# a_2051_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2643 tdc0.w_dly_sig_n[145] tdc0.w_dly_sig[145] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2644 VGND a_26514_6575# clknet_4_11_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2646 VGND a_25870_14709# a_25799_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2647 a_12539_6688# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2648 tdc0.w_dly_sig[58] tdc0.w_dly_sig_n[57] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2649 VGND tdc0.w_dly_sig_n[181] tdc0.w_dly_sig[183] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2651 VPWR clknet_4_10_0_clk a_29559_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2652 tdc0.w_dly_sig[125] tdc0.w_dly_sig_n[123] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2653 tdc0.w_dly_sig[119] tdc0.w_dly_sig_n[117] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2654 VGND clknet_4_11_0_clk a_29375_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2655 tdc0.w_dly_sig_n[123] tdc0.w_dly_sig[122] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2656 VPWR a_7378_13103# clknet_4_5_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2657 VPWR tdc0.w_dly_sig[62] tdc0.w_dly_sig_n[63] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2659 a_25155_3689# a_25026_3433# a_24735_3543# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2660 VGND a_30239_9839# a_30407_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2661 a_2401_9839# a_1867_9845# a_2306_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2663 tdc0.w_dly_sig[64] tdc0.w_dly_sig_n[62] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2664 VPWR a_4866_11989# a_4793_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2665 VGND a_4203_10927# a_4371_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2666 a_16737_9441# _036_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X2667 tdc0.w_dly_sig[106] tdc0.w_dly_sig_n[105] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2668 a_21327_3543# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2669 a_12134_15253# a_11966_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2670 VPWR tdc0.w_dly_sig[74] tdc0.w_dly_sig_n[75] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2671 tdc0.w_dly_sig_n[39] tdc0.w_dly_sig[39] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2672 VPWR _038_ a_19395_3543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2673 VGND tdc0.w_dly_sig[138] tdc0.w_dly_sig_n[139] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2674 VPWR tdc0.w_dly_sig[148] tdc0.w_dly_sig_n[148] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2675 a_9884_10217# a_9485_9845# a_9758_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2676 a_17996_8751# _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X2677 VGND a_26663_4631# tdc0.o_result[188] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2678 VPWR a_4387_4399# a_4555_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2679 VPWR a_24915_8983# _186_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2680 a_4387_4399# a_3689_4405# a_4130_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2681 a_30357_5865# a_29803_5705# a_30010_5764# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2682 VGND _105_ a_17231_8457# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X2683 uo_out[2] a_17937_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2684 VPWR a_23351_14423# _146_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2685 VGND tdc0.w_dly_sig_n[155] tdc0.w_dly_sig[156] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2686 VPWR tdc0.w_dly_sig[15] tdc0.w_dly_sig_n[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2687 a_25571_1653# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2688 VPWR tdc0.o_result[93] a_12539_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2690 a_11785_2229# a_11619_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2691 VPWR a_17010_17429# a_16937_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2692 VGND a_25663_14709# a_25670_15009# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2693 VPWR tdc0.w_dly_sig[33] tdc0.w_dly_sig_n[34] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2694 a_2474_9813# a_2306_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2695 VPWR tdc0.w_dly_sig[82] tdc0.w_dly_sig_n[83] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2696 net6 a_18151_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2697 VPWR a_14675_15253# a_14591_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2698 a_21081_14735# tdc0.w_dly_sig[67] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2699 VPWR a_12391_15279# a_12559_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2700 tdc0.w_dly_sig_n[186] tdc0.w_dly_sig[186] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2702 a_19767_10071# a_20051_10057# a_19986_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2703 VPWR tdc0.w_dly_sig[102] tdc0.w_dly_sig_n[103] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2704 a_12680_8457# _167_ a_12578_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X2705 tdc0.w_dly_sig_n[160] tdc0.w_dly_sig[160] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2706 a_26719_7119# a_26583_7093# a_26299_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2707 VGND a_23455_11145# a_23462_11049# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2708 a_25402_3311# a_25155_3689# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2709 a_18731_16367# a_17949_16373# a_18647_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2710 tdc0.w_dly_sig_n[189] tdc0.w_dly_sig[189] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2712 VPWR tdc0.o_result[66] a_21923_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2713 VPWR tdc0.o_result[134] a_12907_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2714 tdc0.w_dly_sig[138] tdc0.w_dly_sig_n[136] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2715 tdc0.w_dly_sig[129] tdc0.w_dly_sig_n[128] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2717 VPWR clknet_4_0_0_clk a_3247_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2718 VGND tdc0.w_dly_sig[30] tdc0.w_dly_sig_n[30] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2719 VGND tdc0.w_dly_sig[183] tdc0.w_dly_sig_n[183] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2720 tdc0.w_dly_sig_n[137] tdc0.w_dly_sig[137] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2721 VPWR a_14064_7093# _076_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2722 VGND a_27319_10057# a_27326_9961# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2723 VGND tdc0.w_dly_sig_n[161] tdc0.w_dly_sig[162] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2724 a_19211_7271# a_19307_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2725 VGND a_28883_13321# a_28890_13225# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2726 _001_ a_18059_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2728 a_23933_16367# tdc0.w_dly_sig[52] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2730 a_13580_6575# _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X2731 tdc0.w_dly_sig_n[153] tdc0.w_dly_sig[152] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2732 a_5985_15823# a_4995_15823# a_5859_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2733 VGND clknet_4_7_0_clk a_13643_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2734 VPWR a_17937_10927# uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2735 VGND net6 _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2736 a_1113_6031# a_947_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2737 VPWR a_16733_4917# _038_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.75 as=0.135 ps=1.27 w=1 l=0.15
X2738 VGND tdc0.w_dly_sig_n[83] tdc0.w_dly_sig[84] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2739 a_30124_9129# a_29725_8757# a_29998_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2740 tdc0.w_dly_sig[118] tdc0.w_dly_sig_n[116] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2741 a_30186_5487# a_29939_5865# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2742 VPWR a_13997_7637# _023_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2743 VPWR a_5050_8319# a_4977_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2744 VGND a_6476_6549# clknet_4_0_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2745 a_20499_13799# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2746 tdc0.w_dly_sig_n[67] tdc0.w_dly_sig[67] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2747 tdc0.w_dly_sig[44] tdc0.w_dly_sig_n[43] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2748 tdc0.w_dly_sig[151] tdc0.w_dly_sig_n[150] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2749 a_18217_9839# _114_ a_17967_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2750 VGND a_2715_11739# a_2673_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2751 tdc0.w_dly_sig_n[41] tdc0.w_dly_sig[40] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2752 VGND a_8803_2223# a_8971_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2753 VPWR tdc0.w_dly_sig[99] tdc0.w_dly_sig_n[100] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2754 a_30541_11305# a_29987_11145# a_30194_11204# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2755 a_18059_11721# _149_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2756 a_19066_2767# a_18751_2919# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2757 VGND a_11858_1109# a_11816_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2758 a_23947_12335# _170_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2759 a_25467_7119# a_25247_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2760 tdc0.w_dly_sig[90] tdc0.w_dly_sig_n[88] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2761 tdc0.w_dly_sig[80] tdc0.w_dly_sig_n[78] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2762 VPWR tdc0.w_dly_sig_n[76] tdc0.w_dly_sig[77] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2763 clknet_4_10_0_clk a_25428_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2764 VGND a_16127_4943# _060_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2765 VPWR tdc0.w_dly_sig_n[187] tdc0.w_dly_sig[188] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2766 _155_ a_13275_7776# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2767 VGND a_26767_16885# a_26774_17185# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2768 a_20525_1679# a_20359_1679# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2769 VPWR a_6430_5461# a_6357_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2770 a_2122_14013# a_1683_13647# a_2037_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2771 a_11230_2045# a_10791_1679# a_11145_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2772 VPWR ui_in[5] a_17634_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X2773 VGND a_3946_10901# a_3904_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2774 a_6476_6549# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2775 a_24731_14423# tdc0.o_result[51] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2776 VPWR tdc0.w_dly_sig_n[115] tdc0.w_dly_sig[116] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2778 VGND a_12226_2197# a_12184_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2779 VPWR tdc0.w_dly_sig[30] tdc0.w_dly_sig_n[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2780 VPWR a_16210_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2781 VPWR _003_ a_20499_13799# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2782 a_19855_8359# tdc0.o_result[29] a_20089_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2783 a_20292_9071# _010_ a_20172_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X2784 VGND tdc0.w_dly_sig_n[31] tdc0.w_dly_sig[33] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2785 VGND net3 _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X2786 a_1738_5461# a_1570_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2787 VGND a_21104_6005# clknet_4_8_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2790 VGND tdc0.w_dly_sig_n[128] tdc0.w_dly_sig[130] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2791 a_23240_13897# _004_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X2792 a_23193_7669# a_23027_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2793 a_27319_12233# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2794 VGND tdc0.w_dly_sig_n[156] tdc0.w_dly_sig[157] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2795 a_14563_9545# _080_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2796 a_20187_10217# a_20051_10057# a_19767_10071# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2797 VPWR ui_in[7] a_18151_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2798 VGND _051_ a_12325_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2799 VPWR tdc0.w_dly_sig_n[15] tdc0.w_dly_sig[17] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2801 VPWR a_7263_6005# a_7270_6305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2802 tdc0.w_dly_sig_n[182] tdc0.w_dly_sig[182] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2803 tdc0.w_dly_sig[140] tdc0.w_dly_sig_n[139] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2804 tdc0.w_dly_sig[16] tdc0.w_dly_sig_n[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2805 tdc0.w_dly_sig[60] tdc0.w_dly_sig_n[59] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2806 tdc0.w_dly_sig[162] tdc0.w_dly_sig_n[160] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2807 a_25375_8983# _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2808 tdc0.w_dly_sig[128] tdc0.w_dly_sig_n[127] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2809 a_17218_3855# _103_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X2810 a_10861_12559# a_9871_12559# a_10735_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2812 VPWR clknet_4_7_0_clk a_14747_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2814 tdc0.w_dly_sig[7] tdc0.w_dly_sig_n[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2815 VPWR a_9431_8475# a_9347_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2816 tdc0.w_dly_sig_n[12] tdc0.w_dly_sig[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2817 tdc0.w_dly_sig_n[48] tdc0.w_dly_sig[47] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2818 tdc0.w_dly_sig[32] tdc0.w_dly_sig_n[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2819 VPWR net5 a_15885_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X2820 VGND a_14437_8725# _117_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X2821 VPWR a_23903_5095# tdc0.o_result[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2822 tdc0.w_dly_sig_n[17] tdc0.w_dly_sig[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2823 VPWR a_13035_5487# a_13203_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2824 a_13035_5487# a_12337_5493# a_12778_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2825 a_14045_12353# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X2826 tdc0.w_dly_sig[138] tdc0.w_dly_sig_n[137] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2827 a_4222_3967# a_4054_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2828 a_24419_4943# a_24290_5217# a_23999_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2829 a_27455_10217# a_27326_9961# a_27035_10071# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2830 a_14379_7119# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2831 a_2589_7663# tdc0.w_dly_sig[116] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2832 a_11923_14191# a_11141_14197# a_11839_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2833 VPWR tdc0.w_dly_sig[134] tdc0.w_dly_sig_n[135] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2834 _089_ a_12526_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X2835 VPWR _001_ a_17187_13799# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2836 VGND tdc0.w_dly_sig_n[60] tdc0.w_dly_sig[62] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2837 VPWR tdc0.w_dly_sig_n[4] tdc0.w_dly_sig[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2838 a_26571_8359# a_26667_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2839 VPWR tdc0.w_dly_sig_n[96] tdc0.w_dly_sig[98] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2840 a_16658_15101# a_16385_14735# a_16573_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2841 a_24731_14423# tdc0.o_result[51] a_24965_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2842 tdc0.w_dly_sig_n[115] tdc0.w_dly_sig[115] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2843 VPWR a_18703_12559# _003_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R8 VGND uio_out[2] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2845 VPWR tdc0.w_dly_sig[111] tdc0.w_dly_sig_n[111] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2846 tdc0.o_result[68] a_20563_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2847 a_14721_11445# tdc0.o_result[82] a_14974_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X2848 a_19294_8457# _158_ a_18980_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X2849 tdc0.w_dly_sig_n[103] tdc0.w_dly_sig[103] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2850 tdc0.w_dly_sig_n[149] tdc0.w_dly_sig[148] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2851 VGND _007_ a_12693_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2852 VGND a_25295_8181# a_25302_8481# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2853 VPWR clknet_4_15_0_clk a_23579_16373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2854 a_7166_3285# a_6998_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2855 VPWR tdc0.w_dly_sig_n[104] tdc0.w_dly_sig[105] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2856 VGND _194_ a_20175_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2857 VPWR tdc0.o_result[78] a_13367_9952# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2858 VPWR a_25663_14709# a_25670_15009# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2859 VPWR a_11812_13621# clknet_4_7_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2860 tdc0.w_dly_sig[188] tdc0.w_dly_sig_n[187] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2861 VGND tdc0.w_dly_sig[92] tdc0.w_dly_sig_n[92] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2862 tdc0.w_dly_sig[153] tdc0.w_dly_sig_n[151] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2865 clknet_4_10_0_clk a_25428_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X2866 tdc0.w_dly_sig_n[88] tdc0.w_dly_sig[88] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2867 tdc0.w_dly_sig[165] tdc0.w_dly_sig_n[163] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2868 a_24149_1135# a_23811_1367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2869 a_13722_9295# tdc0.o_result[126] a_13641_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X2870 a_9347_16189# a_8565_15823# a_9263_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2871 a_12851_15101# a_11987_14735# a_12594_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2872 VGND tdc0.w_dly_sig_n[87] tdc0.w_dly_sig[88] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2873 VPWR _157_ a_13249_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2874 a_8470_3311# a_8197_3317# a_8385_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2875 VPWR a_22852_7093# clknet_4_9_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2876 tdc0.w_dly_sig[78] tdc0.w_dly_sig_n[77] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2877 a_10819_14013# a_10037_13647# a_10735_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2878 VGND a_16210_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2879 _120_ a_14103_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2880 VGND a_25288_10357# _638_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2881 a_17415_12015# _047_ a_17498_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X2882 clknet_4_11_0_clk a_26514_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2883 a_29621_16745# a_29067_16585# a_29274_16644# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2884 a_9577_2229# a_9411_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2885 VPWR a_11639_5211# a_11555_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2886 VGND net6 a_17703_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2887 a_13968_9545# _179_ a_13866_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X2888 VGND clknet_4_6_0_clk a_14931_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2889 tdc0.w_dly_sig[134] tdc0.w_dly_sig_n[133] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2890 a_23058_13897# _148_ a_22809_13793# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X2891 tdc0.w_dly_sig[124] tdc0.w_dly_sig_n[123] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2893 tdc0.w_dly_sig_n[150] tdc0.w_dly_sig[150] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2895 a_17695_6575# _001_ _064_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2896 VGND clknet_4_13_0_clk a_16219_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2897 tdc0.w_dly_sig_n[123] tdc0.w_dly_sig[123] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2898 VGND a_20074_6005# a_20003_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2899 a_8838_14013# a_8565_13647# a_8753_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2900 VGND tdc0.w_dly_sig_n[80] tdc0.w_dly_sig[81] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2901 VGND a_28883_12233# a_28890_12137# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2902 VGND a_30010_5764# a_29939_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2903 a_19899_3424# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2904 VPWR _026_ a_14379_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2905 a_9673_9839# tdc0.w_dly_sig[79] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2906 VPWR tdc0.w_dly_sig[126] tdc0.w_dly_sig_n[127] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2908 a_4314_17023# a_4146_17277# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2909 tdc0.w_dly_sig[133] tdc0.w_dly_sig_n[132] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2910 tdc0.w_dly_sig_n[91] tdc0.w_dly_sig[91] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2911 a_18659_7895# tdc0.o_result[18] a_18893_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2912 VGND tdc0.w_dly_sig[90] tdc0.w_dly_sig_n[90] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2913 a_16083_8235# _013_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2914 a_7423_3311# a_6725_3317# a_7166_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2915 VPWR tdc0.w_dly_sig[100] tdc0.w_dly_sig_n[101] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2916 a_25318_7093# a_25118_7393# a_25467_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2917 a_30124_8041# a_29725_7669# a_29998_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2918 VPWR a_11455_8475# a_11371_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2919 tdc0.o_result[138] a_10627_4123# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2920 VPWR a_26514_6575# clknet_4_11_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2921 a_7097_7119# tdc0.w_dly_sig[136] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2922 a_15094_16189# a_14655_15823# a_15009_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2923 VPWR a_15837_8181# _014_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2924 tdc0.w_dly_sig[97] tdc0.w_dly_sig_n[95] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2925 VPWR tdc0.w_dly_sig[152] tdc0.w_dly_sig_n[152] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2926 tdc0.o_result[132] a_5475_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2927 a_11356_1679# a_10957_1679# a_11230_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2928 a_15391_3855# _007_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2929 VPWR a_6503_4221# a_6671_4123# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2930 VGND tdc0.w_dly_sig[154] tdc0.w_dly_sig_n[155] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2931 a_16587_11721# _046_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2932 tdc0.w_dly_sig_n[6] tdc0.w_dly_sig[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2933 VGND a_2899_9813# a_2857_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2934 VPWR a_14805_6549# _080_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X2935 a_12693_3677# _025_ a_12621_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2936 a_17996_8751# _095_ a_17894_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X2938 tdc0.w_dly_sig_n[11] tdc0.w_dly_sig[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2939 a_23351_14423# tdc0.o_result[44] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2940 a_27399_4765# a_27179_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2941 a_14645_9545# _089_ a_14563_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2942 a_26217_14735# a_25670_15009# a_25870_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2943 a_29998_7663# a_29725_7669# a_29913_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2944 tdc0.w_dly_sig_n[135] tdc0.w_dly_sig[134] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2945 VPWR tdc0.w_dly_sig[97] tdc0.w_dly_sig_n[97] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2947 a_10129_17999# a_9963_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2948 a_14887_4631# _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2949 VGND clknet_4_5_0_clk a_8399_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2950 VPWR tdc0.w_dly_sig_n[111] tdc0.w_dly_sig[113] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2951 _077_ a_14379_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2952 a_5437_9661# a_4903_9295# a_5342_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2953 VGND tdc0.w_dly_sig_n[35] tdc0.w_dly_sig[36] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2954 VPWR tdc0.w_dly_sig_n[118] tdc0.w_dly_sig[119] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2955 VGND _050_ a_23420_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X2958 a_24547_1501# a_24327_1513# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2959 a_5817_11471# tdc0.o_result[118] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X2960 VPWR a_23155_10749# a_23323_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2961 VGND tdc0.w_dly_sig[136] tdc0.w_dly_sig_n[136] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2962 VGND tdc0.w_dly_sig_n[100] tdc0.w_dly_sig[101] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2963 VGND clknet_4_1_0_clk a_8859_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2964 a_20479_14191# a_19697_14197# a_20395_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2965 VGND _031_ a_17312_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X2966 a_13521_10205# _012_ a_13449_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2967 VGND a_3854_5461# a_3812_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2968 VGND a_1738_5461# a_1696_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2969 a_7699_15101# a_7001_14735# a_7442_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2970 a_13722_8207# _156_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X2971 a_28057_5865# a_27503_5705# a_27710_5764# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2972 a_7274_15101# a_6835_14735# a_7189_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2973 VGND clknet_4_1_0_clk a_6743_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2974 VGND tdc0.w_dly_sig[182] a_22721_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2975 clknet_4_6_0_clk a_12254_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2976 tdc0.w_dly_sig[152] tdc0.w_dly_sig_n[150] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2977 VGND tdc0.w_dly_sig[45] tdc0.w_dly_sig_n[46] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2978 a_25375_5095# a_25471_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2980 tdc0.w_dly_sig_n[118] tdc0.w_dly_sig[118] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2982 tdc0.w_dly_sig[166] tdc0.w_dly_sig_n[165] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2983 a_29423_5719# a_29519_5719# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2985 a_24009_11305# a_23462_11049# a_23662_11204# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2986 VGND a_16495_5487# _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2987 _064_ _001_ a_18479_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2988 clknet_4_0_0_clk a_6476_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X2989 VPWR a_22259_12533# a_22266_12833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2990 tdc0.w_dly_sig_n[7] tdc0.w_dly_sig[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2991 a_2033_9845# a_1867_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2992 a_26951_8181# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2993 tdc0.w_dly_sig[40] tdc0.w_dly_sig_n[39] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2994 tdc0.w_dly_sig[93] tdc0.w_dly_sig_n[92] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2995 a_26859_15497# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2996 a_15472_10159# tdc0.o_result[33] a_14897_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X2997 VPWR _051_ a_11711_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2998 tdc0.w_dly_sig_n[10] tdc0.w_dly_sig[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2999 VGND tdc0.w_dly_sig[70] tdc0.w_dly_sig_n[70] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3000 VGND a_20563_14165# a_20521_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3001 tdc0.w_dly_sig[17] tdc0.w_dly_sig_n[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3002 VGND a_26790_11445# a_26719_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3003 VGND tdc0.w_dly_sig[77] tdc0.w_dly_sig_n[78] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3004 VPWR a_7515_10749# a_7683_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3005 VGND tdc0.w_dly_sig[190] a_27597_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3006 VPWR a_17187_13799# _049_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3008 a_23351_14423# tdc0.o_result[44] a_23585_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3009 a_22546_957# a_22107_591# a_22461_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3010 tdc0.w_dly_sig_n[63] tdc0.w_dly_sig[63] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3011 VPWR tdc0.o_result[68] a_22291_14304# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3012 VPWR a_25428_7637# clknet_4_10_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3013 a_3873_7669# a_3707_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3014 tdc0.w_dly_sig_n[131] tdc0.w_dly_sig[131] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3015 a_25573_3689# a_25026_3433# a_25226_3588# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3016 tdc0.w_dly_sig[75] tdc0.w_dly_sig_n[73] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3017 a_27277_9839# a_26939_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3018 VGND tdc0.w_dly_sig[34] tdc0.w_dly_sig_n[34] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3019 a_17467_10357# _018_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X3022 a_6273_12015# _023_ a_6357_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3024 a_9485_9845# a_9319_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3025 clknet_4_6_0_clk a_12254_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R9 uio_oe[5] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3026 a_24954_3677# a_24639_3543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3027 VPWR _040_ a_20359_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3028 a_20039_13799# tdc0.o_result[43] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3030 tdc0.w_dly_sig_n[54] tdc0.w_dly_sig[53] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3031 a_11159_8864# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3032 VGND a_9263_16189# a_9431_16091# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3033 tdc0.o_result[106] a_2715_13915# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3034 VPWR clknet_4_2_0_clk a_10791_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3035 tdc0.o_result[121] a_5659_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3036 a_7369_3133# a_6835_2767# a_7274_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3037 VPWR a_24283_4917# a_24290_5217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3039 VPWR tdc0.w_dly_sig[74] tdc0.w_dly_sig_n[74] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3040 a_19057_591# tdc0.w_dly_sig[175] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3041 a_22641_957# a_22107_591# a_22546_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3042 VPWR tdc0.w_dly_sig_n[191] tdc0.w_dly_sig[192] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3043 VGND a_12007_7637# a_11965_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3045 a_30357_5865# a_29810_5609# a_30010_5764# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3046 tdc0.w_dly_sig_n[147] tdc0.w_dly_sig[146] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3047 VPWR tdc0.w_dly_sig[119] tdc0.w_dly_sig_n[119] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3049 a_22615_12559# a_22395_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3051 VGND tdc0.w_dly_sig[182] tdc0.w_dly_sig_n[183] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3052 VGND tdc0.w_dly_sig_n[161] tdc0.w_dly_sig[163] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3053 a_15731_7271# net6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X3054 VPWR a_3007_6575# a_3175_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3055 VPWR _003_ a_19289_13441# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3056 a_17194_2197# a_17026_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3057 VPWR clknet_4_13_0_clk a_16219_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3058 a_25665_7119# a_25111_7093# a_25318_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3059 tdc0.o_result[57] a_18171_18267# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3061 a_20359_11471# _063_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3062 a_25339_3855# a_25210_4129# a_24919_3829# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3063 a_9949_3855# tdc0.w_dly_sig[139] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3064 a_19802_6031# a_19487_6183# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3065 _190_ a_19163_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X3066 VGND tdc0.w_dly_sig_n[65] tdc0.w_dly_sig[66] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3067 tdc0.w_dly_sig_n[176] tdc0.w_dly_sig[176] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3068 VGND clknet_4_6_0_clk a_11895_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3069 VPWR tdc0.w_dly_sig_n[14] tdc0.w_dly_sig[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3071 a_24469_12015# tdc0.o_result[5] a_24659_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X3072 a_15094_16189# a_14821_15823# a_15009_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3073 a_22373_14557# tdc0.o_result[68] a_22291_14304# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3074 VGND a_11398_1791# a_11356_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3076 _032_ a_15483_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3077 a_5234_14847# a_5066_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3078 VPWR tdc0.w_dly_sig[167] tdc0.w_dly_sig_n[167] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3079 VGND a_24823_4007# tdc0.o_result[185] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3080 a_12552_15823# a_12153_15823# a_12426_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3081 a_3854_5461# a_3686_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3082 tdc0.w_dly_sig[23] tdc0.w_dly_sig_n[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3083 a_11605_1135# tdc0.w_dly_sig[167] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3084 VPWR clknet_4_5_0_clk a_3707_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3085 a_12241_2767# a_11251_2767# a_12115_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3086 tdc0.w_dly_sig[184] tdc0.w_dly_sig_n[182] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3087 a_14012_9839# tdc0.o_result[97] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X3088 a_20887_12809# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3089 tdc0.w_dly_sig[42] tdc0.w_dly_sig_n[41] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3090 a_19131_2741# clknet_4_8_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3091 a_24363_4007# tdc0.o_result[186] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3092 tdc0.w_dly_sig[70] tdc0.w_dly_sig_n[68] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3093 tdc0.w_dly_sig_n[185] tdc0.w_dly_sig[184] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3094 a_11329_6575# tdc0.w_dly_sig[140] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3095 a_19855_8359# tdc0.o_result[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3097 net1 a_30347_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3098 VGND tdc0.w_dly_sig[101] tdc0.w_dly_sig_n[101] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3099 VPWR a_26583_11445# a_26590_11745# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3100 VPWR tdc0.o_result[46] a_20848_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X3101 _083_ a_14379_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3102 tdc0.w_dly_sig[49] tdc0.w_dly_sig_n[48] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3103 a_15212_11471# _004_ a_14721_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3105 VPWR tdc0.w_dly_sig[113] tdc0.w_dly_sig_n[114] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3106 a_24334_8751# _187_ a_24254_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3107 a_11881_15279# tdc0.w_dly_sig[86] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3108 a_29437_13481# a_28890_13225# a_29090_13380# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3109 VPWR a_5659_15003# a_5575_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3110 a_25571_1653# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3112 tdc0.w_dly_sig[107] tdc0.w_dly_sig_n[106] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3113 tdc0.w_dly_sig_n[60] tdc0.w_dly_sig[60] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3114 VGND a_19954_15253# a_19912_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3115 a_24176_11471# _012_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X3117 VGND a_11471_5309# a_11639_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3118 a_4824_12393# a_4425_12021# a_4698_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3119 VPWR a_21327_17687# tdc0.o_result[54] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3120 VPWR a_29090_13380# a_29019_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3121 a_15496_12559# a_15097_12559# a_15370_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3122 VGND a_26882_12559# clknet_4_14_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3123 a_20204_9545# _175_ a_20102_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X3125 a_29987_11145# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3126 a_14917_2223# tdc0.w_dly_sig[169] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3127 VGND clknet_4_8_0_clk a_22107_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3128 a_24639_3543# a_24735_3543# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3129 a_14931_3855# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3130 tdc0.w_dly_sig_n[188] tdc0.w_dly_sig[187] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3131 VPWR clknet_4_1_0_clk a_8399_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3132 tdc0.w_dly_sig[122] tdc0.w_dly_sig_n[121] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3133 tdc0.w_dly_sig[2] tdc0.w_dly_sig_n[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3134 a_11141_7669# a_10975_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3135 tdc0.w_dly_sig[131] tdc0.w_dly_sig_n[130] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3137 a_11589_7119# _025_ a_11517_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3138 VPWR tdc0.w_dly_sig[23] a_25849_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3139 VPWR a_19773_9441# _177_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X3140 VGND a_22771_17179# a_22729_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3141 tdc0.w_dly_sig[143] tdc0.w_dly_sig_n[142] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3142 a_6261_11247# tdc0.o_result[100] a_5823_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3143 tdc0.w_dly_sig_n[141] tdc0.w_dly_sig[140] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3144 tdc0.w_dly_sig[48] tdc0.w_dly_sig_n[47] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3145 VPWR a_30347_10357# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3146 a_14082_18543# a_13643_18549# a_13997_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3147 tdc0.w_dly_sig[76] tdc0.w_dly_sig_n[75] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3148 tdc0.w_dly_sig[65] tdc0.w_dly_sig_n[64] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3149 a_23055_957# a_22273_591# a_22971_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3150 a_27179_4777# a_27043_4617# a_26759_4631# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3151 tdc0.w_dly_sig[147] tdc0.w_dly_sig_n[145] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3152 tdc0.w_dly_sig_n[148] tdc0.w_dly_sig[147] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3153 a_20421_11305# a_19867_11145# a_20074_11204# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3154 VGND tdc0.w_dly_sig_n[26] tdc0.w_dly_sig[28] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3155 VGND clknet_4_2_0_clk a_11619_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3156 _167_ a_11711_4512# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3157 _001_ a_18059_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3158 VGND a_6476_7637# clknet_4_1_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3159 a_5970_2879# a_5802_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3160 _206_ a_15575_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3161 VGND tdc0.w_dly_sig[168] tdc0.w_dly_sig_n[168] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3162 VPWR clknet_4_0_0_clk a_2051_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3163 tdc0.w_dly_sig_n[87] tdc0.w_dly_sig[86] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3164 a_23844_10159# tdc0.o_result[35] a_23269_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X3165 VGND a_16923_16885# a_16930_17185# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3166 a_13498_13103# _138_ a_13184_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X3167 a_24327_1513# a_24191_1353# a_23907_1367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3168 tdc0.w_dly_sig_n[98] tdc0.w_dly_sig[98] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3169 a_10635_17277# a_9853_16911# a_10551_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3170 VPWR tdc0.w_dly_sig_n[60] tdc0.w_dly_sig[61] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3171 VPWR a_8051_10901# a_7967_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3174 VPWR a_24823_4007# tdc0.o_result[185] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3175 a_8013_7669# a_7847_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3176 a_18847_2741# a_19131_2741# a_19066_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3177 VGND clknet_4_6_0_clk a_9963_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3178 VGND a_9006_8319# a_8964_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3180 VPWR tdc0.w_dly_sig_n[168] tdc0.w_dly_sig[170] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3181 VPWR tdc0.w_dly_sig_n[171] tdc0.w_dly_sig[172] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3182 a_29361_4943# net23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3183 VGND tdc0.w_dly_sig[84] tdc0.w_dly_sig_n[85] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3184 VPWR _064_ a_18127_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3185 a_13530_2223# a_13257_2229# a_13445_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3186 VGND tdc0.w_dly_sig[108] tdc0.w_dly_sig_n[108] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3188 tdc0.w_dly_sig_n[21] tdc0.w_dly_sig[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3189 a_14047_16367# a_13349_16373# a_13790_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3190 tdc0.w_dly_sig_n[65] tdc0.w_dly_sig[64] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3191 tdc0.o_result[145] a_6855_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3192 a_1297_7119# a_1131_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3193 _198_ a_12999_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3194 VPWR tdc0.w_dly_sig_n[156] tdc0.w_dly_sig[158] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3195 VPWR tdc0.w_dly_sig_n[103] tdc0.w_dly_sig[104] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3196 a_4479_4221# a_3615_3855# a_4222_3967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3197 VPWR a_18703_10383# _058_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3198 VPWR tdc0.w_dly_sig[54] a_24837_18921# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3199 VGND _040_ a_14441_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3200 tdc0.w_dly_sig[121] tdc0.w_dly_sig_n[119] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3201 a_29814_9839# a_29375_9845# a_29729_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3202 VGND a_11839_14191# a_12007_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3203 VPWR tdc0.w_dly_sig[72] tdc0.w_dly_sig_n[73] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3205 a_12877_6031# _060_ a_12805_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3206 VPWR _051_ a_11251_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3207 VGND tdc0.w_dly_sig[48] tdc0.w_dly_sig_n[49] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3208 VGND tdc0.w_dly_sig_n[97] tdc0.w_dly_sig[98] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3209 VPWR tdc0.w_dly_sig[27] tdc0.w_dly_sig_n[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3210 VGND a_10570_11583# a_10528_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3211 a_19629_6941# _010_ a_19557_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3212 tdc0.o_result[125] a_7867_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3213 a_9945_2223# a_9411_2229# a_9850_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3214 VGND tdc0.w_dly_sig[187] tdc0.w_dly_sig_n[187] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3215 VPWR tdc0.w_dly_sig_n[180] tdc0.w_dly_sig[181] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3216 tdc0.w_dly_sig[153] tdc0.w_dly_sig_n[152] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3217 VPWR a_4295_11837# a_4463_11739# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3219 VGND tdc0.o_result[59] a_17969_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X3220 VPWR tdc0.w_dly_sig[159] tdc0.w_dly_sig_n[159] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3221 _199_ a_12999_3424# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3222 VPWR clknet_4_3_0_clk a_10423_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3223 a_20887_12809# tdc0.o_result[7] a_20697_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X3224 a_21423_11159# a_21707_11145# a_21642_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3226 a_16109_10633# tdc0.o_result[76] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3227 VPWR a_20258_10116# a_20187_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3228 a_7825_2767# a_6835_2767# a_7699_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
R10 tt_um_hpretl_tt06_tdc_v1_18.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3229 tdc0.w_dly_sig[95] tdc0.w_dly_sig_n[93] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3230 VPWR _043_ a_13459_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3232 a_22787_15279# a_21923_15285# a_22530_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3233 VGND _076_ a_11957_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3234 _081_ a_15023_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3235 VGND _099_ a_14989_8353# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X3236 a_25410_3829# a_25203_3829# a_25586_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3237 _145_ a_18046_4719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X3238 tdc0.w_dly_sig[125] tdc0.w_dly_sig_n[124] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3239 VPWR a_19567_957# a_19735_859# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3240 tdc0.w_dly_sig_n[3] tdc0.w_dly_sig[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3241 VPWR tdc0.w_dly_sig_n[37] tdc0.w_dly_sig[39] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3242 a_29446_5309# a_29007_4943# a_29361_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3244 tdc0.w_dly_sig[68] tdc0.w_dly_sig_n[67] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3246 a_24893_14557# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X3247 a_8914_17429# a_8746_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3248 tdc0.w_dly_sig[84] tdc0.w_dly_sig_n[82] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3249 a_23271_6793# clknet_4_9_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3250 VGND a_22891_6807# tdc0.o_result[24] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3252 a_22457_15279# a_21923_15285# a_22362_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3253 a_19947_7119# a_19727_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3254 VGND tdc0.w_dly_sig[111] tdc0.w_dly_sig_n[112] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3255 a_19131_2741# clknet_4_8_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3256 tdc0.w_dly_sig_n[89] tdc0.w_dly_sig[89] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3259 VPWR a_17451_2223# a_17619_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3260 a_1738_7231# a_1570_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3261 tdc0.w_dly_sig_n[73] tdc0.w_dly_sig[73] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3262 VPWR a_20697_12809# uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3263 a_16757_17455# tdc0.w_dly_sig[59] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3264 a_1849_10927# a_1315_10933# a_1754_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3266 VGND a_11030_8319# a_10988_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3267 a_16293_18549# a_16127_18549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3268 tdc0.w_dly_sig[37] tdc0.w_dly_sig_n[36] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3269 VPWR a_11471_5309# a_11639_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3271 VGND tdc0.w_dly_sig_n[178] tdc0.w_dly_sig[180] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3272 VPWR a_22143_5487# a_22311_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3274 _014_ a_15837_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.38 ps=2.76 w=1 l=0.15
X3275 a_17765_13103# tdc0.o_result[40] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3276 a_22143_5487# a_21445_5493# a_21886_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3277 tdc0.w_dly_sig_n[63] tdc0.w_dly_sig[62] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3278 a_7166_3285# a_6998_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3279 a_9213_8751# tdc0.w_dly_sig[130] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3280 tdc0.w_dly_sig[172] tdc0.w_dly_sig_n[171] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3281 tdc0.w_dly_sig[175] tdc0.w_dly_sig_n[173] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3283 a_26571_8983# a_26667_8983# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3284 _086_ a_11803_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3285 VGND tdc0.w_dly_sig_n[152] tdc0.w_dly_sig[154] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3286 a_1485_5487# tdc0.w_dly_sig[150] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3287 VPWR tdc0.w_dly_sig[61] tdc0.w_dly_sig_n[62] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3288 a_3601_5487# tdc0.w_dly_sig[148] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3289 tdc0.o_result[56] a_17159_18517# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3290 VPWR a_21787_3543# _103_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3292 VGND tdc0.w_dly_sig[47] a_29621_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3294 VGND tdc0.w_dly_sig_n[113] tdc0.w_dly_sig[114] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3295 tdc0.w_dly_sig_n[75] tdc0.w_dly_sig[74] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3296 VGND tdc0.w_dly_sig[174] tdc0.w_dly_sig_n[174] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3297 a_11858_2879# a_11690_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3298 tdc0.o_result[56] a_17159_18517# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3299 a_6729_16367# tdc0.w_dly_sig[99] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3300 tdc0.o_result[166] a_12283_1109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3301 VGND tdc0.w_dly_sig_n[138] tdc0.w_dly_sig[139] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3302 clknet_4_1_0_clk a_6476_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3303 VPWR tdc0.w_dly_sig_n[157] tdc0.w_dly_sig[158] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3304 VGND tdc0.w_dly_sig_n[186] tdc0.w_dly_sig[187] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3305 tdc0.o_result[98] a_7407_16341# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3306 a_23535_17821# a_23315_17833# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3307 a_23903_4007# tdc0.o_result[179] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3308 a_11414_6397# a_11141_6031# a_11329_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3309 tdc0.w_dly_sig_n[76] tdc0.w_dly_sig[76] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3310 VPWR _004_ a_19881_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X3311 a_11141_6581# a_10975_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3312 a_27455_10217# a_27319_10057# a_27035_10071# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3313 tdc0.o_result[98] a_7407_16341# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3314 VPWR tdc0.w_dly_sig[83] tdc0.w_dly_sig_n[83] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3315 VPWR tdc0.w_dly_sig[116] tdc0.w_dly_sig_n[117] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3317 _138_ a_11711_13216# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3318 a_28057_5865# a_27510_5609# a_27710_5764# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3319 VPWR a_25410_13103# clknet_4_15_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3320 VPWR tdc0.w_dly_sig_n[0] tdc0.w_dly_sig[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3321 VGND a_10551_17277# a_10719_17179# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3322 a_18647_16367# a_17783_16373# a_18390_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3323 VPWR tdc0.w_dly_sig[160] tdc0.w_dly_sig_n[160] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3324 tdc0.w_dly_sig_n[68] tdc0.w_dly_sig[68] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3325 VGND _004_ a_19796_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X3326 a_27399_3855# a_27179_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3328 tdc0.o_result[96] a_9339_17429# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3329 VPWR tdc0.w_dly_sig_n[101] tdc0.w_dly_sig[102] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3331 tdc0.w_dly_sig[11] tdc0.w_dly_sig_n[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3332 VPWR tdc0.w_dly_sig[3] tdc0.w_dly_sig_n[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3333 a_23903_15975# a_23999_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3334 tdc0.o_result[96] a_9339_17429# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3335 VPWR a_19890_13103# clknet_4_13_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3336 a_17498_12015# _047_ a_17498_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X3338 _055_ a_20945_13675# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X3339 a_20966_1791# a_20798_2045# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3340 tdc0.w_dly_sig[96] tdc0.w_dly_sig_n[95] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3341 tdc0.w_dly_sig[105] tdc0.w_dly_sig_n[104] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3342 a_17152_14569# a_16753_14197# a_17026_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3343 _016_ a_19715_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X3344 VGND tdc0.w_dly_sig_n[100] tdc0.w_dly_sig[102] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3345 VGND a_12851_15101# a_13019_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3346 a_27035_12247# a_27326_12137# a_27277_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3347 tdc0.w_dly_sig_n[95] tdc0.w_dly_sig[95] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3348 a_25586_4221# a_25339_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3350 a_23947_12335# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3351 tdc0.o_result[82] a_10903_13915# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3352 tdc0.w_dly_sig_n[117] tdc0.w_dly_sig[117] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3353 tdc0.w_dly_sig[114] tdc0.w_dly_sig_n[112] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3354 tdc0.w_dly_sig[55] tdc0.w_dly_sig_n[54] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3356 _105_ a_17218_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X3357 clknet_4_5_0_clk a_7378_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3358 VGND a_27158_9028# a_27087_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3359 a_15737_16911# a_14747_16911# a_15611_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3360 VPWR a_21380_14165# clknet_4_12_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3362 VPWR tdc0.o_result[50] a_15420_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X3363 VGND tdc0.w_dly_sig[65] tdc0.w_dly_sig_n[66] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3364 VPWR tdc0.w_dly_sig_n[117] tdc0.w_dly_sig[119] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3365 VPWR _001_ a_21523_13799# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3366 VGND _170_ a_23947_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X3367 clknet_0_clk a_16210_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3368 VPWR tdc0.w_dly_sig[124] tdc0.w_dly_sig_n[125] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3369 tdc0.w_dly_sig[11] tdc0.w_dly_sig_n[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3370 VGND tdc0.w_dly_sig[73] tdc0.w_dly_sig_n[74] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3371 a_17075_18543# a_16293_18549# a_16991_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3372 VGND tdc0.w_dly_sig[43] tdc0.w_dly_sig_n[43] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3373 tdc0.w_dly_sig[191] tdc0.w_dly_sig_n[190] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3374 tdc0.w_dly_sig[65] tdc0.w_dly_sig_n[63] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3375 a_29572_4943# a_29173_4943# a_29446_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3376 a_16179_7637# a_16355_7969# a_16307_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X3377 VPWR tdc0.o_result[62] a_23855_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3378 VPWR a_13698_2197# a_13625_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3379 VGND tdc0.w_dly_sig_n[61] tdc0.w_dly_sig[63] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3380 a_18037_14735# tdc0.o_result[69] a_17691_14985# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3381 a_6177_13103# tdc0.w_dly_sig[123] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3382 a_12999_12128# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3383 a_23662_11204# a_23462_11049# a_23811_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3384 VPWR tdc0.w_dly_sig_n[132] tdc0.w_dly_sig[133] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3385 VGND tdc0.w_dly_sig_n[90] tdc0.w_dly_sig[91] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3387 a_15365_9545# _121_ a_15293_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3388 VGND tdc0.w_dly_sig_n[45] tdc0.w_dly_sig[47] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3389 VGND tdc0.w_dly_sig[127] tdc0.w_dly_sig_n[128] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3390 a_16713_8235# _021_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X3391 _179_ a_12815_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3392 tdc0.o_result[174] a_19735_859# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3393 a_19867_6005# clknet_4_9_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3395 a_11145_1679# tdc0.w_dly_sig[165] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3396 VPWR clknet_4_0_0_clk a_8031_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3397 VGND tdc0.w_dly_sig[56] tdc0.w_dly_sig_n[57] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3398 VPWR tdc0.w_dly_sig[1] a_25665_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3399 _171_ a_4995_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X3400 clknet_4_1_0_clk a_6476_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X3401 a_18222_16367# a_17949_16373# a_18137_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3403 VGND tdc0.w_dly_sig_n[185] tdc0.w_dly_sig[186] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3404 tdc0.w_dly_sig[13] tdc0.w_dly_sig_n[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3405 VGND a_22259_12533# a_22266_12833# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3406 VGND a_8638_3285# a_8596_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3407 tdc0.o_result[119] a_5291_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3408 a_5639_11471# _023_ a_5817_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X3410 VPWR tdc0.w_dly_sig_n[56] tdc0.w_dly_sig[58] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3411 a_5261_11247# _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X3413 a_5433_6031# a_4443_6031# a_5307_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3414 VGND _058_ a_13521_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3415 a_10827_18365# a_10129_17999# a_10570_18111# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3416 VPWR a_12191_18517# a_12107_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3417 VPWR _019_ a_17139_8759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3418 tdc0.o_result[119] a_5291_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3419 a_29519_5719# a_29810_5609# a_29761_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3420 clknet_4_4_0_clk a_6550_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3421 a_14499_3133# a_13717_2767# a_14415_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3422 VGND a_17159_18517# a_17117_18921# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3423 a_17777_13423# tdc0.o_result[88] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X3424 tdc0.w_dly_sig_n[42] tdc0.w_dly_sig[42] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3425 VGND ui_in[6] a_17507_1143# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3426 a_9255_17455# a_8473_17461# a_9171_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3428 VGND tdc0.w_dly_sig_n[99] tdc0.w_dly_sig[101] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3429 a_7442_2879# a_7274_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3430 tdc0.w_dly_sig_n[68] tdc0.w_dly_sig[67] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3431 tdc0.w_dly_sig[70] tdc0.w_dly_sig_n[69] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3432 VPWR a_19395_6807# _045_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3433 tdc0.w_dly_sig[180] tdc0.w_dly_sig_n[179] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3434 a_28687_16599# a_28783_16599# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3435 tdc0.w_dly_sig[34] tdc0.w_dly_sig_n[33] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3436 VGND _012_ a_20292_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X3438 a_15312_16911# a_14913_16911# a_15186_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3439 VGND net6 a_18196_5719# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X3440 tdc0.w_dly_sig[14] tdc0.w_dly_sig_n[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3441 VGND clknet_4_2_0_clk a_10791_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3442 tdc0.o_result[133] a_5199_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3443 a_25870_14709# a_25670_15009# a_26019_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3445 tdc0.w_dly_sig_n[54] tdc0.w_dly_sig[54] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3446 VPWR tdc0.w_dly_sig[60] tdc0.w_dly_sig_n[61] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3447 VPWR tdc0.w_dly_sig[65] a_17109_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3448 VPWR a_24490_15797# a_24419_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3450 tdc0.o_result[131] a_8879_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3451 tdc0.w_dly_sig[5] tdc0.w_dly_sig_n[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3452 tdc0.w_dly_sig_n[80] tdc0.w_dly_sig[79] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3453 a_15097_12559# a_14931_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3454 a_16665_5487# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3455 VGND tdc0.w_dly_sig_n[133] tdc0.w_dly_sig[135] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3456 VPWR tdc0.w_dly_sig[30] a_21985_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3457 VPWR _010_ a_24915_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3458 VGND tdc0.w_dly_sig[86] tdc0.w_dly_sig_n[86] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3459 VGND _052_ a_16850_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X3460 tdc0.w_dly_sig_n[111] tdc0.w_dly_sig[111] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3462 VPWR tdc0.w_dly_sig_n[51] tdc0.w_dly_sig[53] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3463 a_17109_15823# a_16555_15797# a_16762_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3464 VPWR a_22852_7093# clknet_4_9_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3465 a_18003_18365# a_17305_17999# a_17746_18111# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3466 VPWR a_26387_17063# tdc0.o_result[50] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3467 VGND a_30423_8751# a_30591_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3468 a_17451_2223# a_16587_2229# a_17194_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3469 a_27250_3829# a_27050_4129# a_27399_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3470 a_11509_14191# a_10975_14197# a_11414_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3471 tdc0.w_dly_sig_n[92] tdc0.w_dly_sig[92] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3472 a_14878_11721# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X3473 tdc0.o_result[114] a_5291_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3475 a_27342_7940# a_27135_7881# a_27518_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3476 a_18129_17999# a_17139_17999# a_18003_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3478 a_4333_15285# a_4167_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3479 a_25927_1679# a_25707_1679# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3480 VGND tdc0.w_dly_sig_n[139] tdc0.w_dly_sig[141] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3481 VPWR tdc0.w_dly_sig[37] tdc0.w_dly_sig_n[38] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3482 a_21166_15101# a_20727_14735# a_21081_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3483 clknet_4_7_0_clk a_11812_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3484 tdc0.w_dly_sig[158] tdc0.w_dly_sig_n[157] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3485 tdc0.w_dly_sig[156] tdc0.w_dly_sig_n[155] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3486 VGND tdc0.w_dly_sig_n[8] tdc0.w_dly_sig[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3487 a_25155_13647# a_25026_13921# a_24735_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3488 a_24241_3133# a_23903_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3489 a_10459_4221# a_9761_3855# a_10202_3967# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3490 VPWR a_4647_4123# a_4563_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3491 _638_.X a_25288_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3492 VPWR tdc0.w_dly_sig[131] tdc0.w_dly_sig_n[131] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3493 a_16025_9545# _031_ a_16109_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3495 VPWR tdc0.w_dly_sig[166] tdc0.w_dly_sig_n[166] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3496 VPWR tdc0.w_dly_sig_n[168] tdc0.w_dly_sig[169] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3497 VPWR tdc0.w_dly_sig[11] tdc0.w_dly_sig_n[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3498 a_1995_5487# a_1131_5493# a_1738_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3499 a_5207_12015# a_4425_12021# a_5123_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3500 tdc0.w_dly_sig[178] tdc0.w_dly_sig_n[176] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3501 a_6430_5461# a_6262_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3502 VPWR tdc0.w_dly_sig[53] a_23733_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3503 VGND _172_ a_19255_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3504 a_4698_8751# a_4259_8757# a_4613_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3505 a_3873_10927# a_3339_10933# a_3778_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3506 a_13625_2223# a_13091_2229# a_13530_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3507 VGND tdc0.w_dly_sig_n[183] tdc0.w_dly_sig[185] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3508 a_23082_8725# a_22914_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3509 tdc0.w_dly_sig_n[158] tdc0.w_dly_sig[158] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3510 a_13809_15285# a_13643_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3511 VGND a_10506_7119# clknet_4_3_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X3512 tdc0.w_dly_sig[183] tdc0.w_dly_sig_n[181] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3513 a_6430_4373# a_6262_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3514 a_4088_4777# a_3689_4405# a_3962_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3515 a_6821_15279# tdc0.w_dly_sig[102] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3516 tdc0.w_dly_sig[193] tdc0.w_dly_sig_n[191] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3517 VGND tdc0.w_dly_sig[69] tdc0.w_dly_sig_n[69] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3518 a_6998_14191# a_6725_14197# a_6913_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3519 VPWR tdc0.w_dly_sig[178] tdc0.w_dly_sig_n[178] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3520 _029_ a_17599_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X3521 uo_out[6] a_19777_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3522 VPWR clknet_4_8_0_clk a_16127_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3523 VPWR tdc0.w_dly_sig_n[181] tdc0.w_dly_sig[182] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3525 a_25149_9117# _010_ a_25077_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3526 a_26974_16885# a_26774_17185# a_27123_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3527 VPWR tdc0.w_dly_sig[161] tdc0.w_dly_sig_n[161] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3528 VGND a_22714_703# a_22672_591# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3529 VPWR tdc0.w_dly_sig[33] tdc0.w_dly_sig_n[33] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3532 VGND a_18151_1135# net6 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3533 a_22445_14557# _001_ a_22373_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3534 VGND a_29614_5055# a_29572_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3535 VGND a_27342_7940# a_27271_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3536 VGND a_6550_12559# clknet_4_4_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X3538 a_3394_14165# a_3226_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3539 tdc0.o_result[45] a_30591_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3540 a_14361_10933# a_14195_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3541 a_4882_6397# a_4609_6031# a_4797_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3542 VGND a_4923_3035# a_4881_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3543 VPWR _012_ a_16205_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3544 a_29725_15285# a_29559_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3545 a_1849_12559# a_1683_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3546 a_23229_6575# a_22891_6807# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3547 tdc0.o_result[45] a_30591_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3548 VPWR clknet_4_11_0_clk a_29559_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3549 a_24241_18543# a_23903_18775# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3551 VPWR tdc0.w_dly_sig[127] tdc0.w_dly_sig_n[128] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3553 VGND _019_ a_16799_8235# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3554 VGND clknet_4_1_0_clk a_8399_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3555 a_23155_10749# a_22457_10383# a_22898_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3556 a_22261_11305# a_21714_11049# a_21914_11204# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3557 _011_ a_16495_5487# a_17023_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3558 VPWR tdc0.w_dly_sig_n[62] tdc0.w_dly_sig[63] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3559 VPWR a_24469_12015# uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3560 a_20407_10205# a_20187_10217# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3561 a_19255_12335# _174_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3562 VGND tdc0.o_result[34] a_15212_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X3563 a_1849_13109# a_1683_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3564 a_9834_4373# a_9666_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3566 VPWR a_14151_10535# _074_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3567 a_3689_4405# a_3523_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3568 VPWR _030_ a_19395_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3569 tdc0.w_dly_sig_n[173] tdc0.w_dly_sig[173] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3570 VPWR a_7423_3311# a_7591_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3571 VPWR tdc0.w_dly_sig[121] tdc0.w_dly_sig_n[122] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3573 VPWR a_27250_4676# a_27179_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3574 _010_ a_17691_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3575 a_23082_8725# a_22914_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3576 a_12226_2197# a_12058_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3578 a_24183_15511# tdc0.o_result[41] a_24309_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X3579 VGND _136_ a_19497_5089# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X3580 VGND tdc0.w_dly_sig[39] a_26309_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3581 VGND tdc0.w_dly_sig_n[189] tdc0.w_dly_sig[190] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3582 VGND a_27871_2741# a_27878_3041# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3583 VGND a_10091_4399# a_10259_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3584 a_25891_12559# a_25755_12533# a_25471_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3585 tdc0.w_dly_sig[89] tdc0.w_dly_sig_n[88] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3586 VPWR tdc0.w_dly_sig[75] tdc0.w_dly_sig_n[76] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3587 VGND _152_ a_23947_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3589 VPWR a_24398_1412# a_24327_1513# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3590 a_26794_15645# a_26479_15511# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3591 VGND tdc0.w_dly_sig[38] tdc0.w_dly_sig_n[38] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3592 tdc0.w_dly_sig_n[158] tdc0.w_dly_sig[157] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3593 tdc0.w_dly_sig[169] tdc0.w_dly_sig_n[168] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3594 VGND tdc0.w_dly_sig_n[167] tdc0.w_dly_sig[169] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3595 tdc0.o_result[160] a_9063_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3596 tdc0.w_dly_sig_n[56] tdc0.w_dly_sig[55] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3597 a_28841_13103# a_28503_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3598 VGND a_12007_6299# a_11965_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3599 a_2677_6575# a_2143_6581# a_2582_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3600 a_5805_11721# tdc0.o_result[102] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3601 a_14182_10159# tdc0.o_result[97] a_14101_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X3602 a_14274_13423# _120_ a_14520_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X3603 VGND _016_ a_20359_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3604 VPWR a_11582_6143# a_11509_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3605 VGND _009_ a_17323_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3606 tdc0.w_dly_sig_n[70] tdc0.w_dly_sig[70] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3607 a_27794_13103# a_27547_13481# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3608 a_1297_7119# a_1131_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3609 tdc0.w_dly_sig[182] tdc0.w_dly_sig_n[181] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3610 a_24443_16367# a_23745_16373# a_24186_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3611 clknet_4_6_0_clk a_12254_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3612 a_19255_12015# _172_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3613 tdc0.w_dly_sig_n[161] tdc0.w_dly_sig[161] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3614 _039_ a_15333_4737# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X3615 net25 a_29099_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3616 a_23627_6941# a_23407_6953# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3617 VGND tdc0.w_dly_sig_n[40] tdc0.w_dly_sig[42] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3618 a_19415_11721# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3619 tdc0.w_dly_sig_n[34] tdc0.w_dly_sig[34] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3620 VPWR tdc0.w_dly_sig[179] tdc0.w_dly_sig_n[180] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3621 a_27597_3855# a_27043_3829# a_27250_3829# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3622 VGND tdc0.w_dly_sig_n[27] tdc0.w_dly_sig[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3623 a_21039_3133# a_20175_2767# a_20782_2879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3624 VGND tdc0.w_dly_sig_n[25] tdc0.w_dly_sig[26] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3625 _148_ a_22291_14304# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3626 VPWR tdc0.w_dly_sig_n[163] tdc0.w_dly_sig[164] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3627 a_16560_6935# net4 a_16488_6935# VGND sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X3628 VPWR tdc0.w_dly_sig_n[58] tdc0.w_dly_sig[60] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3629 a_6357_12015# tdc0.o_result[119] a_6273_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3630 a_19629_8029# _030_ a_19557_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3631 a_14533_8207# _025_ a_14461_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3632 a_19969_18921# a_18979_18549# a_19843_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3633 VGND a_30407_12827# a_30365_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3634 a_30507_15279# a_29725_15285# a_30423_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3635 VPWR tdc0.w_dly_sig_n[126] tdc0.w_dly_sig[128] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3636 VGND tdc0.w_dly_sig[72] tdc0.w_dly_sig_n[72] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3637 a_25778_1653# a_25578_1953# a_25927_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3638 VPWR _018_ a_17567_9447# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3639 a_16826_14847# a_16658_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3640 VGND clknet_4_3_0_clk a_10423_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3642 a_24170_11721# tdc0.o_result[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X3643 VPWR a_3946_10901# a_3873_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3644 VPWR a_11260_5461# clknet_4_2_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3645 VPWR a_5491_15101# a_5659_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3646 VGND tdc0.w_dly_sig[184] a_24837_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3648 VGND a_7867_3035# a_7825_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3649 a_19928_5193# _135_ a_19826_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X3650 a_8454_7637# a_8286_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3651 VPWR clknet_4_15_0_clk a_29559_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3652 a_22714_703# a_22546_957# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3653 tdc0.w_dly_sig[141] tdc0.w_dly_sig_n[140] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3654 a_25757_3855# a_25210_4129# a_25410_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3655 a_19505_12015# _190_ a_19777_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3656 tdc0.w_dly_sig[18] tdc0.w_dly_sig_n[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3657 a_14326_9839# _073_ a_14012_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X3659 VPWR a_29515_4631# tdc0.o_result[191] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3660 tdc0.w_dly_sig[27] tdc0.w_dly_sig_n[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3661 VPWR tdc0.w_dly_sig[32] tdc0.w_dly_sig_n[33] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3662 VPWR tdc0.w_dly_sig[91] tdc0.w_dly_sig_n[92] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3663 tdc0.w_dly_sig[43] tdc0.w_dly_sig_n[42] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3664 a_20359_11471# _029_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3665 a_21051_8359# a_21147_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3666 a_4824_9129# a_4425_8757# a_4698_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3667 VPWR _017_ a_24113_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X3669 VGND a_23179_17673# a_23186_17577# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3670 VGND tdc0.w_dly_sig[52] tdc0.w_dly_sig_n[53] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3671 VPWR tdc0.w_dly_sig_n[19] tdc0.w_dly_sig[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3672 VGND _071_ a_24131_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3673 a_2474_9813# a_2306_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3674 VGND a_14675_15253# a_14633_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3675 a_6430_4373# a_6262_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3676 VGND a_6430_5461# a_6388_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3677 clknet_4_0_0_clk a_6476_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3679 tdc0.w_dly_sig[66] tdc0.w_dly_sig_n[65] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3680 tdc0.w_dly_sig_n[172] tdc0.w_dly_sig[172] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3681 VPWR _050_ a_17875_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3682 tdc0.w_dly_sig[104] tdc0.w_dly_sig_n[103] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3683 VGND tdc0.w_dly_sig[57] tdc0.w_dly_sig_n[57] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3684 a_19701_15279# tdc0.w_dly_sig[66] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3686 a_26939_7119# a_26719_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3687 VGND tdc0.w_dly_sig[163] tdc0.w_dly_sig_n[163] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3688 a_21603_4007# tdc0.o_result[182] a_21837_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3690 a_7423_3311# a_6559_3317# a_7166_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3691 a_24965_14557# _003_ a_24893_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3692 VPWR tdc0.w_dly_sig_n[186] tdc0.w_dly_sig[188] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3693 a_20417_4373# _182_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X3694 VPWR _039_ a_14104_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X3695 tdc0.w_dly_sig_n[52] tdc0.w_dly_sig[51] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3696 VGND tdc0.w_dly_sig[87] tdc0.w_dly_sig_n[87] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3697 tdc0.o_result[44] a_30591_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3698 VPWR clknet_0_clk a_6476_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3699 VPWR clknet_4_2_0_clk a_13091_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3700 a_4272_16911# a_3873_16911# a_4146_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3701 a_21923_13647# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3702 clknet_4_9_0_clk a_22852_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3703 a_7952_12393# a_7553_12021# a_7826_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3705 VPWR tdc0.w_dly_sig[68] tdc0.w_dly_sig_n[69] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3706 VPWR a_23339_8751# a_23507_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3707 VGND a_13698_2197# a_13656_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3708 VPWR tdc0.w_dly_sig[145] tdc0.w_dly_sig_n[145] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3709 VPWR tdc0.w_dly_sig_n[129] tdc0.w_dly_sig[131] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3710 a_5893_9295# a_4903_9295# a_5767_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3711 a_18869_591# a_18703_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3712 a_12337_5493# a_12171_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3713 tdc0.w_dly_sig[164] tdc0.w_dly_sig_n[163] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3714 a_6687_4399# a_5989_4405# a_6430_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3715 a_17695_6575# net6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3716 VGND a_17567_9447# _020_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3717 a_17117_591# a_16127_591# a_16991_957# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3718 VGND tdc0.w_dly_sig_n[157] tdc0.w_dly_sig[159] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3719 tdc0.w_dly_sig[93] tdc0.w_dly_sig_n[91] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3720 VGND a_26882_12559# clknet_4_14_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3722 a_6078_4221# a_5805_3855# a_5993_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3723 VPWR a_27526_10116# a_27455_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3724 VGND tdc0.w_dly_sig_n[7] tdc0.w_dly_sig[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3725 VPWR tdc0.w_dly_sig[180] tdc0.w_dly_sig_n[181] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3726 VGND tdc0.w_dly_sig[25] tdc0.w_dly_sig_n[26] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3727 VGND a_22679_4373# a_22637_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3728 VGND tdc0.w_dly_sig_n[23] tdc0.w_dly_sig[25] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3729 a_8385_3311# tdc0.w_dly_sig[161] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3730 uo_out[4] a_19225_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3732 VGND a_5475_6299# a_5433_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3733 tdc0.w_dly_sig[73] tdc0.w_dly_sig_n[71] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3734 tdc0.o_result[66] a_21759_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3735 a_27618_13380# a_27411_13321# a_27794_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3736 a_13392_4719# _025_ a_13272_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X3737 a_25247_7119# a_25118_7393# a_24827_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3738 a_22461_13103# tdc0.w_dly_sig[37] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3739 tdc0.o_result[80] a_10995_11739# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3740 a_14243_8001# _013_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X3741 VPWR a_27871_2741# a_27878_3041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3742 VGND a_23913_8353# _109_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X3744 VGND tdc0.w_dly_sig_n[172] tdc0.w_dly_sig[173] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3745 VGND tdc0.w_dly_sig[13] tdc0.w_dly_sig_n[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3746 VPWR _058_ a_21923_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3747 VGND tdc0.w_dly_sig[3] a_24009_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3748 VGND clknet_4_2_0_clk a_9595_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3749 tdc0.o_result[90] a_14675_17429# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3750 tdc0.w_dly_sig[126] tdc0.w_dly_sig_n[124] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3751 tdc0.w_dly_sig_n[35] tdc0.w_dly_sig[34] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3753 tdc0.w_dly_sig[20] tdc0.w_dly_sig_n[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3754 VGND a_26215_9269# a_26222_9569# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3755 a_25835_9447# a_25931_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3756 tdc0.w_dly_sig[44] tdc0.w_dly_sig_n[42] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3757 VPWR tdc0.o_result[81] a_11803_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3758 tdc0.w_dly_sig[26] tdc0.w_dly_sig_n[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3759 VGND a_24731_7271# tdc0.o_result[21] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3760 a_4774_7231# a_4606_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3761 tdc0.w_dly_sig_n[0] net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3762 a_27547_13481# a_27411_13321# a_27127_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3763 VGND tdc0.w_dly_sig_n[6] tdc0.w_dly_sig[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3764 a_13177_8867# _165_ a_13081_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3765 VGND tdc0.w_dly_sig_n[18] tdc0.w_dly_sig[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3766 a_12502_9813# a_12334_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3767 a_4774_7231# a_4606_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3768 VGND tdc0.w_dly_sig[100] tdc0.w_dly_sig_n[100] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3769 a_20072_4943# tdc0.o_result[188] a_19497_5089# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X3770 VGND tdc0.w_dly_sig[192] a_30449_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3771 tdc0.w_dly_sig_n[31] tdc0.w_dly_sig[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3772 tdc0.w_dly_sig[77] tdc0.w_dly_sig_n[75] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3773 VPWR net3 a_15013_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3774 VGND net6 a_17703_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3775 VPWR a_15611_17277# a_15779_17179# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3776 a_25690_4943# a_25375_5095# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3777 VGND _160_ a_19150_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X3778 VPWR a_3819_3285# a_3735_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3779 tdc0.w_dly_sig_n[173] tdc0.w_dly_sig[172] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3780 a_26203_7271# a_26299_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3781 VPWR a_24653_9545# uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3782 a_9758_9839# a_9485_9845# a_9673_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3783 a_7274_15101# a_7001_14735# a_7189_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3784 tdc0.w_dly_sig[148] tdc0.w_dly_sig_n[147] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3786 _144_ a_17875_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3787 VGND tdc0.w_dly_sig_n[85] tdc0.w_dly_sig[86] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3788 a_19142_957# a_18869_591# a_19057_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3789 VPWR a_20039_13799# _118_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3790 a_18703_11471# _150_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3792 tdc0.w_dly_sig[48] tdc0.w_dly_sig_n[46] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3793 a_2631_12925# a_1849_12559# a_2547_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3794 VPWR tdc0.w_dly_sig_n[175] tdc0.w_dly_sig[176] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3795 VGND a_25428_7637# clknet_4_10_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3796 VGND a_12999_8867# _170_ VGND sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X3797 tdc0.w_dly_sig_n[85] tdc0.w_dly_sig[84] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3798 VGND tdc0.w_dly_sig[143] tdc0.w_dly_sig_n[144] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3799 VGND tdc0.w_dly_sig[14] tdc0.w_dly_sig_n[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3800 a_30507_14191# a_29725_14197# a_30423_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3801 VPWR a_9558_7231# a_9485_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3802 clknet_4_15_0_clk a_25410_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3803 VPWR tdc0.w_dly_sig[184] tdc0.w_dly_sig_n[184] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3804 a_16733_4917# a_16999_4917# a_16945_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3805 VGND a_26514_6575# clknet_4_11_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3806 VPWR a_18171_18267# a_18087_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3807 a_3854_5461# a_3686_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3808 _125_ a_12618_7983# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X3809 VPWR tdc0.w_dly_sig_n[131] tdc0.w_dly_sig[133] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3810 a_30323_12925# a_29541_12559# a_30239_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3811 a_8596_16745# a_8197_16373# a_8470_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3812 VPWR a_6550_12559# clknet_4_4_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3813 VGND a_15963_12827# a_15921_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3814 a_24018_16367# a_23745_16373# a_23933_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3815 a_15477_12335# tdc0.o_result[38] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X3816 VPWR tdc0.w_dly_sig[144] tdc0.w_dly_sig_n[144] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3817 a_29817_6031# a_29651_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3818 VGND a_17251_15003# a_17209_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3819 VPWR a_7699_15101# a_7867_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3820 a_4295_11837# a_3597_11471# a_4038_11583# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3821 _104_ a_17047_3424# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3822 tdc0.w_dly_sig_n[96] tdc0.w_dly_sig[95] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3824 VGND tdc0.w_dly_sig_n[32] tdc0.w_dly_sig[34] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3825 a_12153_15823# a_11987_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3827 VGND a_17559_12711# _112_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X3828 tdc0.o_result[143] a_8327_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3829 tdc0.o_result[152] a_3083_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3830 a_24162_8457# _108_ a_23913_8353# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X3831 clknet_4_11_0_clk a_26514_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3832 a_14591_17455# a_13809_17461# a_14507_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3833 VPWR _058_ a_16495_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3834 _098_ a_14103_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3835 a_23407_6953# a_23271_6793# a_22987_6807# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3836 a_24126_1501# a_23811_1367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3838 tdc0.w_dly_sig_n[159] tdc0.w_dly_sig[158] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3839 VPWR a_24731_14423# _127_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3840 VGND a_10478_13759# a_10436_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3841 a_5123_8751# a_4425_8757# a_4866_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3843 VGND a_19183_2197# a_19141_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3844 a_30641_6031# a_29651_6031# a_30515_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3845 VGND a_27031_13335# tdc0.o_result[40] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3847 a_16762_15797# a_16555_15797# a_16938_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3848 a_10402_11837# a_10129_11471# a_10317_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3849 a_27031_13335# a_27127_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3850 a_29361_4943# net23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3851 a_13600_13103# _139_ a_13498_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X3852 VPWR tdc0.w_dly_sig[163] tdc0.w_dly_sig_n[164] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3853 VPWR _043_ a_14103_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3854 tdc0.w_dly_sig_n[112] tdc0.w_dly_sig[111] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3855 a_10126_17277# a_9853_16911# a_10041_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3856 tdc0.w_dly_sig_n[25] tdc0.w_dly_sig[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3858 tdc0.w_dly_sig_n[24] tdc0.w_dly_sig[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3859 a_22090_17455# a_21843_17833# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3860 VGND a_9431_13915# a_9389_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3861 a_5307_8573# a_4609_8207# a_5050_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3862 VPWR tdc0.w_dly_sig[180] tdc0.w_dly_sig_n[180] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3863 a_25665_11471# a_25111_11445# a_25318_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3864 tdc0.w_dly_sig[139] tdc0.w_dly_sig_n[138] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3865 VGND a_16495_5487# _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3866 VPWR clknet_4_13_0_clk a_16127_18549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3867 a_15097_12559# a_14931_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3868 VGND _054_ a_13889_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3869 a_17599_13103# _020_ a_17777_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X3870 VGND a_14983_7093# _007_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3871 a_5192_14735# a_4793_14735# a_5066_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3872 tdc0.w_dly_sig[89] tdc0.w_dly_sig_n[87] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3873 a_15121_4765# _005_ a_15049_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3874 VPWR a_15687_16091# a_15603_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3875 VPWR tdc0.w_dly_sig[107] tdc0.w_dly_sig_n[107] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3876 a_26851_7895# a_27142_7785# a_27093_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3877 VPWR tdc0.w_dly_sig[98] tdc0.w_dly_sig_n[99] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3878 a_30123_11471# a_29994_11745# a_29703_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3879 VPWR tdc0.w_dly_sig[187] a_25573_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3880 VPWR tdc0.w_dly_sig[46] tdc0.w_dly_sig_n[47] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3881 VPWR tdc0.w_dly_sig[7] tdc0.w_dly_sig_n[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3882 a_10034_3133# a_9595_2767# a_9949_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3883 VPWR a_16991_18543# a_17159_18517# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3885 VGND tdc0.w_dly_sig[130] tdc0.w_dly_sig_n[130] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3886 a_25471_4917# a_25762_5217# a_25713_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3887 tdc0.w_dly_sig_n[126] tdc0.w_dly_sig[126] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3888 VGND a_24639_13799# tdc0.o_result[39] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3889 VPWR tdc0.w_dly_sig_n[91] tdc0.w_dly_sig[92] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3890 tdc0.o_result[169] a_14123_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3891 VGND tdc0.w_dly_sig_n[142] tdc0.w_dly_sig[144] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3892 a_7994_11989# a_7826_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3893 VGND a_6476_6549# clknet_4_0_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3894 a_24419_4943# a_24283_4917# a_23999_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3895 VPWR clknet_4_2_0_clk a_9595_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3896 tdc0.w_dly_sig_n[102] tdc0.w_dly_sig[102] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3897 VPWR a_7239_16367# a_7407_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3898 tdc0.w_dly_sig_n[42] tdc0.w_dly_sig[41] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3900 _022_ a_16547_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3901 a_16845_10927# tdc0.o_result[146] a_16761_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3902 VGND _055_ a_19049_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3904 a_5510_9407# a_5342_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3905 a_17130_16885# a_16930_17185# a_17279_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3906 VGND tdc0.w_dly_sig[104] tdc0.w_dly_sig_n[105] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3907 a_26575_15511# a_26859_15497# a_26794_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3909 a_10570_11583# a_10402_11837# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3910 a_9485_7485# a_8951_7119# a_9390_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3911 VGND a_7239_16367# a_7407_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3912 VPWR tdc0.o_result[86] a_14839_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X3913 VGND a_2290_13077# a_2248_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3914 VPWR a_21207_3035# a_21123_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3916 VPWR clknet_4_0_0_clk a_947_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3917 VPWR a_14215_16341# a_14131_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3918 tdc0.w_dly_sig_n[83] tdc0.w_dly_sig[83] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3919 VGND _015_ a_19715_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3920 VPWR net24 a_30357_5865# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3921 clknet_4_10_0_clk a_25428_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3922 VGND clknet_4_7_0_clk a_11159_18549# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3923 VGND tdc0.w_dly_sig[129] tdc0.w_dly_sig_n[130] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3926 a_17681_13103# _028_ a_17599_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3927 tdc0.w_dly_sig_n[154] tdc0.w_dly_sig[153] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3928 VPWR a_19890_13103# clknet_4_13_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3929 VPWR tdc0.w_dly_sig_n[12] tdc0.w_dly_sig[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3930 VPWR _023_ a_13552_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X3931 VPWR a_9171_17455# a_9339_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3932 a_2309_6581# a_2143_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3933 tdc0.w_dly_sig_n[4] tdc0.w_dly_sig[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3934 VGND a_15609_4971# _008_ VGND sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X3935 a_20315_7895# tdc0.o_result[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3936 VGND tdc0.w_dly_sig[93] tdc0.w_dly_sig_n[93] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3937 tdc0.w_dly_sig[79] tdc0.w_dly_sig_n[78] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3938 a_3643_15279# a_2861_15285# a_3559_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3939 a_2547_13103# a_1849_13109# a_2290_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3940 VPWR a_19289_13441# _017_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X3941 tdc0.w_dly_sig_n[187] tdc0.w_dly_sig[186] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3942 VGND a_21104_6005# clknet_4_8_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3943 tdc0.w_dly_sig[161] tdc0.w_dly_sig_n[159] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3944 tdc0.w_dly_sig[163] tdc0.w_dly_sig_n[162] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3945 tdc0.w_dly_sig[28] tdc0.w_dly_sig_n[26] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3947 a_24191_1353# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3948 _150_ a_18059_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X3949 VPWR _000_ a_18059_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3950 a_1849_12559# a_1683_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3952 VGND a_11766_18517# a_11724_18921# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3953 tdc0.w_dly_sig[102] tdc0.w_dly_sig_n[100] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3954 VPWR tdc0.w_dly_sig[49] a_26309_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3955 a_19813_5853# _030_ a_19741_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3956 VGND clknet_4_7_0_clk a_13183_16373# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3957 a_5805_3855# a_5639_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3958 VPWR a_11839_6397# a_12007_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3959 VGND _154_ a_23947_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3960 tdc0.w_dly_sig_n[129] tdc0.w_dly_sig[128] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3961 VGND a_17565_8725# _097_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X3962 VPWR a_5115_11159# _131_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X3963 a_24639_2767# a_24419_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3964 VPWR tdc0.o_result[35] a_23700_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X3965 tdc0.w_dly_sig[23] tdc0.w_dly_sig_n[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3966 _064_ _001_ a_18479_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3967 _010_ a_17691_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X3969 a_27342_7940# a_27142_7785# a_27491_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3971 VGND tdc0.w_dly_sig_n[127] tdc0.w_dly_sig[129] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3972 tdc0.w_dly_sig[22] tdc0.w_dly_sig_n[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3973 VPWR a_17923_5719# _019_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3974 VGND tdc0.w_dly_sig_n[9] tdc0.w_dly_sig[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3975 a_26309_15823# a_25755_15797# a_25962_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3976 a_7185_10933# a_7019_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3977 a_16577_12559# tdc0.o_result[72] a_16495_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3978 a_21523_13799# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X3979 a_12391_15279# a_11693_15285# a_12134_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3980 _100_ a_14563_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3981 a_2121_7119# a_1131_7119# a_1995_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3982 tdc0.w_dly_sig_n[125] tdc0.w_dly_sig[124] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3983 tdc0.w_dly_sig_n[74] tdc0.w_dly_sig[73] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3984 VGND tdc0.w_dly_sig_n[36] tdc0.w_dly_sig[38] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3985 tdc0.o_result[127] a_8419_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3987 a_11923_6575# a_11141_6581# a_11839_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3988 VGND tdc0.w_dly_sig_n[28] tdc0.w_dly_sig[30] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3989 tdc0.w_dly_sig_n[43] tdc0.w_dly_sig[43] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3990 VPWR a_7591_3285# a_7507_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3991 a_27438_5853# a_27123_5719# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3992 a_6177_5487# tdc0.w_dly_sig[146] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3993 a_13429_8029# _024_ a_13357_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3995 tdc0.w_dly_sig_n[40] tdc0.w_dly_sig[40] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3996 tdc0.o_result[127] a_8419_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3997 a_21914_17732# a_21707_17673# a_22090_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3998 VGND a_10459_3133# a_10627_3035# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3999 a_12483_2223# a_11619_2229# a_12226_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4000 VGND tdc0.w_dly_sig[169] tdc0.w_dly_sig_n[170] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4001 VPWR a_6027_16091# a_5943_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4002 VGND tdc0.w_dly_sig[122] tdc0.w_dly_sig_n[122] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4003 a_24017_8041# a_23027_7669# a_23891_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4005 tdc0.w_dly_sig_n[64] tdc0.w_dly_sig[63] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4006 VGND tdc0.w_dly_sig_n[119] tdc0.w_dly_sig[120] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4007 a_7239_16367# a_6375_16373# a_6982_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4008 a_19583_11159# a_19867_11145# a_19802_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4009 tdc0.w_dly_sig[113] tdc0.w_dly_sig_n[112] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4010 clknet_4_4_0_clk a_6550_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4011 VGND _086_ a_12526_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X4012 a_19777_12015# tdc0.o_result[6] a_19967_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4013 tdc0.w_dly_sig[58] tdc0.w_dly_sig_n[56] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4014 clknet_4_15_0_clk a_25410_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4015 a_16573_14735# tdc0.w_dly_sig[70] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4016 a_23381_7663# tdc0.w_dly_sig[27] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4017 VGND tdc0.w_dly_sig_n[120] tdc0.w_dly_sig[121] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4018 tdc0.w_dly_sig_n[168] tdc0.w_dly_sig[168] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4019 VPWR tdc0.w_dly_sig_n[114] tdc0.w_dly_sig[116] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4020 _030_ a_17323_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X4021 a_12851_11837# a_11987_11471# a_12594_11583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4022 VPWR a_6246_3967# a_6173_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4023 VGND tdc0.w_dly_sig[189] tdc0.w_dly_sig_n[190] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4024 a_26755_7895# a_26851_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4025 a_20187_10217# a_20058_9961# a_19767_10071# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4026 VGND ui_in[5] a_17634_591# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4027 VGND a_10259_4373# a_10217_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4028 VGND tdc0.w_dly_sig[96] tdc0.w_dly_sig_n[96] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4030 tdc0.w_dly_sig_n[179] tdc0.w_dly_sig[179] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4031 VPWR tdc0.w_dly_sig[11] a_27505_9129# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4032 clknet_4_13_0_clk a_19890_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4033 a_17076_12015# _057_ a_16974_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4034 a_13445_2223# tdc0.w_dly_sig[170] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4035 tdc0.w_dly_sig_n[168] tdc0.w_dly_sig[167] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4036 tdc0.w_dly_sig[101] tdc0.w_dly_sig_n[99] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4037 VPWR _085_ a_12264_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X4038 a_10160_2767# a_9761_2767# a_10034_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4039 VPWR a_4571_17277# a_4739_17179# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4040 VGND clknet_4_1_0_clk a_5823_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4041 a_22461_591# tdc0.w_dly_sig[180] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4042 a_26514_6575# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4043 a_29945_11837# a_29607_11623# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4044 VPWR a_15595_18267# a_15511_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4045 a_21665_10927# a_21327_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4046 VGND tdc0.w_dly_sig[26] tdc0.w_dly_sig_n[26] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4047 VPWR a_24183_15511# _067_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X4048 VGND a_3651_14191# a_3819_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4050 a_30258_6143# a_30090_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4051 a_19591_7093# clknet_4_9_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4052 tdc0.w_dly_sig[161] tdc0.w_dly_sig_n[160] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4053 VPWR tdc0.w_dly_sig_n[121] tdc0.w_dly_sig[123] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4054 a_8454_7637# a_8286_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4055 _066_ a_18703_14985# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4056 tdc0.w_dly_sig_n[104] tdc0.w_dly_sig[104] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4057 a_11739_2045# a_10957_1679# a_11655_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4058 VPWR a_11747_9661# a_11915_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4059 a_5069_9295# a_4903_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4060 tdc0.w_dly_sig_n[61] tdc0.w_dly_sig[60] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4061 a_13082_4719# tdc0.o_result[141] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X4062 a_8753_13647# tdc0.w_dly_sig[125] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4063 VPWR tdc0.w_dly_sig[185] tdc0.w_dly_sig_n[185] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4064 a_29446_5309# a_29173_4943# a_29361_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4065 a_13478_6575# _163_ a_13398_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X4066 VGND a_3007_6575# a_3175_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4067 VPWR _064_ a_24843_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4068 tdc0.w_dly_sig_n[32] tdc0.w_dly_sig[32] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4069 tdc0.o_result[55] a_20011_18517# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4070 a_25598_14735# a_25283_14887# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4071 tdc0.w_dly_sig[130] tdc0.w_dly_sig_n[129] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4072 VPWR tdc0.w_dly_sig_n[34] tdc0.w_dly_sig[36] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4073 tdc0.o_result[55] a_20011_18517# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4074 tdc0.w_dly_sig[53] tdc0.w_dly_sig_n[51] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4075 VPWR a_9926_9813# a_9853_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4076 a_24113_14191# tdc0.o_result[53] a_24029_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4077 a_29607_11623# a_29703_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4078 a_2731_9839# a_1867_9845# a_2474_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4079 a_8335_12015# a_7553_12021# a_8251_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4080 clknet_4_1_0_clk a_6476_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4081 a_24137_3855# _060_ a_24065_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4084 tdc0.w_dly_sig[178] tdc0.w_dly_sig_n[177] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4085 VGND clknet_4_5_0_clk a_4167_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4086 a_20109_3855# _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X4087 VGND tdc0.w_dly_sig[50] tdc0.w_dly_sig_n[51] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4088 a_14821_15823# a_14655_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4089 tdc0.w_dly_sig_n[174] tdc0.w_dly_sig[174] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4090 a_30251_4765# a_30031_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X4091 a_27254_10205# a_26939_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4092 VGND _004_ a_15472_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X4093 a_29611_4631# a_29895_4617# a_29830_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4094 VGND a_10995_11739# a_10953_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4096 a_14729_2229# a_14563_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4097 a_29725_8757# a_29559_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4098 tdc0.o_result[126] a_9431_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4100 tdc0.w_dly_sig_n[75] tdc0.w_dly_sig[75] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4101 VPWR tdc0.w_dly_sig[174] tdc0.w_dly_sig_n[175] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4102 VPWR _030_ a_20039_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X4103 VGND tdc0.w_dly_sig[18] tdc0.w_dly_sig_n[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4106 tdc0.o_result[63] a_22955_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4107 a_14645_10383# tdc0.o_result[90] a_14563_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4108 a_24490_2741# a_24290_3041# a_24639_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4109 _054_ a_17139_8759# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X4110 a_14541_2767# a_13551_2767# a_14415_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4111 a_9393_4405# a_9227_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4112 VPWR tdc0.w_dly_sig[109] tdc0.w_dly_sig_n[110] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4113 a_1849_11471# a_1683_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4115 tdc0.w_dly_sig_n[30] tdc0.w_dly_sig[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4116 VPWR tdc0.w_dly_sig_n[86] tdc0.w_dly_sig[88] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4117 a_5805_3855# a_5639_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4118 tdc0.w_dly_sig[180] tdc0.w_dly_sig_n[178] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4119 VPWR a_19777_12015# uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4120 tdc0.o_result[153] a_4647_4123# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4122 VPWR tdc0.w_dly_sig[40] a_25573_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4123 VPWR a_6430_13077# a_6357_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4124 a_2306_9839# a_1867_9845# a_2221_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4125 VPWR tdc0.w_dly_sig_n[92] tdc0.w_dly_sig[94] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4126 a_19526_7119# a_19211_7271# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4127 a_26702_16911# a_26387_17063# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4128 VGND a_7331_15279# a_7499_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4129 tdc0.w_dly_sig[43] tdc0.w_dly_sig_n[41] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4130 tdc0.w_dly_sig[6] tdc0.w_dly_sig_n[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4131 _116_ a_12539_3424# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X4132 tdc0.w_dly_sig_n[41] tdc0.w_dly_sig[41] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4133 VGND clknet_4_6_0_clk a_14195_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4134 a_6173_4221# a_5639_3855# a_6078_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4136 VGND clknet_4_2_0_clk a_11251_1141# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4137 tdc0.w_dly_sig_n[139] tdc0.w_dly_sig[138] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4139 a_9298_8751# a_9025_8757# a_9213_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4140 a_16547_4373# _042_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X4141 a_21445_5493# a_21279_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4142 a_20574_5193# _033_ a_20325_5089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X4143 a_6883_6183# a_6979_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4145 a_20666_4399# _184_ a_20417_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X4146 tdc0.o_result[135] a_7775_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4147 a_16737_9441# _032_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X4149 tdc0.w_dly_sig[171] tdc0.w_dly_sig_n[169] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4150 VGND tdc0.w_dly_sig_n[154] tdc0.w_dly_sig[156] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4152 a_12594_11583# a_12426_11837# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4153 tdc0.w_dly_sig_n[55] tdc0.w_dly_sig[54] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4154 VPWR _050_ a_23027_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X4155 a_20477_8029# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X4156 tdc0.w_dly_sig[63] tdc0.w_dly_sig_n[62] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4157 VGND tdc0.w_dly_sig[183] a_26125_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4158 VPWR a_26663_4631# tdc0.o_result[188] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4159 VPWR tdc0.w_dly_sig[117] tdc0.w_dly_sig_n[118] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4160 VPWR a_19579_5719# _202_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X4161 tdc0.w_dly_sig_n[52] tdc0.w_dly_sig[52] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4162 a_22102_2589# a_21787_2455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4163 VGND a_15163_3543# _123_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X4164 a_14182_10159# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X4166 VGND tdc0.w_dly_sig[136] tdc0.w_dly_sig_n[137] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4167 a_2674_7663# a_2401_7669# a_2589_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4168 a_5307_8573# a_4443_8207# a_5050_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4169 a_15170_18111# a_15002_18365# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4170 uo_out[3] a_18489_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4171 a_25471_12533# a_25762_12833# a_25713_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X4172 VPWR a_23811_1367# tdc0.o_result[180] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4173 tdc0.w_dly_sig_n[76] tdc0.w_dly_sig[75] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4174 tdc0.w_dly_sig_n[188] tdc0.w_dly_sig[188] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4175 VPWR tdc0.w_dly_sig_n[58] tdc0.w_dly_sig[59] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4176 VPWR a_20359_3855# _051_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4177 VPWR net28 a_28057_5865# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4178 a_9853_9839# a_9319_9845# a_9758_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4179 tdc0.w_dly_sig_n[38] tdc0.w_dly_sig[38] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4180 tdc0.w_dly_sig_n[175] tdc0.w_dly_sig[174] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4181 tdc0.w_dly_sig[64] tdc0.w_dly_sig_n[63] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4182 a_2121_5865# a_1131_5493# a_1995_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4183 clknet_4_14_0_clk a_26882_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4184 a_5161_15823# a_4995_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4185 VGND a_20011_18517# a_19969_18921# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4186 VGND a_12115_3133# a_12283_3035# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4188 a_15236_6575# _077_ a_15134_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4189 tdc0.w_dly_sig_n[59] tdc0.w_dly_sig[59] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4190 tdc0.o_result[60] a_18815_16341# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4191 a_6687_5487# a_5823_5493# a_6430_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4192 VPWR a_10506_7119# clknet_4_3_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4194 tdc0.w_dly_sig_n[151] tdc0.w_dly_sig[150] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4195 VGND tdc0.w_dly_sig_n[148] tdc0.w_dly_sig[150] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4196 a_20258_10116# a_20051_10057# a_20434_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4197 a_24283_15797# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4198 tdc0.w_dly_sig_n[164] tdc0.w_dly_sig[164] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4199 VGND tdc0.w_dly_sig_n[109] tdc0.w_dly_sig[111] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4200 a_30347_10357# ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4201 VGND a_22787_3133# a_22955_3035# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4202 a_7331_15279# a_6467_15285# a_7074_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4203 VPWR a_11839_7663# a_12007_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4204 VPWR _064_ a_19415_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4205 VGND tdc0.w_dly_sig_n[19] tdc0.w_dly_sig[21] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4206 tdc0.w_dly_sig[12] tdc0.w_dly_sig_n[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4207 VGND a_29090_12292# a_29019_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4208 a_25835_9447# a_25931_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4210 VGND tdc0.w_dly_sig_n[108] tdc0.w_dly_sig[109] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4211 tdc0.w_dly_sig[75] tdc0.w_dly_sig_n[74] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4212 a_19119_5719# _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X4213 a_17746_18111# a_17578_18365# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4214 _092_ a_7479_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X4215 tdc0.w_dly_sig[128] tdc0.w_dly_sig_n[126] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4216 tdc0.w_dly_sig_n[72] tdc0.w_dly_sig[72] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4217 VGND tdc0.w_dly_sig_n[111] tdc0.w_dly_sig[112] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4219 VGND tdc0.o_result[132] a_5549_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4220 a_18985_4943# _030_ a_18913_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4221 a_17421_13647# _001_ a_17349_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4222 VGND clknet_4_0_0_clk a_3247_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4223 a_23903_2919# a_23999_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4224 VGND tdc0.w_dly_sig_n[104] tdc0.w_dly_sig[106] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4225 a_20625_9545# _069_ a_20709_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4226 VPWR tdc0.w_dly_sig[16] tdc0.w_dly_sig_n[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4227 a_5721_11721# _171_ a_5639_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4228 a_19777_12015# _190_ a_19505_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4229 VPWR a_23478_6852# a_23407_6953# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4230 tdc0.w_dly_sig[112] tdc0.w_dly_sig_n[110] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4231 a_24837_2767# a_24283_2741# a_24490_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4232 VGND _029_ a_20359_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4233 VGND _050_ a_17201_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4234 a_11417_9661# a_10883_9295# a_11322_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4235 VGND a_17619_2197# a_17577_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4236 a_8399_10633# _027_ a_8481_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4237 tdc0.w_dly_sig_n[53] tdc0.w_dly_sig[52] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4238 tdc0.w_dly_sig[87] tdc0.w_dly_sig_n[86] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4239 a_17194_14165# a_17026_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4240 uo_out[3] a_18489_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4241 a_23110_5487# _031_ a_23110_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X4242 a_15299_12015# _004_ a_15477_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X4243 VGND a_20315_7895# _160_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X4244 a_4314_7637# a_4146_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4245 VGND a_11747_9661# a_11915_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4246 a_24309_15279# _014_ a_24511_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4248 a_7733_7119# a_6743_7119# a_7607_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4249 a_15197_9545# _129_ a_15115_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X4251 _154_ a_22751_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X4252 tdc0.w_dly_sig_n[129] tdc0.w_dly_sig[129] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4253 VPWR a_2899_9813# a_2815_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4254 VPWR tdc0.w_dly_sig_n[52] tdc0.w_dly_sig[53] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4256 _009_ net4 a_17329_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4257 tdc0.w_dly_sig_n[57] tdc0.w_dly_sig[57] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4258 a_19057_591# tdc0.w_dly_sig[175] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4259 tdc0.w_dly_sig_n[3] tdc0.w_dly_sig[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4260 a_9666_4399# a_9227_4405# a_9581_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4261 VGND a_11260_5461# clknet_4_2_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4263 _008_ a_15609_4971# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X4264 VPWR a_12651_2197# a_12567_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4265 a_27179_3855# a_27050_4129# a_26759_3829# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4266 a_21104_6005# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4267 a_14983_7093# _006_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X4268 VPWR tdc0.w_dly_sig_n[22] tdc0.w_dly_sig[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4269 VGND a_21707_11145# a_21714_11049# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4270 VPWR a_19310_703# a_19237_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4271 a_14633_15657# a_13643_15285# a_14507_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4272 tdc0.w_dly_sig[83] tdc0.w_dly_sig_n[81] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4273 a_21166_15101# a_20893_14735# a_21081_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4274 tdc0.w_dly_sig_n[11] tdc0.w_dly_sig[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4275 tdc0.w_dly_sig_n[176] tdc0.w_dly_sig[175] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4276 tdc0.w_dly_sig_n[87] tdc0.w_dly_sig[87] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4277 VGND tdc0.w_dly_sig_n[84] tdc0.w_dly_sig[85] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4278 tdc0.o_result[95] a_10719_17179# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4279 VPWR _056_ a_22615_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X4281 VGND a_2290_12671# a_2248_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4282 a_14760_11305# a_14361_10933# a_14634_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4284 a_24005_8725# _188_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X4285 a_3321_14191# a_2787_14197# a_3226_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4287 a_7883_10927# a_7185_10933# a_7626_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4288 tdc0.o_result[126] a_9431_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4289 a_14158_2879# a_13990_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4290 tdc0.o_result[163] a_10443_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4291 VGND a_26663_4007# tdc0.o_result[189] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4292 VGND a_6476_7637# clknet_4_1_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4293 a_27829_3133# a_27491_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4294 a_30031_4777# a_29895_4617# a_29611_4631# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4296 a_15381_12015# _173_ a_15299_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4297 tdc0.w_dly_sig_n[183] tdc0.w_dly_sig[183] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4298 VPWR _024_ a_14011_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4299 VPWR tdc0.w_dly_sig_n[149] tdc0.w_dly_sig[150] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4300 a_13641_8207# _023_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X4301 a_5859_16189# a_5161_15823# a_5602_15935# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4302 tdc0.w_dly_sig[162] tdc0.w_dly_sig_n[161] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4303 VPWR a_26939_10071# tdc0.o_result[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4305 _201_ a_13722_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X4306 _007_ a_14983_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4307 a_5434_16189# a_4995_15823# a_5349_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4308 a_8661_17455# tdc0.w_dly_sig[97] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4309 tdc0.w_dly_sig[15] tdc0.w_dly_sig_n[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4310 VPWR a_18659_7895# _096_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X4312 a_20434_9839# a_20187_10217# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
R11 uio_oe[4] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4313 VGND tdc0.w_dly_sig_n[166] tdc0.w_dly_sig[167] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4314 VGND a_14887_4631# _162_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X4316 a_22077_13647# _001_ a_22005_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4317 tdc0.w_dly_sig_n[126] tdc0.w_dly_sig[125] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4318 a_24170_11721# tdc0.o_result[48] a_24013_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4319 VPWR a_24611_16341# a_24527_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4320 a_16665_5487# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4321 VPWR tdc0.w_dly_sig[133] tdc0.w_dly_sig_n[134] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4322 VGND tdc0.w_dly_sig[49] tdc0.w_dly_sig_n[49] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4323 VPWR a_14507_17455# a_14675_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4324 a_14103_13647# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4325 VGND a_13019_11739# a_12977_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4326 VGND a_22809_13793# _149_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X4327 a_2217_14013# a_1683_13647# a_2122_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4328 VGND a_14507_17455# a_14675_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4329 a_22813_12559# a_22266_12833# a_22466_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4330 VPWR a_10459_3133# a_10627_3035# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4331 VPWR a_29614_5055# a_29541_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4332 a_25962_15797# a_25755_15797# a_26138_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4333 _205_ a_19058_4719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X4334 a_24837_18921# a_24290_18665# a_24490_18820# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4335 VPWR tdc0.w_dly_sig_n[8] tdc0.w_dly_sig[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4336 VPWR tdc0.w_dly_sig_n[122] tdc0.w_dly_sig[124] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4337 a_23591_11305# a_23455_11145# a_23171_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4338 tdc0.w_dly_sig_n[99] tdc0.w_dly_sig[98] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4339 VPWR a_3819_14165# a_3735_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4340 tdc0.w_dly_sig_n[155] tdc0.w_dly_sig[155] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4341 VPWR tdc0.w_dly_sig[53] tdc0.w_dly_sig_n[53] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4343 tdc0.o_result[12] a_30039_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4344 VPWR tdc0.w_dly_sig_n[99] tdc0.w_dly_sig[100] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4346 VPWR _058_ a_13367_9952# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4347 tdc0.o_result[116] a_4371_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4348 tdc0.w_dly_sig[190] tdc0.w_dly_sig_n[189] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4349 VGND a_25428_7637# clknet_4_10_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4350 a_2290_13759# a_2122_14013# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4351 VGND clknet_4_15_0_clk a_23579_16373# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4352 VPWR tdc0.w_dly_sig[184] tdc0.w_dly_sig_n[185] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4353 VPWR tdc0.o_result[157] a_11711_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4355 tdc0.w_dly_sig[33] tdc0.w_dly_sig_n[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4357 VPWR a_24490_18820# a_24419_18921# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4358 a_10317_17999# tdc0.w_dly_sig[95] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4359 VPWR tdc0.w_dly_sig_n[188] tdc0.w_dly_sig[190] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4360 VGND _050_ a_13392_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X4361 VPWR tdc0.w_dly_sig[191] tdc0.w_dly_sig_n[191] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4362 a_22852_7093# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4363 VGND a_4739_17179# a_4697_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4364 a_13790_16341# a_13622_16367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4365 VPWR _035_ a_14103_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4366 VGND tdc0.w_dly_sig_n[178] tdc0.w_dly_sig[179] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4367 tdc0.w_dly_sig_n[140] tdc0.w_dly_sig[140] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4368 clknet_4_15_0_clk a_25410_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4369 VPWR a_16210_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X4371 a_6262_4399# a_5823_4405# a_6177_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4372 a_11509_6575# a_10975_6581# a_11414_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4373 a_2547_12925# a_1683_12559# a_2290_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4374 tdc0.w_dly_sig[19] tdc0.w_dly_sig_n[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4375 a_10735_12925# a_10037_12559# a_10478_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4377 VPWR tdc0.w_dly_sig_n[81] tdc0.w_dly_sig[83] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4378 VPWR tdc0.w_dly_sig[143] tdc0.w_dly_sig_n[143] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4379 a_22809_13793# _148_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X4380 clknet_4_13_0_clk a_19890_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4381 a_26518_11471# a_26203_11623# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4382 VGND clknet_4_7_0_clk a_10055_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4384 a_16669_11721# _062_ a_16587_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X4385 VPWR a_26663_4007# tdc0.o_result[189] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4386 a_24639_3543# a_24735_3543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4388 a_15793_6281# net6 a_15709_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4389 a_15473_3855# tdc0.o_result[154] a_15391_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4390 VPWR tdc0.w_dly_sig_n[174] tdc0.w_dly_sig[175] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4391 a_3041_4777# a_2051_4405# a_2915_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4392 a_9263_16189# a_8565_15823# a_9006_15935# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4393 tdc0.o_result[145] a_6855_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4394 a_15238_8457# _100_ a_14989_8353# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X4395 a_27035_10071# a_27319_10057# a_27254_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4396 tdc0.o_result[57] a_18171_18267# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4397 VGND tdc0.w_dly_sig_n[34] tdc0.w_dly_sig[35] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4398 VPWR a_14437_8725# _117_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X4400 VPWR a_9815_7485# a_9983_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4401 VPWR tdc0.w_dly_sig[8] a_30541_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4402 a_12353_8207# _085_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X4403 tdc0.w_dly_sig_n[181] tdc0.w_dly_sig[181] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4404 a_29945_10927# a_29607_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4405 VPWR net3 a_15530_6077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X4406 a_16649_12559# _012_ a_16577_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4407 VPWR tdc0.w_dly_sig[1] tdc0.w_dly_sig_n[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4408 VGND clknet_4_7_0_clk a_11987_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4409 a_16784_14735# a_16385_14735# a_16658_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4410 a_9792_4777# a_9393_4405# a_9666_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4411 VGND tdc0.w_dly_sig[177] a_19685_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4412 VGND tdc0.w_dly_sig_n[90] tdc0.w_dly_sig[92] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4414 VPWR net4 a_17323_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X4415 VGND a_10662_14847# a_10620_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4416 a_14507_17455# a_13643_17461# a_14250_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4417 net6 a_18151_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4418 tdc0.w_dly_sig[169] tdc0.w_dly_sig_n[167] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4419 _000_ net6 a_17317_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4420 VPWR a_3394_14165# a_3321_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4421 a_17415_12015# _010_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X4422 tdc0.o_result[35] a_23323_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4423 a_11793_4765# tdc0.o_result[157] a_11711_4512# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4424 VGND tdc0.w_dly_sig[87] tdc0.w_dly_sig_n[88] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4425 clknet_4_3_0_clk a_10506_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4426 a_21366_8207# a_21051_8359# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4427 VPWR a_9466_8725# a_9393_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4428 tdc0.o_result[190] a_30591_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4429 a_11690_3133# a_11417_2767# a_11605_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4430 VPWR a_3559_15279# a_3727_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4431 a_25707_1679# a_25578_1953# a_25287_1653# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4432 VGND tdc0.w_dly_sig[26] a_20421_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4434 VGND a_3559_15279# a_3727_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4435 a_23075_11159# a_23171_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4436 tdc0.o_result[131] a_8879_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4437 a_27250_3829# a_27043_3829# a_27426_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4438 a_5391_6397# a_4609_6031# a_5307_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4439 a_14177_17455# a_13643_17461# a_14082_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4440 VGND a_10202_3967# a_10160_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4441 a_22362_3133# a_22089_2767# a_22277_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4442 a_19591_7093# clknet_4_9_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4443 VPWR tdc0.w_dly_sig_n[92] tdc0.w_dly_sig[93] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4444 tdc0.w_dly_sig[62] tdc0.w_dly_sig_n[60] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4445 a_4287_10927# a_3505_10933# a_4203_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4446 tdc0.w_dly_sig_n[43] tdc0.w_dly_sig[42] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4447 tdc0.w_dly_sig[7] tdc0.w_dly_sig_n[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4448 tdc0.w_dly_sig[98] tdc0.w_dly_sig_n[96] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4449 VGND a_2290_11583# a_2248_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4450 a_8711_7663# a_7847_7669# a_8454_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4452 a_2122_12925# a_1849_12559# a_2037_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4453 tdc0.w_dly_sig_n[191] tdc0.w_dly_sig[191] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4455 a_21380_14165# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4456 VPWR tdc0.w_dly_sig[82] tdc0.w_dly_sig_n[82] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4457 a_29541_5309# a_29007_4943# a_29446_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4458 a_8964_13647# a_8565_13647# a_8838_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4459 VPWR tdc0.w_dly_sig[5] tdc0.w_dly_sig_n[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4460 a_5157_7119# a_4167_7119# a_5031_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4461 VPWR a_2842_7637# a_2769_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4462 VPWR a_5475_8475# a_5391_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4463 a_5434_16189# a_5161_15823# a_5349_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4464 tdc0.w_dly_sig[12] tdc0.w_dly_sig_n[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4465 VPWR a_20051_10057# a_20058_9961# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4466 a_20175_12559# _192_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4467 a_24283_4917# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4469 a_21071_11721# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4470 tdc0.o_result[153] a_4647_4123# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4471 tdc0.w_dly_sig_n[17] tdc0.w_dly_sig[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4472 tdc0.w_dly_sig_n[94] tdc0.w_dly_sig[93] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4473 tdc0.w_dly_sig_n[103] tdc0.w_dly_sig[102] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4474 VPWR _017_ a_17765_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X4475 VGND a_25410_13103# clknet_4_15_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4476 tdc0.w_dly_sig_n[47] tdc0.w_dly_sig[46] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4477 a_11003_15101# a_10221_14735# a_10919_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4478 tdc0.w_dly_sig_n[7] tdc0.w_dly_sig[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4479 tdc0.o_result[128] a_7683_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4480 a_16734_18517# a_16566_18543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4481 a_12723_13647# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4482 a_16692_591# a_16293_591# a_16566_957# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4483 a_20661_5853# _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X4484 _070_ a_19982_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X4485 tdc0.w_dly_sig_n[94] tdc0.w_dly_sig[94] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4486 VPWR a_22374_2500# a_22303_2601# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4487 a_25962_4917# a_25755_4917# a_26138_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4488 tdc0.w_dly_sig[144] tdc0.w_dly_sig_n[143] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4489 VPWR tdc0.w_dly_sig[26] tdc0.w_dly_sig_n[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4490 VPWR tdc0.o_result[122] a_17996_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X4491 tdc0.w_dly_sig_n[141] tdc0.w_dly_sig[141] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4493 tdc0.w_dly_sig[92] tdc0.w_dly_sig_n[91] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4494 a_10735_14013# a_9871_13647# a_10478_13759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4495 VPWR a_6855_5461# a_6771_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4496 a_21905_16911# a_21739_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4497 a_26859_15497# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4498 tdc0.w_dly_sig[159] tdc0.w_dly_sig_n[157] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4499 a_14922_13897# tdc0.o_result[94] a_14839_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4500 a_15232_13647# _058_ a_15112_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X4501 a_13722_6031# _045_ a_13968_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X4502 tdc0.w_dly_sig_n[109] tdc0.w_dly_sig[108] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4503 VGND tdc0.w_dly_sig[165] tdc0.w_dly_sig_n[165] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4506 a_4774_15253# a_4606_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4507 tdc0.w_dly_sig[81] tdc0.w_dly_sig_n[80] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4509 tdc0.w_dly_sig_n[21] tdc0.w_dly_sig[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4510 VPWR clknet_4_5_0_clk a_1683_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4511 VPWR a_19890_13103# clknet_4_13_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4512 tdc0.w_dly_sig[139] tdc0.w_dly_sig_n[137] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4513 VGND tdc0.w_dly_sig_n[114] tdc0.w_dly_sig[115] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4514 a_18843_13335# _054_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X4515 VPWR a_16205_10901# _085_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4516 VPWR tdc0.w_dly_sig[186] a_25757_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4517 tdc0.o_result[11] a_30407_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4518 tdc0.w_dly_sig_n[151] tdc0.w_dly_sig[151] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4519 a_14185_13647# tdc0.o_result[83] a_14103_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4520 clknet_4_14_0_clk a_26882_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4521 a_10773_4943# a_10607_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4522 VPWR tdc0.w_dly_sig[50] a_24837_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4523 VGND tdc0.w_dly_sig[21] tdc0.w_dly_sig_n[22] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4524 a_15002_18365# a_14729_17999# a_14917_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4525 VGND a_29895_4617# a_29902_4521# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4526 VGND a_5307_6397# a_5475_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4527 tdc0.w_dly_sig_n[181] tdc0.w_dly_sig[180] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4528 a_21813_4405# a_21647_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4529 a_16858_16911# a_16543_17063# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4530 VPWR _054_ a_12723_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4531 _011_ a_16495_5487# a_17023_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4532 a_12061_9845# a_11895_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4533 a_6246_3967# a_6078_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4534 a_6388_4777# a_5989_4405# a_6262_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4535 tdc0.w_dly_sig_n[163] tdc0.w_dly_sig[163] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4536 net25 a_29099_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4537 a_17117_11247# tdc0.o_result[42] a_16679_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4538 VGND _067_ a_24131_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4539 VGND tdc0.w_dly_sig[138] tdc0.w_dly_sig_n[138] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4540 tdc0.w_dly_sig_n[56] tdc0.w_dly_sig[56] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4541 a_3559_15279# a_2695_15285# a_3302_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4542 _111_ a_17498_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X4543 a_8753_8207# tdc0.w_dly_sig[131] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4544 tdc0.o_result[177] a_21207_3035# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4545 a_19982_8751# tdc0.o_result[137] a_19899_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4547 VPWR tdc0.w_dly_sig_n[179] tdc0.w_dly_sig[180] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4548 a_19307_7093# a_19591_7093# a_19526_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4549 a_19487_6183# a_19583_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4550 tdc0.w_dly_sig[19] tdc0.w_dly_sig_n[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4551 VPWR a_7378_13103# clknet_4_5_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4553 tdc0.w_dly_sig_n[97] tdc0.w_dly_sig[97] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4554 tdc0.w_dly_sig_n[83] tdc0.w_dly_sig[82] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4555 VPWR tdc0.w_dly_sig_n[30] tdc0.w_dly_sig[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4556 a_11414_7663# a_10975_7669# a_11329_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4557 VPWR clknet_4_7_0_clk a_9963_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4558 a_25665_11471# a_25118_11745# a_25318_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4559 VGND a_5659_15003# a_5617_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4560 VPWR tdc0.w_dly_sig[70] tdc0.w_dly_sig_n[71] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4561 tdc0.w_dly_sig[36] tdc0.w_dly_sig_n[35] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4562 VGND clknet_4_8_0_clk a_18703_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4563 tdc0.w_dly_sig_n[10] tdc0.w_dly_sig[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4565 VPWR clknet_4_7_0_clk a_10055_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4566 VPWR a_12115_3133# a_12283_3035# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4567 a_9393_8751# a_8859_8757# a_9298_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4569 a_19163_9545# _189_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X4570 a_20201_13647# _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X4571 VPWR tdc0.w_dly_sig_n[49] tdc0.w_dly_sig[51] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4572 VPWR a_8895_16367# a_9063_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4573 a_26518_7119# a_26203_7271# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4574 VGND _043_ a_12693_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4575 VPWR tdc0.w_dly_sig[55] tdc0.w_dly_sig_n[56] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4577 VGND a_7423_3311# a_7591_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4578 a_29913_7663# tdc0.w_dly_sig[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4579 a_22891_14423# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X4580 _182_ a_14287_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X4581 VGND a_9891_8725# a_9849_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4582 a_16968_17833# a_16569_17461# a_16842_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4583 VGND a_8895_16367# a_9063_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4584 a_27426_4221# a_27179_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4585 VPWR tdc0.w_dly_sig_n[56] tdc0.w_dly_sig[57] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4586 a_10310_14013# a_10037_13647# a_10225_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4587 VPWR a_22787_3133# a_22955_3035# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4588 a_19651_957# a_18869_591# a_19567_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4589 tdc0.o_result[135] a_7775_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4590 a_11679_8983# _025_ a_11853_9089# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4591 tdc0.w_dly_sig[38] tdc0.w_dly_sig_n[36] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4592 VGND tdc0.w_dly_sig_n[158] tdc0.w_dly_sig[159] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4593 VGND _035_ a_23457_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4594 VPWR a_8251_12015# a_8419_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4595 VPWR a_7867_15003# a_7783_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4596 a_29998_15279# a_29725_15285# a_29913_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4597 a_5989_4405# a_5823_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4598 VGND a_7775_7387# a_7733_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4599 tdc0.o_result[62] a_23139_16091# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4601 tdc0.o_result[160] a_9063_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4602 VPWR tdc0.w_dly_sig[85] tdc0.w_dly_sig_n[86] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4603 tdc0.w_dly_sig_n[122] tdc0.w_dly_sig[122] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4604 a_13081_12381# tdc0.o_result[85] a_12999_12128# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4605 a_16355_7969# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X4606 VGND _033_ a_13722_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X4607 a_18758_2197# a_18590_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4608 tdc0.w_dly_sig_n[142] tdc0.w_dly_sig[142] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4609 tdc0.w_dly_sig_n[84] tdc0.w_dly_sig[84] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4610 tdc0.w_dly_sig[120] tdc0.w_dly_sig_n[119] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4611 tdc0.w_dly_sig[130] tdc0.w_dly_sig_n[128] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4612 a_8895_3311# a_8031_3317# a_8638_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4613 VPWR a_7470_6005# a_7399_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4614 a_28007_2767# a_27871_2741# a_27587_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4615 tdc0.w_dly_sig[157] tdc0.w_dly_sig_n[156] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4616 a_4245_2767# tdc0.w_dly_sig[156] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4617 VPWR clknet_4_13_0_clk a_17139_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4618 a_1922_10901# a_1754_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4619 VGND a_22254_4373# a_22212_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4620 tdc0.w_dly_sig_n[4] tdc0.w_dly_sig[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4621 VPWR a_22852_7093# clknet_4_9_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4622 VPWR clknet_4_2_0_clk a_14563_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4623 clknet_4_13_0_clk a_19890_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4624 a_4606_15279# a_4167_15285# a_4521_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4625 tdc0.w_dly_sig[76] tdc0.w_dly_sig_n[74] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4626 VGND tdc0.w_dly_sig_n[77] tdc0.w_dly_sig[79] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4627 VPWR tdc0.w_dly_sig[156] tdc0.w_dly_sig_n[157] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4628 tdc0.w_dly_sig_n[152] tdc0.w_dly_sig[152] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4630 a_20605_10217# a_20058_9961# a_20258_10116# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4631 a_20138_14165# a_19970_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4632 tdc0.w_dly_sig_n[81] tdc0.w_dly_sig[80] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4633 a_10777_8207# tdc0.w_dly_sig[78] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4634 VGND tdc0.w_dly_sig_n[9] tdc0.w_dly_sig[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4635 tdc0.w_dly_sig_n[190] tdc0.w_dly_sig[190] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4637 tdc0.w_dly_sig_n[12] tdc0.w_dly_sig[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4638 a_3226_3311# a_2953_3317# a_3141_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4639 clknet_4_7_0_clk a_11812_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4640 VGND _137_ a_18059_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X4641 a_30323_9839# a_29541_9845# a_30239_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4642 VGND tdc0.w_dly_sig_n[34] tdc0.w_dly_sig[36] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4643 VGND tdc0.w_dly_sig[1] a_25665_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4644 VGND a_2474_9813# a_2432_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4645 a_1570_7485# a_1297_7119# a_1485_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4646 VGND _091_ a_7479_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4647 a_18317_2229# a_18151_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4648 a_30343_7284# tdc0.w_dly_sig[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4649 a_1481_10933# a_1315_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4650 VPWR tdc0.w_dly_sig[92] tdc0.w_dly_sig_n[93] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4651 VPWR tdc0.w_dly_sig[35] tdc0.w_dly_sig_n[35] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4652 a_25019_3529# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4653 tdc0.w_dly_sig[31] tdc0.w_dly_sig_n[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4654 a_12999_12559# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4655 VPWR tdc0.w_dly_sig_n[159] tdc0.w_dly_sig[161] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4656 VGND net2 a_16495_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4657 VPWR tdc0.w_dly_sig_n[190] tdc0.w_dly_sig[191] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4658 tdc0.o_result[92] a_15595_18267# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4659 tdc0.w_dly_sig[123] tdc0.w_dly_sig_n[121] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4660 a_23040_9129# a_22641_8757# a_22914_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4661 a_23733_17833# a_23186_17577# a_23386_17732# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4662 VPWR a_10995_11739# a_10911_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4664 a_12805_13647# tdc0.o_result[124] a_12723_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4666 VGND tdc0.w_dly_sig_n[48] tdc0.w_dly_sig[50] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4667 a_6913_14191# tdc0.w_dly_sig[124] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4668 VPWR tdc0.w_dly_sig[9] tdc0.w_dly_sig_n[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4669 VGND clknet_0_clk a_12254_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4670 a_20074_6005# a_19867_6005# a_20250_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4671 a_29998_15279# a_29559_15285# a_29913_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4672 VPWR tdc0.w_dly_sig[13] tdc0.w_dly_sig_n[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4673 VGND _153_ a_22751_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4674 VPWR a_23386_17732# a_23315_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4676 VGND tdc0.w_dly_sig_n[94] tdc0.w_dly_sig[96] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4677 a_13149_6549# _164_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X4679 VPWR _058_ a_14878_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
R12 tt_um_hpretl_tt06_tdc_v1_10.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4680 tdc0.w_dly_sig_n[51] tdc0.w_dly_sig[50] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4681 a_17187_13799# tdc0.o_result[64] a_17421_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4682 VPWR tdc0.o_result[160] a_13459_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4683 VPWR clknet_4_1_0_clk a_2235_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4685 a_25203_3829# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4686 a_12460_10217# a_12061_9845# a_12334_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4688 tdc0.w_dly_sig_n[164] tdc0.w_dly_sig[163] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4689 a_20201_5853# _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X4690 clknet_4_10_0_clk a_25428_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4691 a_11540_8041# a_11141_7669# a_11414_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4692 tdc0.w_dly_sig_n[191] tdc0.w_dly_sig[190] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4693 VGND tdc0.w_dly_sig_n[28] tdc0.w_dly_sig[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4694 VPWR tdc0.w_dly_sig[120] tdc0.w_dly_sig_n[121] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4695 a_15128_2601# a_14729_2229# a_15002_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4696 VPWR tdc0.w_dly_sig_n[112] tdc0.w_dly_sig[113] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4697 VPWR tdc0.w_dly_sig_n[84] tdc0.w_dly_sig[86] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4698 tdc0.o_result[118] a_4463_11739# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4699 a_10551_17277# a_9853_16911# a_10294_17023# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4700 VGND a_20138_14165# a_20096_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4701 VPWR a_4279_5461# a_4195_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4702 a_3141_14191# tdc0.w_dly_sig[106] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4703 tdc0.w_dly_sig_n[180] tdc0.w_dly_sig[180] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4704 VPWR tdc0.w_dly_sig[149] tdc0.w_dly_sig_n[149] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4705 tdc0.o_result[156] a_6395_3035# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4706 tdc0.w_dly_sig_n[58] tdc0.w_dly_sig[58] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4708 tdc0.w_dly_sig_n[157] tdc0.w_dly_sig[156] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4709 a_22641_8757# a_22475_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4710 a_16639_16885# a_16930_17185# a_16881_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X4711 a_13349_16373# a_13183_16373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4712 a_17047_3424# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4713 tdc0.w_dly_sig[88] tdc0.w_dly_sig_n[86] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4715 a_27411_13321# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4716 VPWR _040_ a_19931_4737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4717 a_15553_17999# a_14563_17999# a_15427_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4718 VPWR tdc0.w_dly_sig[165] tdc0.w_dly_sig_n[166] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4720 VGND tdc0.w_dly_sig_n[170] tdc0.w_dly_sig[172] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4722 a_20325_5089# _033_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X4723 a_22917_12015# tdc0.o_result[61] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4724 VPWR a_26939_12247# tdc0.o_result[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4725 a_22254_4373# a_22086_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4726 tdc0.o_result[58] a_17435_17429# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4727 a_2217_13103# a_1683_13109# a_2122_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4728 tdc0.w_dly_sig[192] tdc0.w_dly_sig_n[191] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4729 VGND a_21603_4007# _183_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X4730 a_30166_14165# a_29998_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4732 VGND tdc0.w_dly_sig_n[112] tdc0.w_dly_sig[114] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4733 VGND tdc0.w_dly_sig_n[93] tdc0.w_dly_sig[94] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4734 VPWR a_29987_11145# a_29994_11049# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4736 tdc0.w_dly_sig_n[78] tdc0.w_dly_sig[77] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4737 a_2037_13647# tdc0.w_dly_sig[107] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4738 a_29998_14191# a_29725_14197# a_29913_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4740 a_4981_14735# tdc0.w_dly_sig[122] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4741 a_19487_2767# a_19267_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X4742 a_19982_8751# _039_ a_19982_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X4743 VPWR a_22530_2879# a_22457_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4744 VPWR a_1995_7485# a_2163_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4745 VPWR tdc0.w_dly_sig_n[102] tdc0.w_dly_sig[104] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4746 a_9389_8207# a_8399_8207# a_9263_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4747 a_22194_12559# a_21879_12711# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4748 VPWR clknet_4_14_0_clk a_22291_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4749 VGND tdc0.w_dly_sig[186] tdc0.w_dly_sig_n[187] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4750 VPWR tdc0.o_result[25] a_15236_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X4751 tdc0.w_dly_sig[122] tdc0.w_dly_sig_n[120] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4752 VGND net6 a_16560_6935# VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
X4753 a_16691_15823# a_16562_16097# a_16271_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4755 a_13541_3677# tdc0.o_result[160] a_13459_3424# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4756 VGND tdc0.w_dly_sig[77] tdc0.w_dly_sig_n[77] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4757 net1 a_30347_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4758 VPWR net27 a_27689_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4759 a_29814_12925# a_29541_12559# a_29729_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4760 VGND a_24490_15797# a_24419_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4761 tdc0.w_dly_sig_n[14] tdc0.w_dly_sig[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4762 VGND tdc0.w_dly_sig_n[47] tdc0.w_dly_sig[49] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4763 VPWR _076_ a_11803_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4764 a_23903_4007# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X4765 a_16293_18549# a_16127_18549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4767 VPWR tdc0.w_dly_sig[94] tdc0.w_dly_sig_n[95] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4769 VGND _056_ a_14349_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4770 VGND a_26790_7093# a_26719_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4771 VGND a_12651_2197# a_12609_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4772 VPWR tdc0.w_dly_sig[17] tdc0.w_dly_sig_n[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4773 VPWR clknet_4_1_0_clk a_4443_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4774 a_27271_8041# a_27142_7785# a_26851_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4776 VGND _058_ a_22077_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4777 a_10225_12559# tdc0.w_dly_sig[82] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4778 VGND a_18383_8983# _095_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X4779 VGND tdc0.w_dly_sig_n[106] tdc0.w_dly_sig[108] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4780 VGND tdc0.w_dly_sig[14] tdc0.w_dly_sig_n[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4781 a_10528_17999# a_10129_17999# a_10402_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4782 a_20250_6397# a_20003_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4783 VPWR tdc0.w_dly_sig_n[61] tdc0.w_dly_sig[62] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4784 VGND a_28595_7284# net27 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4785 a_8565_13647# a_8399_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4786 tdc0.w_dly_sig_n[127] tdc0.w_dly_sig[126] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4787 VPWR clknet_4_5_0_clk a_4995_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4788 _053_ a_16850_13423# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X4789 _151_ a_17691_14985# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4790 a_29331_7284# tdc0.w_dly_sig[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4791 VPWR _072_ a_5805_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X4792 VPWR tdc0.w_dly_sig[9] a_30541_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4793 VPWR a_10018_2197# a_9945_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4794 VGND clknet_4_10_0_clk a_29007_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4795 a_24659_12015# tdc0.o_result[5] a_24469_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X4796 VPWR tdc0.w_dly_sig[147] tdc0.w_dly_sig_n[147] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4797 VPWR tdc0.w_dly_sig_n[54] tdc0.w_dly_sig[56] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4798 tdc0.w_dly_sig_n[73] tdc0.w_dly_sig[72] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4799 a_11141_6581# a_10975_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4800 a_12526_9295# _088_ a_12772_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X4802 tdc0.w_dly_sig[47] tdc0.w_dly_sig_n[46] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4803 tdc0.w_dly_sig[111] tdc0.w_dly_sig_n[109] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4804 a_19825_10927# a_19487_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4805 VPWR a_30347_10357# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4806 VPWR a_24490_4917# a_24419_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4807 VGND tdc0.w_dly_sig[153] tdc0.w_dly_sig_n[153] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4808 a_13081_12559# tdc0.o_result[87] a_12999_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4810 a_17351_17455# a_16569_17461# a_17267_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4811 tdc0.w_dly_sig[179] tdc0.w_dly_sig_n[177] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4812 tdc0.o_result[107] a_2715_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4813 a_13997_7637# _013_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X4814 VGND a_5050_8319# a_5008_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4816 a_17695_6575# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X4818 VGND tdc0.w_dly_sig[95] tdc0.w_dly_sig_n[96] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4819 VPWR tdc0.o_result[80] a_16679_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4820 a_16623_3133# a_15925_2767# a_16366_2879# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4821 VGND a_12191_18517# a_12149_18921# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4822 VGND tdc0.w_dly_sig[44] tdc0.w_dly_sig_n[44] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4823 tdc0.w_dly_sig_n[170] tdc0.w_dly_sig[169] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4825 VGND _026_ a_12877_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4826 tdc0.w_dly_sig[100] tdc0.w_dly_sig_n[99] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4827 a_24218_2767# a_23903_2919# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4828 tdc0.w_dly_sig[39] tdc0.w_dly_sig_n[37] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4829 a_1937_6031# a_947_6031# a_1811_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4831 VGND tdc0.w_dly_sig[25] tdc0.w_dly_sig_n[25] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4832 VGND net3 a_15293_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4833 VPWR tdc0.w_dly_sig[124] tdc0.w_dly_sig_n[124] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4834 a_17937_10927# tdc0.o_result[2] a_18127_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4836 a_22261_17833# a_21707_17673# a_21914_17732# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4837 a_25203_3829# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4838 tdc0.w_dly_sig[40] tdc0.w_dly_sig_n[38] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4839 a_3946_10901# a_3778_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4840 a_15105_10383# tdc0.o_result[105] a_15023_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4841 a_21147_8181# a_21431_8181# a_21366_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4842 a_22603_17277# a_21739_16911# a_22346_17023# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4843 VGND a_22346_17023# a_22304_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4844 tdc0.w_dly_sig_n[183] tdc0.w_dly_sig[182] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4845 a_24266_11471# _010_ a_24176_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X4846 tdc0.w_dly_sig[163] tdc0.w_dly_sig_n[161] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4847 a_14082_15279# a_13643_15285# a_13997_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4848 a_24241_16189# a_23903_15975# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4850 tdc0.o_result[122] a_6855_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4851 VPWR a_21914_11204# a_21843_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4852 a_2490_4399# a_2217_4405# a_2405_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4854 VGND a_14215_16341# a_14173_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4855 VGND tdc0.w_dly_sig[55] tdc0.w_dly_sig_n[55] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4856 a_6550_12559# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4857 a_27597_3855# a_27050_4129# a_27250_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4859 a_22273_17277# a_21739_16911# a_22178_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4860 VGND tdc0.w_dly_sig[114] tdc0.w_dly_sig_n[115] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4861 tdc0.w_dly_sig[53] tdc0.w_dly_sig_n[52] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4862 a_22929_12335# tdc0.o_result[37] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4863 a_23466_7663# a_23193_7669# a_23381_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4864 a_30541_11471# a_29987_11445# a_30194_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4865 VPWR tdc0.w_dly_sig[57] tdc0.w_dly_sig_n[58] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4866 tdc0.w_dly_sig[189] tdc0.w_dly_sig_n[188] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4867 VGND tdc0.w_dly_sig_n[68] tdc0.w_dly_sig[69] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4868 VPWR tdc0.w_dly_sig_n[69] tdc0.w_dly_sig[71] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4869 tdc0.w_dly_sig_n[36] tdc0.w_dly_sig[36] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4870 VGND clknet_4_4_0_clk a_1867_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4871 VGND _076_ a_14533_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4872 VGND a_5199_7387# a_5157_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4873 a_14729_10927# a_14195_10933# a_14634_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4874 tdc0.w_dly_sig[91] tdc0.w_dly_sig_n[89] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4876 VGND _054_ a_21031_13675# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4877 tdc0.o_result[169] a_14123_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4878 VGND tdc0.w_dly_sig_n[51] tdc0.w_dly_sig[52] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4879 VPWR tdc0.w_dly_sig_n[76] tdc0.w_dly_sig[78] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4880 tdc0.w_dly_sig_n[174] tdc0.w_dly_sig[173] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4881 a_23903_15975# a_23999_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4882 VGND tdc0.w_dly_sig[189] tdc0.w_dly_sig_n[189] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4883 a_19338_2741# a_19138_3041# a_19487_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4884 a_7373_10927# tdc0.w_dly_sig[80] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4885 VPWR tdc0.o_result[167] a_12999_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4886 tdc0.o_result[177] a_21207_3035# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4887 a_16307_8029# net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X4889 _145_ a_18046_4719# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X4890 VGND _069_ a_20072_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X4891 a_13955_2223# a_13091_2229# a_13698_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4892 VPWR tdc0.w_dly_sig_n[55] tdc0.w_dly_sig[56] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4893 VGND a_15427_18365# a_15595_18267# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4895 a_24569_16745# a_23579_16373# a_24443_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4896 tdc0.w_dly_sig_n[139] tdc0.w_dly_sig[139] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4897 VGND tdc0.w_dly_sig_n[88] tdc0.w_dly_sig[90] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4898 VPWR tdc0.w_dly_sig_n[174] tdc0.w_dly_sig[176] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4900 VGND tdc0.w_dly_sig[144] tdc0.w_dly_sig_n[145] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4902 VPWR tdc0.w_dly_sig[80] tdc0.w_dly_sig_n[80] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4904 a_8711_7663# a_8013_7669# a_8454_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4905 VPWR tdc0.o_result[120] a_15483_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4906 a_19629_3677# _038_ a_19557_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4907 _064_ net5 a_17703_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4908 tdc0.w_dly_sig_n[156] tdc0.w_dly_sig[156] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4909 tdc0.w_dly_sig_n[77] tdc0.w_dly_sig[76] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4910 VPWR a_3394_3285# a_3321_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4911 VGND tdc0.w_dly_sig[152] tdc0.w_dly_sig_n[153] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4912 VPWR tdc0.w_dly_sig_n[10] tdc0.w_dly_sig[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4913 VGND clknet_4_5_0_clk a_1683_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4916 tdc0.w_dly_sig_n[18] tdc0.w_dly_sig[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4917 a_14813_9545# _080_ a_14741_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4918 VPWR tdc0.w_dly_sig_n[57] tdc0.w_dly_sig[58] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4919 VPWR tdc0.w_dly_sig[122] tdc0.w_dly_sig_n[123] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4920 VPWR a_22511_4399# a_22679_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4923 tdc0.w_dly_sig[102] tdc0.w_dly_sig_n[101] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4924 VPWR a_30166_3285# a_30093_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4925 VGND tdc0.w_dly_sig_n[62] tdc0.w_dly_sig[64] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4926 VGND a_23903_15975# tdc0.o_result[49] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4927 a_14721_11445# _004_ a_14878_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X4928 tdc0.o_result[116] a_4371_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4929 VGND a_23903_2919# tdc0.o_result[183] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4930 VGND clknet_0_clk a_26514_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4931 a_19049_14735# tdc0.o_result[57] a_18703_14985# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4932 VPWR a_16301_6575# a_16401_6691# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X4934 VGND tdc0.w_dly_sig_n[24] tdc0.w_dly_sig[25] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4935 a_15465_12015# tdc0.o_result[142] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4936 a_12552_11471# a_12153_11471# a_12426_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4937 VGND a_30515_6397# a_30683_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4938 VPWR tdc0.w_dly_sig[39] tdc0.w_dly_sig_n[39] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4939 tdc0.o_result[83] a_11087_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4940 _005_ a_15203_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4941 a_10478_13759# a_10310_14013# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4942 tdc0.w_dly_sig[183] tdc0.w_dly_sig_n[182] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4943 VPWR a_14250_18517# a_14177_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4944 a_27618_13380# a_27418_13225# a_27767_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4945 VPWR a_17937_10927# uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4946 a_23171_11159# a_23462_11049# a_23413_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X4947 a_12525_5487# tdc0.w_dly_sig[145] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4948 a_14897_9813# _081_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X4949 VGND _122_ a_12618_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X4950 VGND a_10735_14013# a_10903_13915# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4951 tdc0.w_dly_sig_n[137] tdc0.w_dly_sig[136] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4952 a_27491_2919# a_27587_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4953 a_14257_13647# _058_ a_14185_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4954 a_25410_13103# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4955 a_12539_10383# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4956 a_13081_3677# tdc0.o_result[167] a_12999_3424# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4957 VPWR a_23139_859# a_23055_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4959 a_6629_12335# tdc0.o_result[103] a_6191_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4960 VPWR _043_ a_12999_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4962 tdc0.o_result[178] a_21391_1947# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4963 a_26299_7093# a_26583_7093# a_26518_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4964 tdc0.w_dly_sig[17] tdc0.w_dly_sig_n[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4965 a_12618_7983# _124_ a_12864_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X4966 VPWR tdc0.w_dly_sig_n[66] tdc0.w_dly_sig[68] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4967 a_22254_4373# a_22086_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4968 a_23913_8353# _108_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X4969 clknet_4_13_0_clk a_19890_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4970 VPWR _064_ a_20887_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4971 tdc0.o_result[108] a_2715_11739# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4972 VPWR _038_ a_16635_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X4973 _181_ a_13722_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X4975 a_2305_11305# a_1315_10933# a_2179_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4976 a_9815_7485# a_9117_7119# a_9558_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4978 a_22971_16189# a_22273_15823# a_22714_15935# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4979 VPWR tdc0.w_dly_sig[21] tdc0.w_dly_sig_n[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4980 VPWR tdc0.o_result[9] a_19899_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X4981 a_19912_15657# a_19513_15285# a_19786_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4983 VPWR a_25191_1831# tdc0.o_result[182] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4984 tdc0.w_dly_sig[91] tdc0.w_dly_sig_n[90] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4985 a_8838_9661# a_8399_9295# a_8753_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4986 tdc0.w_dly_sig[174] tdc0.w_dly_sig_n[172] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4988 VGND tdc0.w_dly_sig_n[134] tdc0.w_dly_sig[136] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4989 a_29814_9839# a_29541_9845# a_29729_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4990 a_29738_5853# a_29423_5719# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4991 a_23097_15823# a_22107_15823# a_22971_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4992 a_27319_10057# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4993 VPWR a_22346_17023# a_22273_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4994 VGND a_11812_13621# clknet_4_7_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4995 a_13809_15285# a_13643_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4996 a_20273_13647# _011_ a_20201_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4997 VPWR a_5123_12015# a_5291_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4999 VGND tdc0.w_dly_sig_n[144] tdc0.w_dly_sig[145] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5000 a_18659_7895# tdc0.o_result[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5001 VGND tdc0.w_dly_sig_n[79] tdc0.w_dly_sig[81] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5002 VPWR clknet_4_4_0_clk a_3431_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5004 a_9117_7119# a_8951_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5006 VPWR tdc0.w_dly_sig[67] tdc0.w_dly_sig_n[67] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5007 VPWR tdc0.w_dly_sig_n[43] tdc0.w_dly_sig[44] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5008 a_29982_12671# a_29814_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5009 VGND a_5123_12015# a_5291_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5010 tdc0.w_dly_sig_n[157] tdc0.w_dly_sig[157] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5011 tdc0.w_dly_sig_n[1] tdc0.w_dly_sig[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5012 a_12539_3424# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5013 VGND tdc0.w_dly_sig[104] tdc0.w_dly_sig_n[104] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5014 tdc0.o_result[67] a_15687_16091# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5015 a_22511_4399# a_21813_4405# a_22254_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5016 tdc0.w_dly_sig[92] tdc0.w_dly_sig_n[90] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5017 tdc0.w_dly_sig_n[134] tdc0.w_dly_sig[134] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5018 VGND _014_ a_20348_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X5019 VGND tdc0.w_dly_sig_n[78] tdc0.w_dly_sig[80] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5020 a_5802_3133# a_5363_2767# a_5717_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5021 a_17121_14191# a_16587_14197# a_17026_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5022 VPWR a_23903_2919# tdc0.o_result[183] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5023 a_17220_12335# tdc0.o_result[56] a_16645_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X5024 a_19947_4007# tdc0.o_result[190] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5025 tdc0.w_dly_sig_n[127] tdc0.w_dly_sig[127] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5027 a_3321_3311# a_2787_3317# a_3226_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5028 a_26767_16885# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5029 a_19685_2767# a_19131_2741# a_19338_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X5030 a_16916_4373# _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X5031 VPWR a_28687_16599# tdc0.o_result[46] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5032 a_13153_12381# _034_ a_13081_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5033 VGND _026_ a_14533_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5034 a_4479_4221# a_3781_3855# a_4222_3967# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5035 VGND a_24490_2741# a_24419_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X5036 tdc0.w_dly_sig_n[79] tdc0.w_dly_sig[79] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5038 a_24735_13621# a_25019_13621# a_24954_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5039 VPWR a_23075_11159# tdc0.o_result[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5040 VGND tdc0.w_dly_sig_n[163] tdc0.w_dly_sig[165] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5041 a_15203_5309# a_15023_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5043 a_30093_3311# a_29559_3317# a_29998_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5044 VPWR tdc0.w_dly_sig[155] tdc0.w_dly_sig_n[155] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5045 VGND tdc0.w_dly_sig[172] tdc0.w_dly_sig_n[172] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5046 a_27491_2919# a_27587_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5048 a_20499_13799# tdc0.o_result[55] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5049 VGND a_11823_1947# a_11781_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5050 a_7189_14735# tdc0.w_dly_sig[126] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5051 a_19885_14191# tdc0.w_dly_sig[69] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5052 a_6262_13103# a_5823_13109# a_6177_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5054 a_21334_14847# a_21166_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5055 VGND clknet_0_clk a_25410_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5056 a_16734_703# a_16566_957# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5057 a_19899_8751# _039_ a_19982_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X5058 tdc0.w_dly_sig_n[5] tdc0.w_dly_sig[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5059 VPWR a_25318_11445# a_25247_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5060 _026_ a_15351_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5061 VGND _192_ a_20175_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5062 tdc0.w_dly_sig[25] tdc0.w_dly_sig_n[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5063 a_9558_7231# a_9390_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5064 VGND a_19890_13103# clknet_4_13_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5065 tdc0.w_dly_sig[3] tdc0.w_dly_sig_n[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5066 a_6246_3967# a_6078_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5067 VPWR a_17619_14165# a_17535_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5068 VGND tdc0.w_dly_sig_n[127] tdc0.w_dly_sig[128] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5069 a_24490_2741# a_24283_2741# a_24666_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5070 a_11214_5055# a_11046_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5071 VPWR tdc0.w_dly_sig_n[27] tdc0.w_dly_sig[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5072 a_19586_18517# a_19418_18543# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5073 a_10919_15101# a_10055_14735# a_10662_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5074 _119_ a_13735_14304# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5076 VGND tdc0.w_dly_sig_n[6] tdc0.w_dly_sig[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5077 VPWR tdc0.w_dly_sig[19] tdc0.w_dly_sig_n[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5078 VGND tdc0.w_dly_sig[47] tdc0.w_dly_sig_n[48] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5079 VPWR tdc0.w_dly_sig[153] tdc0.w_dly_sig_n[154] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5080 a_29997_4943# a_29007_4943# a_29871_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5081 a_3183_7663# a_2401_7669# a_3099_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5082 VPWR a_21759_15003# a_21675_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5083 tdc0.w_dly_sig_n[66] tdc0.w_dly_sig[65] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5084 clknet_4_14_0_clk a_26882_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5085 a_24525_3855# _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X5086 a_22277_15279# tdc0.w_dly_sig[64] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5089 a_24653_9545# _090_ a_24381_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5090 VPWR a_19671_10071# tdc0.o_result[33] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5091 a_25287_1653# a_25578_1953# a_25529_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5092 a_20022_9545# _033_ a_19773_9441# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5093 VPWR a_10570_18111# a_10497_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5094 a_10589_15101# a_10055_14735# a_10494_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5095 VGND _010_ a_18479_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5096 tdc0.w_dly_sig_n[114] tdc0.w_dly_sig[114] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5097 VGND tdc0.w_dly_sig_n[53] tdc0.w_dly_sig[54] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5098 VGND tdc0.w_dly_sig[130] tdc0.w_dly_sig_n[131] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5099 uo_out[4] a_19225_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5100 a_26571_8983# a_26667_8983# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5101 VPWR a_6476_7637# clknet_4_1_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5102 tdc0.w_dly_sig_n[117] tdc0.w_dly_sig[116] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5103 a_20625_9545# _070_ a_20543_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5104 a_12877_13647# _022_ a_12805_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5105 VGND tdc0.w_dly_sig_n[143] tdc0.w_dly_sig[145] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5106 VGND tdc0.w_dly_sig_n[141] tdc0.w_dly_sig[143] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5107 VGND a_4774_15253# a_4732_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5108 a_19893_10383# tdc0.o_result[144] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X5109 tdc0.w_dly_sig_n[33] tdc0.w_dly_sig[33] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5110 VGND tdc0.w_dly_sig[54] a_24837_18921# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5111 a_23745_16373# a_23579_16373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5112 a_20881_11721# _063_ a_20609_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5113 a_20175_12559# _194_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5114 a_10662_14847# a_10494_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5115 tdc0.w_dly_sig_n[134] tdc0.w_dly_sig[133] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5116 tdc0.w_dly_sig_n[65] tdc0.w_dly_sig[65] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5117 VGND tdc0.w_dly_sig_n[69] tdc0.w_dly_sig[70] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5118 a_2037_13103# tdc0.w_dly_sig[112] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5119 VPWR a_19867_11145# a_19874_11049# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5120 uo_out[3] a_18489_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5121 tdc0.o_result[103] a_6027_16091# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5122 VPWR a_30423_15279# a_30591_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5123 a_27135_7881# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5125 VPWR a_17691_6281# _033_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5126 VGND clknet_4_15_0_clk a_29559_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5127 a_26299_11445# a_26590_11745# a_26541_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5128 VPWR tdc0.w_dly_sig[135] tdc0.w_dly_sig_n[136] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5129 a_12935_15101# a_12153_14735# a_12851_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5130 a_8964_9295# a_8565_9295# a_8838_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5132 a_22511_4399# a_21647_4405# a_22254_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5135 VGND a_30423_15279# a_30591_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5136 VPWR _011_ a_19807_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X5137 a_10543_3133# a_9761_2767# a_10459_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5139 tdc0.o_result[109] a_1979_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5140 VPWR tdc0.w_dly_sig[178] tdc0.w_dly_sig_n[179] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5141 a_2953_3317# a_2787_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5142 VGND tdc0.w_dly_sig_n[25] tdc0.w_dly_sig[27] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5143 a_2248_13647# a_1849_13647# a_2122_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5144 VGND tdc0.w_dly_sig_n[165] tdc0.w_dly_sig[166] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5145 a_13735_14304# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5146 a_16385_14735# a_16219_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5148 VPWR tdc0.w_dly_sig[123] tdc0.w_dly_sig_n[123] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5149 a_22005_13647# tdc0.o_result[66] a_21923_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5150 a_21389_8573# a_21051_8359# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5151 VGND a_9431_8475# a_9389_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5152 VPWR a_17194_14165# a_17121_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5153 VPWR a_24639_13799# tdc0.o_result[39] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5154 VPWR a_30258_6143# a_30185_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5155 a_9006_15935# a_8838_16189# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5156 _135_ a_12999_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5157 VPWR a_23634_7637# a_23561_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5158 VGND tdc0.w_dly_sig_n[151] tdc0.w_dly_sig[153] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5159 VPWR tdc0.w_dly_sig[188] tdc0.w_dly_sig_n[189] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5160 VPWR tdc0.w_dly_sig[59] tdc0.w_dly_sig_n[59] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5162 a_5928_2767# a_5529_2767# a_5802_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5163 VPWR a_21787_2455# tdc0.o_result[181] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5164 tdc0.o_result[178] a_21391_1947# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5165 VGND tdc0.w_dly_sig_n[72] tdc0.w_dly_sig[73] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5166 VPWR tdc0.w_dly_sig_n[33] tdc0.w_dly_sig[35] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5168 VPWR tdc0.w_dly_sig_n[95] tdc0.w_dly_sig[97] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5169 clknet_4_2_0_clk a_11260_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5170 VGND clknet_4_1_0_clk a_4443_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5171 a_9171_17455# a_8473_17461# a_8914_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5172 _174_ a_15299_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X5173 a_13866_6281# _041_ a_13552_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X5174 VPWR tdc0.w_dly_sig[5] tdc0.w_dly_sig_n[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5175 a_19418_18543# a_18979_18549# a_19333_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5176 tdc0.w_dly_sig[88] tdc0.w_dly_sig_n[87] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5177 tdc0.w_dly_sig_n[86] tdc0.w_dly_sig[85] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5178 a_19221_13793# _206_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X5179 a_17741_9323# _019_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X5180 VGND a_20051_10057# a_20058_9961# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5181 a_3969_3855# tdc0.w_dly_sig[154] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5182 tdc0.w_dly_sig[147] tdc0.w_dly_sig_n[146] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5183 a_12445_9295# _085_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X5184 VPWR tdc0.w_dly_sig_n[44] tdc0.w_dly_sig[45] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5185 tdc0.w_dly_sig_n[19] tdc0.w_dly_sig[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5186 a_18137_16367# tdc0.w_dly_sig[61] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5187 tdc0.w_dly_sig_n[161] tdc0.w_dly_sig[160] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5188 a_28503_12247# a_28599_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5189 a_24666_3133# a_24419_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5190 a_8565_13647# a_8399_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5191 VPWR tdc0.w_dly_sig_n[153] tdc0.w_dly_sig[155] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5193 VGND a_14415_3133# a_14583_3035# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5194 a_27321_16911# a_26774_17185# a_26974_16885# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5195 VPWR tdc0.w_dly_sig_n[184] tdc0.w_dly_sig[185] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5196 VGND a_11839_7663# a_12007_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5197 tdc0.o_result[35] a_23323_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5198 VGND a_25375_8983# _106_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X5199 a_17218_3855# tdc0.o_result[138] a_17137_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X5200 VPWR clknet_0_clk a_11260_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5201 tdc0.w_dly_sig_n[116] tdc0.w_dly_sig[115] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5202 VGND tdc0.w_dly_sig_n[7] tdc0.w_dly_sig[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5203 a_15645_15823# a_14655_15823# a_15519_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5204 VPWR tdc0.o_result[162] a_14103_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5205 a_11141_7669# a_10975_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5206 tdc0.w_dly_sig_n[90] tdc0.w_dly_sig[90] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5208 VGND tdc0.w_dly_sig_n[39] tdc0.w_dly_sig[41] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5211 a_30365_10217# a_29375_9845# a_30239_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5213 tdc0.w_dly_sig[104] tdc0.w_dly_sig_n[102] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5214 a_22546_957# a_22273_591# a_22461_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5215 a_20614_3133# a_20175_2767# a_20529_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5216 VPWR _007_ a_12907_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5218 a_23478_6852# a_23271_6793# a_23654_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5219 VPWR tdc0.w_dly_sig_n[149] tdc0.w_dly_sig[151] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5220 clknet_4_5_0_clk a_7378_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5221 a_11839_6397# a_11141_6031# a_11582_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5222 tdc0.w_dly_sig[36] tdc0.w_dly_sig_n[34] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5225 VPWR clknet_4_4_0_clk a_1315_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5226 tdc0.w_dly_sig_n[35] tdc0.w_dly_sig[35] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5227 VPWR _040_ a_13735_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5228 VGND a_11582_6549# a_11540_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5229 a_13722_6031# tdc0.o_result[136] a_13641_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X5230 VGND a_3394_3285# a_3352_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5231 a_13149_6549# _162_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
R13 VPWR tt_um_hpretl_tt06_tdc_v1_9.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5232 a_19470_13897# _208_ a_19221_13793# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5233 VGND _118_ a_14274_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X5234 VPWR a_5031_7485# a_5199_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5235 VGND tdc0.w_dly_sig[88] tdc0.w_dly_sig_n[88] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5236 VPWR tdc0.w_dly_sig[110] tdc0.w_dly_sig_n[111] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5237 VGND a_11455_8475# a_11413_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5239 VGND a_25502_8181# a_25431_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X5241 a_23999_2741# a_24283_2741# a_24218_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5242 a_8013_7669# a_7847_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5243 a_22259_12533# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5244 VGND tdc0.w_dly_sig[3] tdc0.w_dly_sig_n[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5245 VGND tdc0.w_dly_sig[6] tdc0.w_dly_sig_n[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5247 VPWR tdc0.w_dly_sig_n[39] tdc0.w_dly_sig[40] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5248 VPWR tdc0.w_dly_sig_n[169] tdc0.w_dly_sig[171] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5250 a_25891_15823# a_25762_16097# a_25471_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5251 VPWR a_24013_11445# _015_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X5252 tdc0.w_dly_sig_n[192] tdc0.w_dly_sig[192] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5253 a_17923_5719# a_18196_5719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5254 tdc0.o_result[128] a_7683_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5255 tdc0.w_dly_sig[101] tdc0.w_dly_sig_n[100] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5256 tdc0.w_dly_sig[62] tdc0.w_dly_sig_n[61] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5257 a_22461_591# tdc0.w_dly_sig[180] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5258 a_22291_14304# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5259 a_13153_12559# _034_ a_13081_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5261 VGND tdc0.w_dly_sig[63] tdc0.w_dly_sig_n[63] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5262 a_16301_6575# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5263 a_11679_8983# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X5264 a_12517_15657# a_11527_15285# a_12391_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5265 clknet_4_10_0_clk a_25428_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5266 VGND a_23339_8751# a_23507_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5267 a_25573_13647# a_25026_13921# a_25226_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5268 VGND tdc0.w_dly_sig[8] tdc0.w_dly_sig_n[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5269 VPWR tdc0.w_dly_sig_n[82] tdc0.w_dly_sig[83] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5270 VGND tdc0.w_dly_sig_n[59] tdc0.w_dly_sig[61] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5271 VGND a_24611_16341# a_24569_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5272 a_26755_7895# a_26851_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5273 clknet_0_clk a_16210_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5274 a_12334_9839# a_12061_9845# a_12249_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5275 tdc0.w_dly_sig[96] tdc0.w_dly_sig_n[94] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5276 VPWR a_13790_16341# a_13717_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5277 a_4701_15279# a_4167_15285# a_4606_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5278 a_15419_4737# _038_ a_15333_4737# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X5279 tdc0.o_result[78] a_10351_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5280 a_14549_10927# tdc0.w_dly_sig[77] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5281 a_20153_10383# tdc0.o_result[32] a_19715_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5282 clknet_4_9_0_clk a_22852_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5283 a_30185_6397# a_29651_6031# a_30090_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5284 a_7479_11471# _023_ a_7657_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
R14 VGND uio_out[5] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5285 tdc0.w_dly_sig_n[72] tdc0.w_dly_sig[71] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5286 VGND a_21380_14165# clknet_4_12_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5287 VPWR a_29982_9813# a_29909_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5288 tdc0.o_result[99] a_9431_16091# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5289 _175_ a_18151_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5290 a_23561_7663# a_23027_7669# a_23466_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5291 a_26817_15279# a_26479_15511# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5292 tdc0.w_dly_sig_n[46] tdc0.w_dly_sig[45] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5293 a_21843_17833# a_21707_17673# a_21423_17687# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5294 VGND tdc0.w_dly_sig_n[136] tdc0.w_dly_sig[137] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5295 a_15220_15823# a_14821_15823# a_15094_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5296 VPWR a_30423_14191# a_30591_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5297 VPWR a_22167_2441# a_22174_2345# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5298 a_11490_9407# a_11322_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5299 tdc0.w_dly_sig[86] tdc0.w_dly_sig_n[84] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5301 a_15177_10383# _022_ a_15105_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5302 a_17967_10159# _064_ a_18489_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5303 a_29423_16733# a_29203_16745# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X5304 VGND a_15575_591# net2 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5305 VPWR tdc0.w_dly_sig[137] tdc0.w_dly_sig_n[138] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5306 a_22825_10749# a_22291_10383# a_22730_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5307 a_29913_8751# tdc0.w_dly_sig[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5308 VGND a_16737_9441# _037_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X5310 a_13968_12809# _199_ a_13866_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X5311 tdc0.w_dly_sig[185] tdc0.w_dly_sig_n[184] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5312 tdc0.o_result[163] a_10443_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5313 VGND tdc0.w_dly_sig[98] tdc0.w_dly_sig_n[98] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5314 VPWR _058_ a_22291_14304# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5315 VGND _056_ a_20053_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5316 VPWR tdc0.w_dly_sig_n[153] tdc0.w_dly_sig[154] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5317 tdc0.o_result[13] a_30591_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5318 a_11141_14197# a_10975_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5319 tdc0.o_result[28] a_22311_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5320 VGND tdc0.w_dly_sig_n[116] tdc0.w_dly_sig[117] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5321 a_16385_14735# a_16219_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5322 tdc0.w_dly_sig_n[37] tdc0.w_dly_sig[37] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5323 a_10091_4399# a_9393_4405# a_9834_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5324 VPWR clknet_4_6_0_clk a_11895_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5325 a_17415_11247# _092_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5326 VGND tdc0.w_dly_sig[149] tdc0.w_dly_sig_n[150] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5327 VPWR a_17267_17455# a_17435_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5328 VGND tdc0.w_dly_sig_n[144] tdc0.w_dly_sig[146] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5329 VPWR tdc0.o_result[91] a_14868_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X5331 VGND a_5970_2879# a_5928_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5332 VPWR tdc0.w_dly_sig_n[45] tdc0.w_dly_sig[46] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5333 a_19746_5193# _033_ a_19497_5089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5335 tdc0.o_result[84] a_12007_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5336 VGND a_17267_17455# a_17435_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5337 VGND a_7699_3133# a_7867_3035# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5338 a_21787_3543# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X5339 a_8573_10927# tdc0.o_result[135] a_8491_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5340 VGND tdc0.w_dly_sig_n[16] tdc0.w_dly_sig[18] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5341 _178_ a_12907_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5342 VGND tdc0.w_dly_sig[128] tdc0.w_dly_sig_n[129] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5343 VGND a_23269_9813# _129_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X5344 a_7400_14735# a_7001_14735# a_7274_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5346 VPWR a_10506_7119# clknet_4_3_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5347 net5 a_17507_1143# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5348 VPWR tdc0.w_dly_sig_n[130] tdc0.w_dly_sig[131] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5349 tdc0.w_dly_sig_n[165] tdc0.w_dly_sig[165] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5350 a_23654_6575# a_23407_6953# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5351 a_20697_12809# tdc0.o_result[7] a_20887_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X5352 tdc0.w_dly_sig_n[82] tdc0.w_dly_sig[82] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5353 _057_ a_16311_3424# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5354 _079_ a_14195_3424# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5355 tdc0.w_dly_sig_n[98] tdc0.w_dly_sig[97] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5357 VPWR a_16219_1143# net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5358 VGND tdc0.w_dly_sig_n[68] tdc0.w_dly_sig[70] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5359 VGND a_14250_15253# a_14208_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5360 VPWR tdc0.w_dly_sig_n[70] tdc0.w_dly_sig[71] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5361 VGND tdc0.w_dly_sig[177] tdc0.w_dly_sig_n[178] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5362 VPWR _177_ a_19413_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5363 a_6814_16367# a_6541_16373# a_6729_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5365 VGND a_8546_2197# a_8504_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5366 a_6227_3133# a_5529_2767# a_5970_2879# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5367 VGND clknet_4_13_0_clk a_16127_18549# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5368 VPWR a_9431_16091# a_9347_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5370 VGND a_7607_7485# a_7775_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5371 tdc0.w_dly_sig_n[167] tdc0.w_dly_sig[166] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5372 tdc0.w_dly_sig[159] tdc0.w_dly_sig_n[158] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5373 a_20740_2767# a_20341_2767# a_20614_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5374 VPWR tdc0.w_dly_sig_n[106] tdc0.w_dly_sig[107] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5375 a_15226_9839# _082_ a_15146_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X5376 a_18413_591# a_18236_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X5377 VGND tdc0.w_dly_sig_n[29] tdc0.w_dly_sig[30] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5378 tdc0.w_dly_sig[86] tdc0.w_dly_sig_n[85] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5379 uo_out[7] a_20697_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5380 a_26541_7485# a_26203_7271# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5381 tdc0.w_dly_sig[108] tdc0.w_dly_sig_n[106] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5382 a_25755_4917# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5383 clknet_4_0_0_clk a_6476_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5384 VPWR tdc0.w_dly_sig[139] tdc0.w_dly_sig_n[139] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5385 tdc0.w_dly_sig_n[108] tdc0.w_dly_sig[107] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5387 a_13249_8867# _161_ a_13177_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5388 tdc0.w_dly_sig_n[26] tdc0.w_dly_sig[26] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5389 VPWR clknet_4_9_0_clk a_23027_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5390 a_24283_18761# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5391 a_21327_17687# a_21423_17687# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5392 VPWR tdc0.w_dly_sig[31] tdc0.w_dly_sig_n[32] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5393 a_16665_5487# net6 a_17023_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5395 tdc0.w_dly_sig_n[169] tdc0.w_dly_sig[169] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5396 _041_ a_13735_4512# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5397 a_17168_9545# _031_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X5398 VGND tdc0.w_dly_sig_n[0] tdc0.w_dly_sig[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5399 a_18390_16341# a_18222_16367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5400 a_20017_8207# _054_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X5401 a_8838_8573# a_8565_8207# a_8753_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5402 a_22546_13103# a_22107_13109# a_22461_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5404 VPWR tdc0.w_dly_sig_n[138] tdc0.w_dly_sig[140] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5405 VGND tdc0.w_dly_sig[62] tdc0.w_dly_sig_n[63] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5406 a_15695_4971# _005_ a_15609_4971# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X5407 VPWR a_4774_15253# a_4701_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5410 tdc0.w_dly_sig_n[101] tdc0.w_dly_sig[101] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5411 a_2290_12671# a_2122_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5412 VPWR tdc0.w_dly_sig_n[47] tdc0.w_dly_sig[48] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5413 VGND tdc0.w_dly_sig_n[75] tdc0.w_dly_sig[76] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5414 VGND tdc0.w_dly_sig_n[64] tdc0.w_dly_sig[65] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5415 _153_ a_13082_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X5416 a_17267_17455# a_16403_17461# a_17010_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5417 a_18233_10383# tdc0.o_result[70] a_18151_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5418 VGND a_11260_5461# clknet_4_2_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5419 VPWR tdc0.w_dly_sig_n[175] tdc0.w_dly_sig[177] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5420 a_22466_12533# a_22266_12833# a_22615_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5421 tdc0.o_result[154] a_3819_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5423 VGND tdc0.w_dly_sig[148] tdc0.w_dly_sig_n[148] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5424 VGND tdc0.w_dly_sig[15] tdc0.w_dly_sig_n[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5425 a_9117_7119# a_8951_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5426 tdc0.w_dly_sig_n[116] tdc0.w_dly_sig[116] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5427 a_24827_11445# a_25111_11445# a_25046_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5428 tdc0.w_dly_sig_n[44] tdc0.w_dly_sig[44] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5429 VPWR a_22898_10495# a_22825_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5431 VPWR a_24283_15797# a_24290_16097# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5432 a_11681_3855# _026_ a_11609_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5433 VPWR a_29067_16585# a_29074_16489# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5434 a_28883_13321# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5435 tdc0.o_result[190] a_30591_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5436 VPWR a_10903_12827# a_10819_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5437 a_13552_12809# tdc0.o_result[127] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X5438 a_14887_4631# tdc0.o_result[181] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5439 VGND tdc0.w_dly_sig[32] tdc0.w_dly_sig_n[32] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5440 a_21081_14735# tdc0.w_dly_sig[67] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5441 a_7549_3689# a_6559_3317# a_7423_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5442 tdc0.w_dly_sig[149] tdc0.w_dly_sig_n[148] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5443 tdc0.w_dly_sig_n[124] tdc0.w_dly_sig[124] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5444 VPWR a_20563_14165# a_20479_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5445 a_24191_1353# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5446 VGND a_23811_1367# tdc0.o_result[180] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5447 net3 a_16219_1143# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5448 VGND a_9466_8725# a_9424_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5449 VPWR a_6687_13103# a_6855_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5450 VGND tdc0.w_dly_sig[102] tdc0.w_dly_sig_n[103] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5451 a_13990_3133# a_13717_2767# a_13905_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5452 a_27702_12015# a_27455_12393# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5453 a_21567_8207# a_21431_8181# a_21147_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5454 a_10294_17023# a_10126_17277# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5455 a_12851_16189# a_11987_15823# a_12594_15935# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5456 VGND a_12594_15935# a_12552_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5459 VGND tdc0.w_dly_sig_n[119] tdc0.w_dly_sig[121] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5460 a_20039_13799# tdc0.o_result[43] a_20273_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5461 VGND a_6687_13103# a_6855_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5462 a_18590_2223# a_18151_2229# a_18505_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5464 a_20250_10927# a_20003_11305# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5465 a_14913_16911# a_14747_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5466 a_21039_3133# a_20341_2767# a_20782_2879# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5467 a_16941_2223# tdc0.w_dly_sig[173] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5468 VGND a_25191_1831# tdc0.o_result[182] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5469 VGND a_12007_14165# a_11965_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5470 VGND tdc0.w_dly_sig[131] tdc0.w_dly_sig_n[132] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5473 tdc0.w_dly_sig[181] tdc0.w_dly_sig_n[180] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5474 tdc0.w_dly_sig_n[159] tdc0.w_dly_sig[159] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5475 tdc0.o_result[118] a_4463_11739# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5476 VPWR clknet_4_4_0_clk a_3339_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5477 tdc0.w_dly_sig[136] tdc0.w_dly_sig_n[135] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5478 tdc0.w_dly_sig_n[107] tdc0.w_dly_sig[107] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5479 VGND tdc0.w_dly_sig_n[93] tdc0.w_dly_sig[95] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5480 VGND a_16733_4917# _038_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0878 ps=0.92 w=0.65 l=0.15
X5481 a_5342_9661# a_5069_9295# a_5257_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5482 a_11693_15285# a_11527_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5483 VPWR tdc0.w_dly_sig_n[124] tdc0.w_dly_sig[125] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5484 a_17665_10927# _110_ a_17937_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5485 VPWR tdc0.w_dly_sig[2] tdc0.w_dly_sig_n[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5487 tdc0.w_dly_sig_n[108] tdc0.w_dly_sig[108] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5488 tdc0.w_dly_sig[13] tdc0.w_dly_sig_n[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5489 VPWR tdc0.w_dly_sig_n[67] tdc0.w_dly_sig[68] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5490 a_24837_2767# a_24290_3041# a_24490_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5491 a_25428_7637# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5492 a_4425_8757# a_4259_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5493 tdc0.w_dly_sig[172] tdc0.w_dly_sig_n[170] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5495 VGND tdc0.w_dly_sig[28] a_20145_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5496 VGND a_25428_7637# clknet_4_10_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5497 a_13997_18543# tdc0.w_dly_sig[92] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5498 VGND a_15538_12671# a_15496_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5499 tdc0.w_dly_sig[90] tdc0.w_dly_sig_n[88] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5500 a_17194_2197# a_17026_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5501 a_14887_4631# tdc0.o_result[181] a_15121_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5502 VPWR tdc0.w_dly_sig[134] tdc0.w_dly_sig_n[134] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5503 tdc0.w_dly_sig[60] tdc0.w_dly_sig_n[58] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5504 VPWR tdc0.w_dly_sig_n[23] tdc0.w_dly_sig[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5505 VPWR tdc0.w_dly_sig[89] tdc0.w_dly_sig_n[89] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5506 VPWR tdc0.w_dly_sig_n[80] tdc0.w_dly_sig[82] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5507 VGND tdc0.w_dly_sig[71] tdc0.w_dly_sig_n[71] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5508 a_19579_5719# tdc0.o_result[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5509 VGND a_15101_7637# _047_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X5510 VPWR tdc0.w_dly_sig[12] tdc0.w_dly_sig_n[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5511 tdc0.w_dly_sig[165] tdc0.w_dly_sig_n[164] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5512 a_14369_3855# tdc0.o_result[158] a_14287_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5513 a_10129_17999# a_9963_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5514 VPWR tdc0.w_dly_sig[16] tdc0.w_dly_sig_n[17] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5515 VPWR tdc0.w_dly_sig_n[73] tdc0.w_dly_sig[74] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5516 VGND tdc0.w_dly_sig_n[36] tdc0.w_dly_sig[37] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5517 a_14208_18921# a_13809_18549# a_14082_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5518 VGND a_30166_14165# a_30124_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5520 VPWR tdc0.w_dly_sig[191] tdc0.w_dly_sig_n[192] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5521 tdc0.w_dly_sig[117] tdc0.w_dly_sig_n[116] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5522 a_17306_17277# a_17059_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5523 VPWR a_17565_8725# _097_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X5524 a_29607_11623# a_29703_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5525 a_4571_7663# a_3873_7669# a_4314_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5526 VPWR tdc0.w_dly_sig_n[50] tdc0.w_dly_sig[51] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5527 VPWR tdc0.w_dly_sig[150] tdc0.w_dly_sig_n[150] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5528 VPWR tdc0.w_dly_sig_n[165] tdc0.w_dly_sig[167] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5531 VGND a_10919_15101# a_11087_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5532 tdc0.o_result[161] a_8971_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5533 a_12434_8207# tdc0.o_result[77] a_12353_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X5535 VPWR a_15351_7093# _026_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5537 a_11471_5309# a_10607_4943# a_11214_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5538 VGND a_9006_13759# a_8964_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5539 a_3141_3311# tdc0.w_dly_sig[155] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5540 a_17493_17999# tdc0.w_dly_sig[58] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5541 a_23855_14735# _055_ a_24033_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5544 VGND _054_ a_12877_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5545 VGND tdc0.w_dly_sig[76] tdc0.w_dly_sig_n[76] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5546 tdc0.w_dly_sig[37] tdc0.w_dly_sig_n[35] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5547 tdc0.o_result[152] a_3083_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5548 tdc0.w_dly_sig[10] tdc0.w_dly_sig_n[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5549 tdc0.w_dly_sig[16] tdc0.w_dly_sig_n[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5550 VPWR a_12502_9813# a_12429_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5551 VPWR a_14415_3133# a_14583_3035# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5552 VGND clknet_4_0_0_clk a_7295_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5554 a_2290_11583# a_2122_11837# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5555 a_19715_10383# _008_ a_19893_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5556 VGND tdc0.w_dly_sig_n[130] tdc0.w_dly_sig[132] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5557 a_29940_10217# a_29541_9845# a_29814_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5559 a_7274_3133# a_7001_2767# a_7189_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5560 tdc0.w_dly_sig[68] tdc0.w_dly_sig_n[66] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5561 a_10506_7119# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5562 VPWR _050_ a_12999_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X5564 tdc0.w_dly_sig[1] tdc0.w_dly_sig_n[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5565 a_11417_2767# a_11251_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5566 a_19579_5719# tdc0.o_result[15] a_19813_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5568 VGND tdc0.w_dly_sig_n[41] tdc0.w_dly_sig[42] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5569 tdc0.w_dly_sig_n[135] tdc0.w_dly_sig[135] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5570 VPWR tdc0.w_dly_sig[68] tdc0.w_dly_sig_n[68] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5571 VPWR tdc0.w_dly_sig_n[40] tdc0.w_dly_sig[41] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5572 a_16635_4007# tdc0.o_result[173] a_16869_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5573 a_24977_3311# a_24639_3543# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5574 a_27526_12292# a_27319_12233# a_27702_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5575 VPWR tdc0.w_dly_sig_n[185] tdc0.w_dly_sig[187] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5576 a_18217_9839# _130_ a_18489_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5577 VGND tdc0.w_dly_sig_n[107] tdc0.w_dly_sig[108] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5578 VGND a_11812_13621# clknet_4_7_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5579 _093_ a_13551_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5580 a_15795_12925# a_14931_12559# a_15538_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5581 a_14081_2601# a_13091_2229# a_13955_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5582 VGND _140_ a_13354_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X5583 a_20074_11204# a_19867_11145# a_20250_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5584 VGND a_26974_16885# a_26903_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X5585 a_27070_8029# a_26755_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5586 tdc0.w_dly_sig_n[71] tdc0.w_dly_sig[70] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5587 VGND _132_ a_18703_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5588 a_22089_2767# a_21923_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5590 VGND a_30407_9813# a_30365_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5591 a_12429_9839# a_11895_9845# a_12334_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5593 a_28883_12233# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5594 VPWR clknet_4_1_0_clk a_3707_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5595 VPWR tdc0.w_dly_sig_n[95] tdc0.w_dly_sig[96] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5596 VGND tdc0.w_dly_sig_n[104] tdc0.w_dly_sig[105] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5597 VGND tdc0.w_dly_sig_n[67] tdc0.w_dly_sig[69] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5598 clknet_4_5_0_clk a_7378_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5599 a_8009_11305# a_7019_10933# a_7883_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5601 a_16765_11721# _053_ a_16669_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X5602 tdc0.w_dly_sig[168] tdc0.w_dly_sig_n[166] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5603 VPWR a_5767_9661# a_5935_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5604 tdc0.w_dly_sig[66] tdc0.w_dly_sig_n[64] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5605 tdc0.o_result[71] a_13019_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5606 a_27455_12393# a_27319_12233# a_27035_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5607 a_18716_2601# a_18317_2229# a_18590_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5608 VPWR tdc0.w_dly_sig[95] tdc0.w_dly_sig_n[95] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5609 VGND a_19119_5719# _078_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X5610 a_8753_9295# tdc0.w_dly_sig[127] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5611 a_19967_12015# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5612 a_25778_1653# a_25571_1653# a_25954_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5613 a_15465_12925# a_14931_12559# a_15370_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5614 tdc0.w_dly_sig[81] tdc0.w_dly_sig_n[79] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5615 a_26759_4631# a_27043_4617# a_26978_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5616 VPWR tdc0.w_dly_sig_n[54] tdc0.w_dly_sig[55] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5617 VGND clknet_4_11_0_clk a_29559_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5618 VPWR tdc0.w_dly_sig_n[7] tdc0.w_dly_sig[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5619 VPWR a_21591_15101# a_21759_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5620 tdc0.w_dly_sig[186] tdc0.w_dly_sig_n[184] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5622 VGND tdc0.w_dly_sig_n[1] tdc0.w_dly_sig[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5623 tdc0.w_dly_sig[111] tdc0.w_dly_sig_n[110] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5624 VPWR _051_ a_11527_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5625 tdc0.w_dly_sig_n[23] tdc0.w_dly_sig[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5626 VPWR a_15519_16189# a_15687_16091# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5627 VPWR a_22633_4917# _133_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X5628 a_17923_5719# a_18196_5719# a_18154_5847# VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5629 VGND clknet_0_clk a_22852_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5630 a_21642_11293# a_21327_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5631 a_21431_8181# clknet_4_9_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5632 VPWR _012_ a_17415_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X5633 a_23825_6953# a_23278_6697# a_23478_6852# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5634 VGND a_6855_5461# a_6813_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5635 VPWR _038_ a_15163_3543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5636 a_11214_5055# a_11046_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5637 VGND a_12559_15253# a_12517_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5638 VGND a_11582_7637# a_11540_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5639 a_11049_9295# a_10883_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5640 a_5717_2767# tdc0.w_dly_sig[157] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5641 a_11747_9661# a_10883_9295# a_11490_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5642 VGND tdc0.w_dly_sig[8] a_30541_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5645 a_26667_8983# a_26951_8969# a_26886_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5646 tdc0.o_result[129] a_9891_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5647 VPWR tdc0.w_dly_sig_n[182] tdc0.w_dly_sig[183] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5648 tdc0.o_result[112] a_2899_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5649 a_19396_8457# _159_ a_19294_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X5650 a_17130_16885# a_16923_16885# a_17306_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5651 VPWR _056_ a_16311_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5652 VPWR _056_ a_14195_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5653 a_22259_12533# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5654 VPWR tdc0.w_dly_sig_n[30] tdc0.w_dly_sig[32] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5655 a_24837_15823# a_24290_16097# a_24490_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5656 VPWR a_24731_11623# tdc0.o_result[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5657 VPWR tdc0.w_dly_sig[132] tdc0.w_dly_sig_n[133] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5658 a_26309_12559# a_25755_12533# a_25962_12533# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X5659 a_30449_4777# a_29895_4617# a_30102_4676# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X5660 tdc0.w_dly_sig[179] tdc0.w_dly_sig_n[178] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5661 VGND a_5031_7485# a_5199_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5662 VPWR _007_ a_15333_4737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5663 VGND tdc0.w_dly_sig_n[176] tdc0.w_dly_sig[178] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5664 tdc0.o_result[134] a_9983_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5665 a_15420_8457# _098_ a_15318_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X5666 a_11812_13621# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5667 VPWR _002_ a_18383_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5668 VGND a_12502_9813# a_12460_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5669 VPWR tdc0.w_dly_sig[42] tdc0.w_dly_sig_n[42] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5671 a_13082_4399# _039_ a_13082_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X5672 a_3133_6953# a_2143_6581# a_3007_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5673 a_11241_9117# tdc0.o_result[129] a_11159_8864# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5674 a_17059_16911# a_16923_16885# a_16639_16885# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5675 a_12153_11471# a_11987_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5676 a_8293_2223# tdc0.w_dly_sig[162] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5677 a_6913_3311# tdc0.w_dly_sig[159] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5678 a_22913_15657# a_21923_15285# a_22787_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5679 VGND a_10183_9839# a_10351_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5680 VGND tdc0.w_dly_sig[67] tdc0.w_dly_sig_n[68] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5681 a_28687_16599# a_28783_16599# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5682 VPWR clknet_4_0_0_clk a_1131_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5683 VPWR tdc0.w_dly_sig[185] tdc0.w_dly_sig_n[186] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5684 tdc0.w_dly_sig_n[146] tdc0.w_dly_sig[146] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5685 tdc0.w_dly_sig[63] tdc0.w_dly_sig_n[61] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5686 VPWR a_7699_3133# a_7867_3035# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5688 a_17695_6575# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5689 a_22645_10383# tdc0.w_dly_sig[36] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5691 _124_ a_11435_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5692 VGND a_7378_13103# clknet_4_5_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5693 a_26939_12247# a_27035_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5694 a_9389_15823# a_8399_15823# a_9263_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5695 VGND _054_ a_18857_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5696 tdc0.w_dly_sig[132] tdc0.w_dly_sig_n[131] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5697 a_28599_12247# a_28890_12137# a_28841_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5698 tdc0.w_dly_sig[54] tdc0.w_dly_sig_n[53] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5699 a_19267_2767# a_19138_3041# a_18847_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5701 VGND tdc0.w_dly_sig[6] a_27873_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5702 tdc0.w_dly_sig_n[144] tdc0.w_dly_sig[143] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5705 tdc0.w_dly_sig[142] tdc0.w_dly_sig_n[141] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5709 a_19119_5719# tdc0.o_result[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5710 a_3873_16911# a_3707_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5711 a_26909_8751# a_26571_8983# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5712 VGND a_18751_2919# tdc0.o_result[176] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5713 a_30278_4399# a_30031_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5714 VPWR _010_ a_20315_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5715 VGND clknet_4_0_0_clk a_7939_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5716 tdc0.w_dly_sig_n[163] tdc0.w_dly_sig[162] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5717 a_29913_15279# tdc0.w_dly_sig[46] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5718 VPWR tdc0.w_dly_sig[156] tdc0.w_dly_sig_n[156] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5719 VPWR tdc0.w_dly_sig[190] a_27597_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5720 tdc0.w_dly_sig_n[37] tdc0.w_dly_sig[36] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5721 VPWR a_22714_703# a_22641_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5722 VPWR a_5859_16189# a_6027_16091# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5723 VGND tdc0.w_dly_sig[22] tdc0.w_dly_sig_n[22] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5724 a_18617_9117# _002_ a_18545_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5725 VPWR tdc0.w_dly_sig[39] a_26309_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5726 a_11417_2767# a_11251_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5727 a_19967_12015# tdc0.o_result[6] a_19777_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X5728 VGND _017_ a_17117_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X5729 VPWR a_25111_7093# a_25118_7393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5730 tdc0.w_dly_sig[6] tdc0.w_dly_sig_n[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5731 a_10585_2767# a_9595_2767# a_10459_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5732 VPWR a_15538_12671# a_15465_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5733 a_8159_4399# a_7295_4405# a_7902_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5734 VGND tdc0.w_dly_sig_n[63] tdc0.w_dly_sig[65] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5735 a_22714_15935# a_22546_16189# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5736 VGND tdc0.w_dly_sig[73] tdc0.w_dly_sig_n[73] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5737 a_17498_12335# tdc0.o_result[107] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X5738 a_20529_2767# tdc0.w_dly_sig[178] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5739 VGND _017_ a_24293_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X5740 VPWR tdc0.o_result[39] a_19652_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X5741 a_23937_14985# _193_ a_23855_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5742 a_7005_10383# tdc0.w_dly_sig[129] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5743 a_27806_2767# a_27491_2919# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5744 VGND a_23903_4007# _128_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X5745 VGND _011_ a_15177_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5746 VGND a_12283_1109# a_12241_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5747 _000_ net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5748 VGND a_23891_7663# a_24059_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5749 VGND tdc0.w_dly_sig[20] tdc0.w_dly_sig_n[20] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5751 a_22089_2767# a_21923_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5753 a_9850_2223# a_9577_2229# a_9765_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5754 VPWR tdc0.w_dly_sig_n[158] tdc0.w_dly_sig[160] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5755 VGND a_16210_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5756 a_29203_16745# a_29074_16489# a_28783_16599# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5757 _208_ a_18703_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5758 VPWR tdc0.o_result[123] a_13735_14304# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5759 VPWR a_24653_9545# uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5761 a_11141_6031# a_10975_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5762 a_11260_5461# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5763 a_29450_16367# a_29203_16745# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5764 VPWR tdc0.w_dly_sig_n[29] tdc0.w_dly_sig[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5765 _169_ a_12434_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X5766 VPWR tdc0.w_dly_sig[132] tdc0.w_dly_sig_n[132] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5768 a_9213_8751# tdc0.w_dly_sig[130] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5769 VGND a_14721_11445# _091_ VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X5770 a_14703_3543# tdc0.o_result[169] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5771 a_9263_9661# a_8399_9295# a_9006_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5772 a_3962_4399# a_3689_4405# a_3877_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5773 VPWR a_19777_12015# uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5774 a_29922_11471# a_29607_11623# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5775 a_11839_6575# a_10975_6581# a_11582_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5776 tdc0.w_dly_sig[30] tdc0.w_dly_sig_n[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5777 VPWR tdc0.w_dly_sig[151] tdc0.w_dly_sig_n[151] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5778 VPWR a_12254_13103# clknet_4_6_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5779 VPWR a_5510_9407# a_5437_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5780 a_18773_16745# a_17783_16373# a_18647_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5781 tdc0.w_dly_sig[73] tdc0.w_dly_sig_n[72] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5782 a_13633_11471# tdc0.o_result[74] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5783 VPWR a_16739_7895# _021_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X5784 a_22167_2441# clknet_4_8_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5785 _126_ a_23303_3424# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5786 a_20549_8029# _010_ a_20477_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5787 _194_ a_23855_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5788 a_19119_5719# tdc0.o_result[17] a_19353_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5789 VPWR a_19395_3543# _204_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X5790 clknet_4_1_0_clk a_6476_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5791 a_9949_3855# tdc0.w_dly_sig[139] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5792 a_19015_2223# a_18317_2229# a_18758_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5793 a_14917_17999# tdc0.w_dly_sig[93] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5794 tdc0.w_dly_sig[149] tdc0.w_dly_sig_n[147] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5795 tdc0.w_dly_sig_n[146] tdc0.w_dly_sig[145] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5796 tdc0.w_dly_sig[55] tdc0.w_dly_sig_n[53] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5797 a_11858_2879# a_11690_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5798 a_22269_5865# a_21279_5493# a_22143_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5800 VPWR a_28503_12247# tdc0.o_result[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5801 VGND a_22971_13103# a_23139_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5802 a_30507_8751# a_29725_8757# a_30423_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5803 a_7001_2767# a_6835_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5804 VPWR a_30166_7637# a_30093_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5806 a_15731_7271# net6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X5807 tdc0.w_dly_sig_n[190] tdc0.w_dly_sig[189] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5809 a_15611_17277# a_14747_16911# a_15354_17023# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5810 VGND a_15354_17023# a_15312_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5811 a_27413_15657# a_26866_15401# a_27066_15556# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5812 _143_ a_12171_4512# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5813 a_25375_5095# a_25471_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5814 VGND a_5767_9661# a_5935_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5815 clknet_4_5_0_clk a_7378_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5816 a_5077_10633# tdc0.o_result[110] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5817 tdc0.w_dly_sig_n[140] tdc0.w_dly_sig[139] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5818 tdc0.w_dly_sig[144] tdc0.w_dly_sig_n[142] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5819 VGND tdc0.w_dly_sig_n[79] tdc0.w_dly_sig[80] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5820 tdc0.w_dly_sig[24] tdc0.w_dly_sig_n[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5821 a_8933_8573# a_8399_8207# a_8838_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5822 a_22530_2879# a_22362_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5823 tdc0.w_dly_sig_n[9] tdc0.w_dly_sig[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5824 a_23937_13647# tdc0.o_result[62] a_23855_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5825 tdc0.w_dly_sig[41] tdc0.w_dly_sig_n[39] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5826 a_22829_8751# tdc0.w_dly_sig[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5827 a_12426_15101# a_12153_14735# a_12341_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5829 a_26217_14735# a_25663_14709# a_25870_14709# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X5830 VPWR a_18751_2919# tdc0.o_result[176] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5831 _203_ a_11527_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5832 VPWR tdc0.w_dly_sig_n[3] tdc0.w_dly_sig[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5833 a_18190_4399# _142_ a_17876_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X5834 a_13817_14557# tdc0.o_result[123] a_13735_14304# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5835 VGND a_2715_13915# a_2673_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5836 tdc0.w_dly_sig[182] tdc0.w_dly_sig_n[180] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5837 VGND a_6687_4399# a_6855_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5838 a_15281_17277# a_14747_16911# a_15186_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5839 tdc0.w_dly_sig_n[152] tdc0.w_dly_sig[151] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5840 a_19225_11721# _150_ a_18953_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5842 VGND tdc0.w_dly_sig[171] tdc0.w_dly_sig_n[171] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5843 tdc0.w_dly_sig_n[192] tdc0.w_dly_sig[191] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5844 VPWR tdc0.w_dly_sig_n[88] tdc0.w_dly_sig[89] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5845 a_16623_3133# a_15759_2767# a_16366_2879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5846 a_14703_3543# tdc0.o_result[169] a_14937_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5847 a_1386_6397# a_947_6031# a_1301_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5848 tdc0.w_dly_sig[106] tdc0.w_dly_sig_n[104] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5849 tdc0.w_dly_sig_n[175] tdc0.w_dly_sig[175] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5850 a_11858_1109# a_11690_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5851 VGND a_22615_4007# _163_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X5852 a_10225_13647# tdc0.w_dly_sig[83] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5853 VPWR tdc0.w_dly_sig[177] tdc0.w_dly_sig_n[177] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5854 a_21292_14735# a_20893_14735# a_21166_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5855 a_29913_3311# tdc0.w_dly_sig[191] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5856 a_19513_18543# a_18979_18549# a_19418_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5857 VPWR tdc0.w_dly_sig_n[159] tdc0.w_dly_sig[160] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5858 _043_ a_17231_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X5859 clknet_0_clk a_16210_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5860 clknet_4_9_0_clk a_22852_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5861 a_19505_12015# _174_ a_19255_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5862 VPWR tdc0.w_dly_sig[190] tdc0.w_dly_sig_n[191] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5863 VGND a_24469_12015# uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5864 VPWR a_7442_2879# a_7369_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5865 a_19567_957# a_18703_591# a_19310_703# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5866 a_9723_8751# a_9025_8757# a_9466_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5867 a_20798_2045# a_20359_1679# a_20713_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5868 tdc0.w_dly_sig[137] tdc0.w_dly_sig_n[135] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5869 clknet_4_4_0_clk a_6550_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5870 a_19338_2741# a_19131_2741# a_19514_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5871 _044_ a_13459_3424# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5872 a_19225_11721# tdc0.o_result[4] a_19415_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X5873 a_1922_10901# a_1754_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5875 tdc0.w_dly_sig_n[29] tdc0.w_dly_sig[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5876 tdc0.w_dly_sig[61] tdc0.w_dly_sig_n[59] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5877 a_1895_6397# a_1113_6031# a_1811_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5878 a_22721_2601# a_22174_2345# a_22374_2500# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5879 VPWR tdc0.w_dly_sig_n[9] tdc0.w_dly_sig[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5880 a_27321_16911# a_26767_16885# a_26974_16885# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X5881 tdc0.w_dly_sig[48] tdc0.w_dly_sig_n[47] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5882 tdc0.w_dly_sig_n[2] tdc0.w_dly_sig[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5883 VPWR tdc0.w_dly_sig_n[167] tdc0.w_dly_sig[168] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5884 VPWR tdc0.w_dly_sig[48] tdc0.w_dly_sig_n[48] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5885 a_29913_14191# tdc0.w_dly_sig[45] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5886 a_11766_18517# a_11598_18543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5887 a_21423_17687# a_21714_17577# a_21665_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5888 a_29274_16644# a_29067_16585# a_29450_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5889 _031_ a_18737_6059# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X5890 a_4793_14735# a_4627_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5891 VPWR a_2715_11739# a_2631_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5892 a_4609_6031# a_4443_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5893 a_10957_8573# a_10423_8207# a_10862_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5895 a_7641_10383# a_6651_10383# a_7515_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5896 VPWR _019_ a_18737_6059# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5897 a_24436_8751# _186_ a_24334_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X5898 tdc0.w_dly_sig_n[66] tdc0.w_dly_sig[66] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5899 a_19497_5089# _033_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X5900 VPWR a_23269_9813# _129_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X5901 tdc0.w_dly_sig_n[98] tdc0.w_dly_sig[98] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5903 VGND tdc0.w_dly_sig_n[60] tdc0.w_dly_sig[61] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5904 VPWR tdc0.w_dly_sig[41] a_27965_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5905 a_21051_8359# a_21147_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5906 VPWR tdc0.w_dly_sig[96] tdc0.w_dly_sig_n[97] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5907 VPWR tdc0.w_dly_sig_n[98] tdc0.w_dly_sig[99] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5908 VPWR tdc0.w_dly_sig[140] tdc0.w_dly_sig_n[141] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5909 VGND tdc0.w_dly_sig_n[52] tdc0.w_dly_sig[54] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5910 a_19954_15253# a_19786_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5911 VPWR clknet_4_6_0_clk a_10975_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5912 tdc0.w_dly_sig[192] tdc0.w_dly_sig_n[190] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5913 VPWR tdc0.w_dly_sig[112] tdc0.w_dly_sig_n[112] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5914 tdc0.w_dly_sig_n[142] tdc0.w_dly_sig[141] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5915 a_24183_15511# _066_ a_24511_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5916 a_14274_13423# _119_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X5917 VPWR tdc0.w_dly_sig_n[148] tdc0.w_dly_sig[149] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5918 tdc0.o_result[112] a_2899_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5919 VGND _092_ a_17415_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5920 tdc0.w_dly_sig[71] tdc0.w_dly_sig_n[69] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5921 VPWR a_30711_6794# net24 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5922 tdc0.w_dly_sig[46] tdc0.w_dly_sig_n[45] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5923 a_30093_7663# a_29559_7669# a_29998_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5924 VGND tdc0.w_dly_sig_n[103] tdc0.w_dly_sig[104] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5925 VPWR a_11839_14191# a_12007_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5926 _072_ a_14045_12353# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X5928 VPWR a_27135_7881# a_27142_7785# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5929 VPWR _055_ a_22917_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X5930 VPWR clknet_4_3_0_clk a_10607_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5931 VGND tdc0.w_dly_sig[9] tdc0.w_dly_sig_n[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5932 VPWR _030_ a_19855_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5933 VGND tdc0.w_dly_sig_n[118] tdc0.w_dly_sig[119] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5934 tdc0.w_dly_sig_n[23] tdc0.w_dly_sig[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5935 tdc0.w_dly_sig[157] tdc0.w_dly_sig_n[155] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5937 VPWR a_11915_9563# a_11831_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5938 a_8895_16367# a_8031_16373# a_8638_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5939 a_10202_2879# a_10034_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5940 VGND a_4279_5461# a_4237_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5941 VGND a_30591_7637# a_30549_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5942 _188_ a_23303_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5943 VPWR tdc0.w_dly_sig[26] a_20421_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5945 VGND a_9263_8573# a_9431_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5946 VGND tdc0.w_dly_sig[51] tdc0.w_dly_sig_n[52] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5947 a_14104_13103# tdc0.o_result[139] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X5949 a_24029_14191# _151_ a_23947_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5950 a_17362_4105# _102_ a_17048_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X5951 a_17967_10159# tdc0.o_result[3] a_18489_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X5952 VPWR _007_ a_12539_6688# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5953 tdc0.w_dly_sig[124] tdc0.w_dly_sig_n[122] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5954 a_24735_3543# a_25026_3433# a_24977_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5955 a_22530_15253# a_22362_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5956 tdc0.w_dly_sig[109] tdc0.w_dly_sig_n[107] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5957 a_3785_11471# tdc0.w_dly_sig[119] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5958 VGND a_4571_7663# a_4739_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5959 a_8565_16367# a_8031_16373# a_8470_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5960 a_27859_5853# a_27639_5865# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X5961 a_15351_7093# _006_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X5963 VPWR a_15354_17023# a_15281_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5964 a_7001_2767# a_6835_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5967 VGND tdc0.w_dly_sig_n[38] tdc0.w_dly_sig[39] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5968 VPWR tdc0.w_dly_sig[1] tdc0.w_dly_sig_n[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5969 a_19798_7093# a_19598_7393# a_19947_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5970 VPWR _060_ a_21327_3543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5971 VGND tdc0.w_dly_sig_n[91] tdc0.w_dly_sig[93] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5972 VPWR a_2290_11583# a_2217_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5973 VPWR a_14045_12353# _072_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X5975 VPWR a_28078_2741# a_28007_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5976 _051_ a_20359_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X5977 tdc0.w_dly_sig_n[89] tdc0.w_dly_sig[89] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5978 a_11973_2223# tdc0.w_dly_sig[166] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5979 a_1512_6031# a_1113_6031# a_1386_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5980 VPWR a_5291_11989# a_5207_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5981 VPWR a_19586_18517# a_19513_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5982 tdc0.w_dly_sig[45] tdc0.w_dly_sig_n[43] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5983 a_20089_8029# _030_ a_20017_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5984 a_19514_3133# a_19267_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5985 VGND a_12254_13103# clknet_4_6_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X5986 a_10677_16911# a_9687_16911# a_10551_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5987 a_20425_12809# _210_ a_20697_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5988 VPWR tdc0.w_dly_sig[6] tdc0.w_dly_sig_n[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5991 VPWR tdc0.w_dly_sig_n[124] tdc0.w_dly_sig[126] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5992 VGND tdc0.w_dly_sig[34] tdc0.w_dly_sig_n[35] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5993 tdc0.o_result[113] a_2163_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5995 VGND tdc0.w_dly_sig[15] tdc0.w_dly_sig_n[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5996 VGND a_4222_3967# a_4180_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5997 a_4655_7663# a_3873_7669# a_4571_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5998 tdc0.w_dly_sig_n[63] tdc0.w_dly_sig[62] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5999 a_10401_2601# a_9411_2229# a_10275_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6000 a_11803_12559# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6002 a_20003_6031# a_19874_6305# a_19583_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6003 a_12851_15101# a_12153_14735# a_12594_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6004 VPWR tdc0.w_dly_sig_n[42] tdc0.w_dly_sig[44] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6005 VPWR tdc0.w_dly_sig[127] tdc0.w_dly_sig_n[127] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6006 VPWR tdc0.w_dly_sig_n[187] tdc0.w_dly_sig[189] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6007 VGND a_23139_859# a_23097_591# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6008 VPWR a_24731_7271# tdc0.o_result[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6011 VGND a_7867_15003# a_7825_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6012 VPWR a_14802_10901# a_14729_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6013 tdc0.w_dly_sig[35] tdc0.w_dly_sig_n[34] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6014 a_20924_1679# a_20525_1679# a_20798_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6015 _205_ a_19058_4719# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X6016 a_6476_7637# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6017 a_3394_3285# a_3226_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6018 VPWR tdc0.w_dly_sig[113] tdc0.w_dly_sig_n[113] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6019 a_30449_4777# a_29902_4521# a_30102_4676# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6020 a_12434_8207# _167_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X6021 a_30423_14191# a_29725_14197# a_30166_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6022 a_26125_1679# a_25578_1953# a_25778_1653# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6023 _056_ a_16547_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6024 a_1995_7485# a_1297_7119# a_1738_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6025 a_12226_2197# a_12058_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6026 VGND _085_ a_8837_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6027 VPWR tdc0.w_dly_sig_n[75] tdc0.w_dly_sig[77] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6028 VGND a_11287_8573# a_11455_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6029 uo_out[1] a_24653_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6030 tdc0.w_dly_sig_n[0] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6031 a_15545_3855# _007_ a_15473_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6032 VPWR a_8327_4373# a_8243_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6033 VGND a_2658_4373# a_2616_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6035 a_7826_12015# a_7553_12021# a_7741_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6036 tdc0.w_dly_sig[177] tdc0.w_dly_sig_n[176] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6037 VPWR _060_ a_21603_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X6038 tdc0.w_dly_sig_n[16] tdc0.w_dly_sig[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6039 VGND tdc0.w_dly_sig_n[46] tdc0.w_dly_sig[48] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6040 _004_ a_21313_13441# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X6041 a_1738_5461# a_1570_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6042 VPWR clknet_4_11_0_clk a_29375_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6043 VGND tdc0.w_dly_sig_n[94] tdc0.w_dly_sig[95] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6044 tdc0.w_dly_sig_n[137] tdc0.w_dly_sig[137] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6045 VGND a_14064_7093# _076_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6047 VPWR tdc0.w_dly_sig[155] tdc0.w_dly_sig_n[156] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6048 VPWR tdc0.w_dly_sig_n[14] tdc0.w_dly_sig[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6049 a_21431_8181# clknet_4_9_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6050 VGND a_17451_14191# a_17619_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6051 a_20359_11471# tdc0.o_result[0] a_20881_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X6052 a_4793_14735# a_4627_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6053 a_16837_11721# _046_ a_16765_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6055 a_10861_13647# a_9871_13647# a_10735_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6056 a_26882_12559# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X6057 tdc0.w_dly_sig[44] tdc0.w_dly_sig_n[43] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6058 a_11865_4765# _026_ a_11793_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6059 a_25318_7093# a_25111_7093# a_25494_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6060 VGND clknet_4_7_0_clk a_14747_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6061 VPWR a_9431_9563# a_9347_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6062 VPWR _008_ a_17876_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X6063 tdc0.w_dly_sig_n[8] tdc0.w_dly_sig[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6064 tdc0.w_dly_sig[193] tdc0.w_dly_sig_n[192] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6065 a_4571_17277# a_3707_16911# a_4314_17023# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6066 VGND a_4314_17023# a_4272_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6067 VPWR _009_ a_17691_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6068 a_4881_2767# a_3891_2767# a_4755_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6069 tdc0.w_dly_sig_n[165] tdc0.w_dly_sig[164] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6070 VGND tdc0.w_dly_sig[192] tdc0.w_dly_sig_n[192] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6072 a_6982_16341# a_6814_16367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6074 tdc0.w_dly_sig[137] tdc0.w_dly_sig_n[136] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6075 VGND tdc0.w_dly_sig_n[109] tdc0.w_dly_sig[110] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6076 VGND a_6027_16091# a_5985_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6077 a_14379_8207# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6079 VPWR tdc0.w_dly_sig[133] tdc0.w_dly_sig_n[133] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6080 tdc0.w_dly_sig[57] tdc0.w_dly_sig_n[55] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6081 a_20417_4373# _184_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X6083 VPWR tdc0.w_dly_sig_n[20] tdc0.w_dly_sig[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6084 VPWR clknet_4_7_0_clk a_11527_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6087 a_26790_11445# a_26583_11445# a_26966_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6088 VPWR _051_ a_23303_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6089 VGND tdc0.w_dly_sig_n[115] tdc0.w_dly_sig[116] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6090 a_4241_17277# a_3707_16911# a_4146_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6091 VPWR a_8638_16341# a_8565_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6092 a_19954_15253# a_19786_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6093 VPWR _097_ a_17481_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X6095 VGND tdc0.w_dly_sig_n[97] tdc0.w_dly_sig[99] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6096 a_27031_13335# a_27127_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6097 tdc0.w_dly_sig[189] tdc0.w_dly_sig_n[187] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6098 VGND a_18935_3543# _061_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X6100 tdc0.w_dly_sig[150] tdc0.w_dly_sig_n[149] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6102 tdc0.w_dly_sig[82] tdc0.w_dly_sig_n[80] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6103 a_10662_14847# a_10494_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6104 tdc0.w_dly_sig_n[71] tdc0.w_dly_sig[71] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6105 VGND a_25410_13103# clknet_4_15_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X6106 VPWR _010_ a_25375_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X6107 a_20733_5853# _030_ a_20661_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6108 VPWR a_30591_15253# a_30507_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6109 VPWR a_12778_5461# a_12705_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6110 tdc0.w_dly_sig[15] tdc0.w_dly_sig_n[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6111 a_20145_7119# a_19591_7093# a_19798_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6112 VGND tdc0.w_dly_sig[48] a_27413_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6113 VPWR _003_ a_18843_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X6114 tdc0.w_dly_sig[167] tdc0.w_dly_sig_n[166] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6115 VGND _055_ a_17220_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X6116 a_11145_1679# tdc0.w_dly_sig[165] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6117 tdc0.w_dly_sig[140] tdc0.w_dly_sig_n[139] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6118 a_16684_9071# _068_ a_16193_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X6119 VPWR tdc0.w_dly_sig[49] tdc0.w_dly_sig_n[50] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6120 tdc0.w_dly_sig[150] tdc0.w_dly_sig_n[148] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6121 tdc0.w_dly_sig[145] tdc0.w_dly_sig_n[143] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6122 a_26203_7271# a_26299_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6123 VGND a_26422_9269# a_26351_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6124 tdc0.w_dly_sig[74] tdc0.w_dly_sig_n[73] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6126 VGND a_1554_6143# a_1512_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6127 a_16175_15975# a_16271_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6128 VGND a_29607_11623# tdc0.o_result[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6129 VPWR a_16791_3035# a_16707_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6130 a_25962_12533# a_25755_12533# a_26138_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6131 a_2582_6575# a_2309_6581# a_2497_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6132 a_16350_8751# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X6133 tdc0.o_result[102] a_5199_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6134 VGND tdc0.w_dly_sig_n[87] tdc0.w_dly_sig[89] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6135 VGND _012_ a_15729_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6136 tdc0.w_dly_sig_n[156] tdc0.w_dly_sig[155] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6137 VPWR _076_ a_14379_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6138 tdc0.w_dly_sig_n[15] tdc0.w_dly_sig[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6139 VGND _178_ a_13722_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X6143 _048_ a_16219_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6144 VGND net5 _006_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X6145 VPWR tdc0.w_dly_sig[8] tdc0.w_dly_sig_n[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6146 a_24170_11721# _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X6148 tdc0.w_dly_sig[51] tdc0.w_dly_sig_n[50] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6149 net2 a_15575_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X6150 tdc0.o_result[102] a_5199_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6151 a_8546_2197# a_8378_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6152 VGND a_22511_4399# a_22679_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6153 a_12537_7983# _023_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X6154 tdc0.w_dly_sig[138] tdc0.w_dly_sig_n[137] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6155 VPWR tdc0.w_dly_sig[126] tdc0.w_dly_sig_n[126] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6156 _173_ a_14922_13897# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X6157 a_24639_13799# a_24735_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6158 VGND a_25111_7093# a_25118_7393# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6159 VPWR _039_ a_15465_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X6160 a_22523_2589# a_22303_2601# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6161 tdc0.o_result[170] a_17159_859# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6162 a_23075_4007# tdc0.o_result[184] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6163 a_24218_15823# a_23903_15975# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6164 VGND a_10627_3035# a_10585_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6165 VPWR a_19947_4007# _176_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6166 VGND clknet_4_2_0_clk a_15759_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6167 VPWR tdc0.w_dly_sig[41] tdc0.w_dly_sig_n[42] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6168 a_27587_2741# a_27871_2741# a_27806_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6169 VGND a_20966_1791# a_20924_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6170 tdc0.w_dly_sig[51] tdc0.w_dly_sig_n[49] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6171 VGND a_20881_11721# uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6172 a_17083_15101# a_16219_14735# a_16826_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6173 VGND _158_ a_19150_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X6174 a_25609_9117# _010_ a_25537_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6175 a_22787_3133# a_21923_2767# a_22530_2879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6176 VGND tdc0.w_dly_sig[161] tdc0.w_dly_sig_n[162] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6177 VGND a_16179_7637# _002_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X6178 VGND tdc0.w_dly_sig[170] tdc0.w_dly_sig_n[170] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6179 tdc0.w_dly_sig[30] tdc0.w_dly_sig_n[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6180 a_29998_8751# a_29725_8757# a_29913_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6182 VGND a_11812_13621# clknet_4_7_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6183 VGND _072_ a_6629_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X6184 tdc0.w_dly_sig_n[133] tdc0.w_dly_sig[133] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6185 a_4797_8207# tdc0.w_dly_sig[133] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6186 VPWR clknet_4_5_0_clk a_8399_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6190 _099_ a_14379_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6191 a_17765_13103# tdc0.o_result[88] a_17681_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6193 tdc0.w_dly_sig[21] tdc0.w_dly_sig_n[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6195 VPWR _003_ a_22891_14423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X6196 a_27639_5865# a_27503_5705# a_27219_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6197 a_25494_7485# a_25247_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6198 VGND a_23634_7637# a_23592_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6199 VGND tdc0.w_dly_sig[60] tdc0.w_dly_sig_n[61] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6200 a_11885_12559# tdc0.o_result[81] a_11803_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6201 tdc0.w_dly_sig[108] tdc0.w_dly_sig_n[107] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6202 VGND a_22852_7093# clknet_4_9_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6203 VGND a_11582_6143# a_11540_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6204 VPWR tdc0.w_dly_sig_n[78] tdc0.w_dly_sig[79] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6205 VPWR _056_ a_19899_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6206 a_4146_7663# a_3707_7669# a_4061_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6207 tdc0.w_dly_sig[69] tdc0.w_dly_sig_n[67] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6208 a_21223_2045# a_20525_1679# a_20966_1791# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6209 tdc0.w_dly_sig_n[123] tdc0.w_dly_sig[123] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6210 VGND net1 tdc0.w_dly_sig_n[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6211 tdc0.w_dly_sig[175] tdc0.w_dly_sig_n[174] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6212 VGND tdc0.w_dly_sig[121] tdc0.w_dly_sig_n[121] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6213 VPWR a_19183_2197# a_19099_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6214 tdc0.w_dly_sig[174] tdc0.w_dly_sig_n[173] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6215 VGND tdc0.w_dly_sig[181] tdc0.w_dly_sig_n[181] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6216 VPWR tdc0.w_dly_sig_n[21] tdc0.w_dly_sig[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6217 a_13349_16373# a_13183_16373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6218 VPWR _064_ a_19967_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6219 a_17451_2223# a_16753_2229# a_17194_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6221 a_9263_14013# a_8399_13647# a_9006_13759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6222 tdc0.w_dly_sig_n[105] tdc0.w_dly_sig[104] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6225 VGND a_22466_12533# a_22395_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6226 VGND tdc0.w_dly_sig_n[189] tdc0.w_dly_sig[191] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6227 tdc0.w_dly_sig[2] tdc0.w_dly_sig_n[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6228 tdc0.w_dly_sig[4] tdc0.w_dly_sig_n[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6229 a_16850_13423# _052_ a_17096_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X6231 VPWR a_4314_17023# a_4241_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6232 tdc0.w_dly_sig_n[115] tdc0.w_dly_sig[114] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6234 tdc0.w_dly_sig[170] tdc0.w_dly_sig_n[168] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6235 VGND a_15837_8181# _014_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X6236 VPWR tdc0.o_result[95] a_18703_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6237 a_5115_15279# a_4333_15285# a_5031_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6238 a_6771_13103# a_5989_13109# a_6687_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6239 VPWR a_19497_5089# _137_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X6240 tdc0.w_dly_sig[67] tdc0.w_dly_sig_n[65] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6241 a_12705_5487# a_12171_5493# a_12610_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6242 a_15325_3677# _056_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X6243 tdc0.w_dly_sig[158] tdc0.w_dly_sig_n[156] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6244 a_15085_3855# _038_ a_15013_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6245 a_1995_5487# a_1297_5493# a_1738_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6247 VPWR tdc0.w_dly_sig_n[146] tdc0.w_dly_sig[147] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6248 VPWR tdc0.w_dly_sig[40] tdc0.w_dly_sig_n[40] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6249 VPWR clknet_4_3_0_clk a_10883_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6250 a_8399_10633# _027_ a_8481_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6252 VGND a_5234_14847# a_5192_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6253 _077_ a_14379_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X6254 clknet_4_3_0_clk a_10506_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6255 tdc0.w_dly_sig[14] tdc0.w_dly_sig_n[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6256 VPWR a_15427_18365# a_15595_18267# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6257 VPWR tdc0.w_dly_sig[63] tdc0.w_dly_sig_n[64] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6258 VGND tdc0.w_dly_sig_n[177] tdc0.w_dly_sig[178] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6260 VGND tdc0.w_dly_sig_n[169] tdc0.w_dly_sig[170] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6261 a_21718_5487# a_21445_5493# a_21633_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6262 a_19333_18543# tdc0.w_dly_sig[56] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6263 tdc0.o_result[123] a_7591_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6264 VPWR tdc0.w_dly_sig[71] tdc0.w_dly_sig_n[72] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6265 a_23947_12015# _152_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6266 a_27087_8207# a_26951_8181# a_26667_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6267 a_23700_9839# _126_ a_23598_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6268 VPWR clknet_4_2_0_clk a_9411_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6269 VGND tdc0.w_dly_sig[119] tdc0.w_dly_sig_n[119] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6270 tdc0.w_dly_sig[129] tdc0.w_dly_sig_n[127] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6271 VGND a_24283_4917# a_24290_5217# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6273 a_11405_4765# _026_ a_11333_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6274 a_16665_5487# net6 a_17023_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6275 a_12935_11837# a_12153_11471# a_12851_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6276 a_17383_5095# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X6277 VGND tdc0.w_dly_sig_n[162] tdc0.w_dly_sig[164] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6278 VGND tdc0.w_dly_sig_n[171] tdc0.w_dly_sig[173] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6279 VPWR a_30591_14165# a_30507_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6280 a_4498_2879# a_4330_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6281 VGND tdc0.w_dly_sig[173] tdc0.w_dly_sig_n[174] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6282 a_13889_14557# _022_ a_13817_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6283 tdc0.w_dly_sig_n[120] tdc0.w_dly_sig[119] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6284 a_15427_18365# a_14729_17999# a_15170_18111# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6286 a_17477_16911# a_16923_16885# a_17130_16885# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6287 VPWR tdc0.w_dly_sig[45] tdc0.w_dly_sig_n[45] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6288 VGND clknet_4_6_0_clk a_11987_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6289 a_19685_2767# a_19138_3041# a_19338_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6290 VPWR _076_ a_12999_12128# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6291 VGND tdc0.w_dly_sig[33] a_20421_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6292 a_22987_6807# a_23271_6793# a_23206_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6293 VGND clknet_0_clk a_7378_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6294 VGND a_28687_16599# tdc0.o_result[46] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6295 tdc0.w_dly_sig_n[107] tdc0.w_dly_sig[106] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6296 VGND _048_ a_16850_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X6297 tdc0.w_dly_sig[156] tdc0.w_dly_sig_n[154] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6298 _010_ a_17691_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6299 tdc0.o_result[105] a_3819_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6300 a_15009_15823# tdc0.w_dly_sig[68] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6301 tdc0.w_dly_sig[40] tdc0.w_dly_sig_n[39] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6302 tdc0.w_dly_sig_n[121] tdc0.w_dly_sig[120] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6303 a_24197_12015# _170_ a_24469_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6304 VPWR tdc0.w_dly_sig_n[2] tdc0.w_dly_sig[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6305 a_24131_9295# _090_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6307 VGND a_17187_13799# _049_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X6308 _201_ a_13722_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X6309 _156_ a_12999_12128# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6310 VGND tdc0.w_dly_sig_n[18] tdc0.w_dly_sig[20] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6312 tdc0.o_result[13] a_30591_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6313 a_5989_5493# a_5823_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6314 VPWR a_12007_6299# a_11923_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6315 tdc0.w_dly_sig[89] tdc0.w_dly_sig_n[88] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6316 VPWR clknet_4_2_0_clk a_15759_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6317 a_16271_15797# a_16555_15797# a_16490_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6318 VPWR _026_ a_11159_8864# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6319 VGND a_29274_16644# a_29203_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6320 VGND a_27043_4617# a_27050_4521# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6321 a_20273_5853# _030_ a_20201_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6322 tdc0.w_dly_sig_n[105] tdc0.w_dly_sig[105] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6323 VPWR a_19807_12559# _012_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6324 VPWR a_18130_591# a_18236_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X6325 VGND clknet_4_5_0_clk a_3707_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6326 a_9347_8573# a_8565_8207# a_9263_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6327 VPWR tdc0.w_dly_sig[97] tdc0.w_dly_sig_n[98] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6328 a_24029_14191# _014_ a_24113_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6330 clknet_4_2_0_clk a_11260_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6331 a_19341_9545# _185_ a_19245_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6332 a_11329_7663# tdc0.w_dly_sig[138] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6333 a_25931_9269# a_26215_9269# a_26150_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6334 a_17578_18365# a_17139_17999# a_17493_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6335 VGND tdc0.w_dly_sig[35] tdc0.w_dly_sig_n[36] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6336 VPWR a_20499_5719# _196_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6337 VGND clk a_16210_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6338 clknet_4_12_0_clk a_21380_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6340 a_27767_13469# a_27547_13481# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6341 a_6909_7119# a_6743_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6342 VGND a_16210_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6343 VGND clknet_0_clk a_6550_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6344 a_1995_7485# a_1131_7119# a_1738_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6345 a_11858_1109# a_11690_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6346 VPWR _068_ a_20709_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X6347 VGND a_21787_2455# tdc0.o_result[181] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6348 VPWR tdc0.w_dly_sig_n[145] tdc0.w_dly_sig[146] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6350 a_4272_8041# a_3873_7669# a_4146_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6351 tdc0.o_result[157] a_6671_4123# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6352 tdc0.w_dly_sig_n[147] tdc0.w_dly_sig[146] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6353 VPWR tdc0.w_dly_sig[75] tdc0.w_dly_sig_n[75] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6354 a_15293_4943# a_15023_5309# a_15203_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X6355 a_2405_4399# tdc0.w_dly_sig[153] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6356 tdc0.w_dly_sig_n[59] tdc0.w_dly_sig[58] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6357 VGND tdc0.w_dly_sig[170] tdc0.w_dly_sig_n[171] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6358 a_21949_3677# _056_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X6359 a_10175_4399# a_9393_4405# a_10091_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6361 VPWR a_9006_13759# a_8933_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6362 VGND _017_ a_20992_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X6363 a_24186_16341# a_24018_16367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6364 VPWR a_12254_13103# clknet_4_6_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6365 VPWR tdc0.w_dly_sig[184] a_24837_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6366 a_23465_9129# a_22475_8757# a_23339_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6367 a_14686_8751# _033_ a_14437_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X6368 tdc0.w_dly_sig[155] tdc0.w_dly_sig_n[154] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6369 a_5249_9129# a_4259_8757# a_5123_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6370 VGND tdc0.w_dly_sig[46] tdc0.w_dly_sig_n[46] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6371 VPWR clknet_4_1_0_clk a_8399_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6372 a_19497_5089# _135_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X6373 VGND clknet_4_0_0_clk a_3615_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6375 _200_ a_13643_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6376 VGND tdc0.w_dly_sig[183] tdc0.w_dly_sig_n[184] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6377 VGND _176_ a_19773_9441# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X6378 a_6227_3133# a_5363_2767# a_5970_2879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6379 VGND tdc0.w_dly_sig_n[164] tdc0.w_dly_sig[166] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6380 a_18659_7895# _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X6381 VGND tdc0.w_dly_sig_n[172] tdc0.w_dly_sig[174] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6382 VPWR a_19735_859# a_19651_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6383 a_11965_14569# a_10975_14197# a_11839_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6384 tdc0.w_dly_sig[120] tdc0.w_dly_sig_n[118] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6385 VGND tdc0.w_dly_sig_n[4] tdc0.w_dly_sig[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6386 a_29611_4631# a_29902_4521# a_29853_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6387 a_21380_14165# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6388 VPWR tdc0.w_dly_sig[41] tdc0.w_dly_sig_n[41] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6389 a_18888_4399# tdc0.o_result[151] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X6390 tdc0.w_dly_sig[25] tdc0.w_dly_sig_n[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6391 a_27123_5719# a_27219_5719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6392 tdc0.w_dly_sig_n[22] tdc0.w_dly_sig[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6394 a_15101_7637# _022_ a_15347_8001# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6395 a_19947_4007# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X6396 VGND a_16734_18517# a_16692_18921# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6397 _063_ a_16587_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X6398 VPWR clknet_0_clk a_25428_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6399 a_11965_8041# a_10975_7669# a_11839_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6400 a_5349_15823# tdc0.w_dly_sig[104] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6401 _105_ a_17218_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X6402 a_2658_4373# a_2490_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6403 tdc0.w_dly_sig_n[31] tdc0.w_dly_sig[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6404 _083_ a_14379_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X6405 a_3049_15279# tdc0.w_dly_sig[105] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6407 clknet_4_10_0_clk a_25428_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6408 a_19802_11293# a_19487_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6410 VGND tdc0.w_dly_sig[54] tdc0.w_dly_sig_n[55] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6411 VPWR tdc0.w_dly_sig[23] tdc0.w_dly_sig_n[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6412 a_21787_8207# a_21567_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6413 VGND _116_ a_14437_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X6414 tdc0.w_dly_sig[107] tdc0.w_dly_sig_n[106] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6415 tdc0.w_dly_sig[80] tdc0.w_dly_sig_n[79] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6416 _102_ a_15391_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6417 a_7399_6031# a_7263_6005# a_6979_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6418 VPWR tdc0.w_dly_sig[105] tdc0.w_dly_sig_n[106] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6419 VPWR tdc0.w_dly_sig_n[140] tdc0.w_dly_sig[142] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6421 tdc0.o_result[154] a_3819_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6422 tdc0.w_dly_sig[4] tdc0.w_dly_sig_n[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6423 clknet_0_clk a_16210_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6424 a_16753_2229# a_16587_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6425 a_30239_9839# a_29375_9845# a_29982_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6426 a_16991_18543# a_16293_18549# a_16734_18517# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6427 VPWR a_2750_6549# a_2677_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6428 VGND tdc0.w_dly_sig[52] tdc0.w_dly_sig_n[52] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6429 a_3651_3311# a_2787_3317# a_3394_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6430 a_17957_3855# tdc0.o_result[172] a_17875_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6431 a_14428_9839# _074_ a_14326_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X6432 VGND a_18489_9839# uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6433 a_17117_18921# a_16127_18549# a_16991_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6434 VGND tdc0.w_dly_sig[145] tdc0.w_dly_sig_n[145] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6435 a_17688_12335# tdc0.o_result[11] a_17498_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X6436 VGND _000_ a_18059_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6437 VPWR tdc0.w_dly_sig_n[63] tdc0.w_dly_sig[64] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6440 a_28503_12247# a_28599_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6441 a_1301_6031# tdc0.w_dly_sig[110] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6442 a_9390_7485# a_9117_7119# a_9305_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6443 a_16179_7637# net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X6444 a_14064_7093# _013_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6445 a_7365_16745# a_6375_16373# a_7239_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6446 clknet_4_4_0_clk a_6550_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6447 a_2915_4399# a_2217_4405# a_2658_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6449 _046_ a_13722_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X6450 VPWR a_19855_7895# _115_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6451 VPWR tdc0.o_result[30] a_24436_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X6452 VPWR a_22955_3035# a_22871_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
R15 VPWR tt_um_hpretl_tt06_tdc_v1_11.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6454 a_7090_10749# a_6651_10383# a_7005_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6455 uo_out[5] a_24469_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6457 VPWR ui_in[0] a_30347_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6458 a_5050_6143# a_4882_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6459 a_24018_16367# a_23579_16373# a_23933_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6460 _206_ a_15575_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X6461 a_25665_7119# a_25118_7393# a_25318_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6462 a_26663_4631# a_26759_4631# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6463 tdc0.o_result[148] a_4555_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6464 a_12999_8867# _169_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X6465 VGND ui_in[4] a_16219_1143# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6466 a_5433_8207# a_4443_8207# a_5307_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6467 a_9297_17833# a_8307_17461# a_9171_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6469 a_20713_1679# tdc0.w_dly_sig[179] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6470 VPWR clknet_0_clk a_10506_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6471 tdc0.w_dly_sig_n[119] tdc0.w_dly_sig[118] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6472 VPWR tdc0.w_dly_sig_n[42] tdc0.w_dly_sig[43] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6473 VGND tdc0.w_dly_sig_n[101] tdc0.w_dly_sig[103] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6474 tdc0.w_dly_sig[29] tdc0.w_dly_sig_n[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6475 tdc0.w_dly_sig_n[34] tdc0.w_dly_sig[33] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6476 a_9853_16911# a_9687_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6477 tdc0.w_dly_sig_n[48] tdc0.w_dly_sig[48] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6478 a_21031_13675# _003_ a_20945_13675# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X6479 a_7626_10901# a_7458_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6481 VPWR tdc0.w_dly_sig_n[32] tdc0.w_dly_sig[33] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6482 VGND clknet_4_5_0_clk a_4627_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6483 a_2432_10217# a_2033_9845# a_2306_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6484 VPWR tdc0.w_dly_sig[186] tdc0.w_dly_sig_n[186] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6485 VPWR tdc0.w_dly_sig[81] tdc0.w_dly_sig_n[81] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6486 a_5805_11721# tdc0.o_result[118] a_5721_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6487 a_15553_2601# a_14563_2229# a_15427_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6490 VPWR tdc0.w_dly_sig[27] tdc0.w_dly_sig_n[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6491 a_23381_7663# tdc0.w_dly_sig[27] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6493 VPWR clknet_4_12_0_clk a_21923_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6494 VPWR tdc0.w_dly_sig_n[110] tdc0.w_dly_sig[112] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6495 VPWR tdc0.w_dly_sig[25] a_23825_6953# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6496 a_14250_17429# a_14082_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6497 VPWR tdc0.w_dly_sig[3] a_24009_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6498 tdc0.w_dly_sig_n[97] tdc0.w_dly_sig[96] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6499 a_15354_17023# a_15186_17277# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6500 a_7458_10927# a_7185_10933# a_7373_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6501 tdc0.w_dly_sig[54] tdc0.w_dly_sig_n[52] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6502 _012_ a_19807_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6503 VGND tdc0.w_dly_sig[27] tdc0.w_dly_sig_n[28] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6504 VGND tdc0.w_dly_sig[11] a_27505_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6505 VGND clknet_4_4_0_clk a_7019_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6506 VPWR tdc0.w_dly_sig_n[128] tdc0.w_dly_sig[129] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6507 a_28783_16599# a_29074_16489# a_29025_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6508 VGND _003_ a_21399_13441# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X6509 a_2673_12559# a_1683_12559# a_2547_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6511 a_24511_15279# tdc0.o_result[49] a_24309_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6512 VPWR tdc0.w_dly_sig_n[21] tdc0.w_dly_sig[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6513 VGND a_17231_4399# _043_ VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6514 VPWR tdc0.w_dly_sig[137] tdc0.w_dly_sig_n[137] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6515 a_4866_8725# a_4698_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6516 a_29266_12015# a_29019_12393# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6517 a_21914_11204# a_21714_11049# a_22063_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6518 a_21883_2455# a_22167_2441# a_22102_2589# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6519 VPWR a_16762_15797# a_16691_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6520 VGND a_21759_15003# a_21717_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6521 VPWR clknet_4_0_0_clk a_3615_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6522 VGND _043_ a_13153_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6523 tdc0.w_dly_sig[125] tdc0.w_dly_sig_n[124] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6525 a_24385_14511# tdc0.o_result[45] a_23947_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6526 VGND a_16635_4007# _168_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X6527 VGND tdc0.w_dly_sig_n[116] tdc0.w_dly_sig[118] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6529 tdc0.w_dly_sig[119] tdc0.w_dly_sig_n[118] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6530 VPWR a_20039_5719# _136_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6531 tdc0.w_dly_sig_n[166] tdc0.w_dly_sig[166] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6532 tdc0.w_dly_sig[115] tdc0.w_dly_sig_n[113] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6533 VPWR tdc0.w_dly_sig[175] tdc0.w_dly_sig_n[175] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6534 VGND tdc0.w_dly_sig[144] tdc0.w_dly_sig_n[144] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6535 VGND _113_ a_15943_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6536 a_2179_10927# a_1481_10933# a_1922_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6537 tdc0.w_dly_sig[134] tdc0.w_dly_sig_n[132] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6538 a_21707_11145# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6539 tdc0.o_result[161] a_8971_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6540 VPWR a_21886_5461# a_21813_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6541 a_12023_18543# a_11325_18549# a_11766_18517# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
R16 VGND uio_out[6] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6542 _152_ a_23947_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X6543 a_6998_3311# a_6725_3317# a_6913_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6545 a_8803_2223# a_7939_2229# a_8546_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6547 _210_ a_19255_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6548 tdc0.w_dly_sig_n[178] tdc0.w_dly_sig[178] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6549 VGND tdc0.w_dly_sig[129] tdc0.w_dly_sig_n[129] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6550 a_26939_11471# a_26719_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6551 a_24241_5309# a_23903_5095# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6552 a_21638_8181# a_21438_8481# a_21787_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6554 a_20096_14569# a_19697_14197# a_19970_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6555 a_21489_3677# _056_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X6556 a_15002_18365# a_14563_17999# a_14917_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6557 a_15465_12015# tdc0.o_result[38] a_15381_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6558 a_24344_8457# _031_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X6559 VPWR tdc0.w_dly_sig[166] tdc0.w_dly_sig_n[167] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6560 tdc0.w_dly_sig_n[18] tdc0.w_dly_sig[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6561 tdc0.w_dly_sig_n[2] tdc0.w_dly_sig[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6562 a_26903_16911# a_26767_16885# a_26483_16885# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6563 a_2915_4399# a_2051_4405# a_2658_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6564 _014_ a_15837_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.247 ps=2.06 w=0.65 l=0.15
X6565 a_18127_10927# tdc0.o_result[2] a_17937_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X6566 VGND a_12851_16189# a_13019_16091# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6570 VGND a_20074_11204# a_20003_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6571 a_24919_3829# a_25210_4129# a_25161_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6572 VPWR tdc0.w_dly_sig[125] tdc0.w_dly_sig_n[126] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6573 a_7124_3689# a_6725_3317# a_6998_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6574 VGND _075_ a_14563_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6575 a_6913_14191# tdc0.w_dly_sig[124] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6576 a_13153_3677# _025_ a_13081_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6577 VGND tdc0.w_dly_sig[42] a_26217_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6578 tdc0.o_result[90] a_14675_17429# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6579 VGND tdc0.w_dly_sig[109] tdc0.w_dly_sig_n[109] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6580 a_13717_2767# a_13551_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6581 tdc0.w_dly_sig_n[27] tdc0.w_dly_sig[27] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6582 a_9765_2223# tdc0.w_dly_sig[164] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6583 VPWR a_27710_5764# a_27639_5865# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6584 tdc0.o_result[111] a_2715_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6585 a_20697_12809# _210_ a_20425_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6586 VPWR net6 a_17773_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X6587 tdc0.w_dly_sig[85] tdc0.w_dly_sig_n[84] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6588 VPWR tdc0.w_dly_sig[162] tdc0.w_dly_sig_n[162] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6589 a_25069_11837# a_24731_11623# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6590 VPWR clknet_4_12_0_clk a_17783_16373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6591 VGND tdc0.w_dly_sig[182] tdc0.w_dly_sig_n[182] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6592 VPWR tdc0.o_result[152] a_13735_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6594 VGND _047_ a_13897_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6595 VGND tdc0.w_dly_sig_n[160] tdc0.w_dly_sig[162] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6597 a_29729_12559# tdc0.w_dly_sig[44] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6598 VGND tdc0.w_dly_sig[98] tdc0.w_dly_sig_n[99] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6599 tdc0.w_dly_sig[97] tdc0.w_dly_sig_n[96] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6600 VPWR clknet_4_3_0_clk a_10975_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6601 VPWR tdc0.w_dly_sig_n[31] tdc0.w_dly_sig[32] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6602 VGND tdc0.w_dly_sig[83] tdc0.w_dly_sig_n[83] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6603 VPWR a_21327_11159# tdc0.o_result[34] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6604 a_15538_12671# a_15370_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6605 tdc0.w_dly_sig_n[169] tdc0.w_dly_sig[168] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6606 tdc0.w_dly_sig[52] tdc0.w_dly_sig_n[50] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6607 tdc0.w_dly_sig_n[171] tdc0.w_dly_sig[171] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6608 VGND tdc0.w_dly_sig[43] a_29437_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6609 VGND tdc0.w_dly_sig[78] tdc0.w_dly_sig_n[79] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6610 VGND a_7263_6005# a_7270_6305# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6611 a_23745_16373# a_23579_16373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6612 VPWR tdc0.w_dly_sig[20] tdc0.w_dly_sig_n[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6613 VGND a_15795_12925# a_15963_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6614 _195_ a_14931_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6615 VPWR tdc0.w_dly_sig_n[137] tdc0.w_dly_sig[138] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6616 a_3141_14191# tdc0.w_dly_sig[106] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6618 a_18130_591# a_17953_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6619 a_25375_15975# a_25471_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6620 VGND net1 tdc0.w_dly_sig_n[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6621 tdc0.w_dly_sig_n[89] tdc0.w_dly_sig[88] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6622 a_8638_3285# a_8470_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6623 a_11957_12559# _034_ a_11885_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6624 VPWR tdc0.w_dly_sig_n[77] tdc0.w_dly_sig[78] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6625 a_19890_13103# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X6626 tdc0.w_dly_sig_n[113] tdc0.w_dly_sig[112] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6627 VPWR a_20011_18517# a_19927_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6628 _003_ a_18703_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X6630 tdc0.w_dly_sig_n[49] tdc0.w_dly_sig[49] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6631 a_4333_7119# a_4167_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6632 tdc0.w_dly_sig[95] tdc0.w_dly_sig_n[94] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6633 a_6725_3317# a_6559_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6634 a_2221_9839# tdc0.w_dly_sig[113] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6635 tdc0.w_dly_sig_n[28] tdc0.w_dly_sig[28] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6636 tdc0.w_dly_sig[117] tdc0.w_dly_sig_n[115] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6637 a_23903_5095# a_23999_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6638 VPWR a_14250_15253# a_14177_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6639 VPWR a_14158_2879# a_14085_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6640 VPWR _051_ a_12171_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6642 VPWR clknet_4_5_0_clk a_4627_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6643 a_11582_14165# a_11414_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6645 a_29090_12292# a_28883_12233# a_29266_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6646 a_5077_10383# tdc0.o_result[150] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6649 VPWR a_5123_8751# a_5291_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6650 VPWR tdc0.w_dly_sig[79] tdc0.w_dly_sig_n[80] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6651 VGND _131_ a_5823_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6652 a_19974_7485# a_19727_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6653 tdc0.w_dly_sig_n[180] tdc0.w_dly_sig[179] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6654 a_15801_7369# a_15731_7271# _006_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X6655 VPWR a_19395_7895# _158_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6656 a_21813_5487# a_21279_5493# a_21718_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6657 VPWR a_6395_3035# a_6311_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6658 a_13817_4765# tdc0.o_result[152] a_13735_4512# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6659 VPWR tdc0.w_dly_sig[38] tdc0.w_dly_sig_n[39] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6661 a_23269_9813# _128_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X6662 a_6541_16373# a_6375_16373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6663 VGND tdc0.w_dly_sig[124] tdc0.w_dly_sig_n[125] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6664 _035_ a_14255_6835# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6665 tdc0.w_dly_sig[110] tdc0.w_dly_sig_n[109] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6666 a_29019_12393# a_28883_12233# a_28599_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6667 a_2673_11471# a_1683_11471# a_2547_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6668 _010_ a_17691_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6669 _064_ _010_ a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6670 VPWR _023_ a_8481_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6671 a_8895_3311# a_8197_3317# a_8638_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6672 VGND a_16547_4373# _056_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X6673 tdc0.w_dly_sig_n[60] tdc0.w_dly_sig[59] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6674 tdc0.w_dly_sig[72] tdc0.w_dly_sig_n[71] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6675 VGND tdc0.w_dly_sig_n[132] tdc0.w_dly_sig[133] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6676 a_5560_15823# a_5161_15823# a_5434_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6677 a_4471_4399# a_3689_4405# a_4387_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6678 a_1570_7485# a_1131_7119# a_1485_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6679 VGND a_27411_13321# a_27418_13225# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6680 a_22273_591# a_22107_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6681 VPWR a_18843_13335# _140_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6682 VGND clknet_4_0_0_clk a_5363_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6683 a_15837_8181# _002_ a_16083_8235# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6684 tdc0.w_dly_sig[56] tdc0.w_dly_sig_n[54] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6685 VPWR a_2347_10901# a_2263_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6686 a_9673_9839# tdc0.w_dly_sig[79] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6687 tdc0.w_dly_sig[99] tdc0.w_dly_sig_n[97] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6688 a_8473_17461# a_8307_17461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6689 VGND a_2547_12925# a_2715_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6690 tdc0.w_dly_sig[27] tdc0.w_dly_sig_n[26] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6691 tdc0.w_dly_sig[85] tdc0.w_dly_sig_n[83] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6692 VGND a_27043_3829# a_27050_4129# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6693 a_23137_17455# a_22799_17687# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6694 tdc0.w_dly_sig[135] tdc0.w_dly_sig_n[134] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6695 a_17066_9545# _033_ a_16986_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X6697 a_21985_8207# a_21431_8181# a_21638_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6698 tdc0.o_result[157] a_6671_4123# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6699 a_25891_4943# a_25762_5217# a_25471_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6700 a_16941_14191# tdc0.w_dly_sig[71] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6701 VGND tdc0.w_dly_sig_n[5] tdc0.w_dly_sig[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6702 a_11690_1135# a_11251_1141# a_11605_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6703 VGND tdc0.w_dly_sig[42] tdc0.w_dly_sig_n[43] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6704 VPWR a_30407_9813# a_30323_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6705 VPWR clknet_4_5_0_clk a_5823_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6706 VGND tdc0.w_dly_sig[10] tdc0.w_dly_sig_n[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6707 _018_ a_17503_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X6708 tdc0.w_dly_sig_n[114] tdc0.w_dly_sig[113] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6709 tdc0.w_dly_sig[171] tdc0.w_dly_sig_n[170] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6710 a_16937_17455# a_16403_17461# a_16842_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6711 a_25247_11471# a_25118_11745# a_24827_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6712 a_9581_4399# tdc0.w_dly_sig[142] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6713 tdc0.w_dly_sig_n[64] tdc0.w_dly_sig[63] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6714 a_17685_12559# _072_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X6715 a_24597_3855# _050_ a_24525_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6716 tdc0.w_dly_sig_n[50] tdc0.w_dly_sig[49] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6717 VGND tdc0.w_dly_sig_n[57] tdc0.w_dly_sig[59] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6718 a_12483_2223# a_11785_2229# a_12226_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6719 VPWR a_12483_2223# a_12651_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6720 tdc0.w_dly_sig_n[143] tdc0.w_dly_sig[142] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6721 a_11766_18517# a_11598_18543# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6722 a_12134_15253# a_11966_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6723 a_16025_10633# _133_ a_15943_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6724 tdc0.w_dly_sig[142] tdc0.w_dly_sig_n[140] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6725 _065_ a_16713_8235# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X6726 tdc0.w_dly_sig[70] tdc0.w_dly_sig_n[69] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6727 tdc0.w_dly_sig[168] tdc0.w_dly_sig_n[167] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6728 VGND a_16175_15975# tdc0.o_result[64] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6729 a_22125_2223# a_21787_2455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6730 tdc0.w_dly_sig[188] tdc0.w_dly_sig_n[186] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6731 VPWR tdc0.w_dly_sig[93] tdc0.w_dly_sig_n[94] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6732 a_13119_5487# a_12337_5493# a_13035_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6733 tdc0.o_result[76] a_15227_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6734 a_6430_5461# a_6262_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6735 VPWR tdc0.w_dly_sig_n[12] tdc0.w_dly_sig[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6736 tdc0.w_dly_sig_n[88] tdc0.w_dly_sig[87] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6737 VPWR tdc0.w_dly_sig[94] tdc0.w_dly_sig_n[94] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6739 VGND a_8159_4399# a_8327_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6740 VPWR clknet_4_6_0_clk a_9871_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6741 tdc0.w_dly_sig_n[29] tdc0.w_dly_sig[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6742 tdc0.w_dly_sig[118] tdc0.w_dly_sig_n[116] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6743 a_13717_2767# a_13551_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6744 VPWR _030_ a_20499_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X6745 a_11598_18543# a_11325_18549# a_11513_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6746 a_6909_7119# a_6743_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6747 tdc0.w_dly_sig_n[177] tdc0.w_dly_sig[176] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6748 VGND clknet_4_1_0_clk a_2235_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6749 tdc0.w_dly_sig_n[160] tdc0.w_dly_sig[159] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6750 a_7645_11721# tdc0.o_result[98] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6751 a_16913_8001# net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X6752 tdc0.w_dly_sig_n[123] tdc0.w_dly_sig[122] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6753 VPWR tdc0.w_dly_sig[108] tdc0.w_dly_sig_n[109] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6755 VPWR tdc0.w_dly_sig_n[150] tdc0.w_dly_sig[151] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6756 uo_out[0] a_20881_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6757 tdc0.w_dly_sig_n[58] tdc0.w_dly_sig[57] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6758 VPWR tdc0.w_dly_sig_n[150] tdc0.w_dly_sig[152] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6759 a_1849_13647# a_1683_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6761 VGND tdc0.w_dly_sig[118] tdc0.w_dly_sig_n[118] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6762 a_12434_8207# _168_ a_12680_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X6763 a_12594_14847# a_12426_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6764 VGND a_22852_7093# clknet_4_9_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6765 VPWR tdc0.w_dly_sig[164] tdc0.w_dly_sig_n[165] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6766 a_14085_3133# a_13551_2767# a_13990_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6768 a_18935_3543# tdc0.o_result[176] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6769 VPWR clknet_4_11_0_clk a_29559_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6770 a_29803_5705# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6771 a_5123_8751# a_4259_8757# a_4866_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6772 a_15519_16189# a_14821_15823# a_15262_15935# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6773 VPWR a_23903_15975# tdc0.o_result[49] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6774 a_4425_12021# a_4259_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6775 VGND tdc0.w_dly_sig[10] tdc0.w_dly_sig_n[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6776 VGND tdc0.w_dly_sig[7] a_29437_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6777 tdc0.w_dly_sig_n[61] tdc0.w_dly_sig[60] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6778 a_30239_9839# a_29541_9845# a_29982_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6779 VPWR tdc0.w_dly_sig_n[59] tdc0.w_dly_sig[60] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6781 a_4203_10927# a_3505_10933# a_3946_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6783 VGND tdc0.w_dly_sig[56] tdc0.w_dly_sig_n[56] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6784 a_10041_16911# tdc0.w_dly_sig[96] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6785 VGND a_23351_14423# _146_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X6786 VPWR a_24363_4007# _108_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6787 a_19899_8751# _010_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X6788 a_11322_9661# a_11049_9295# a_11237_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6789 VGND clknet_4_8_0_clk a_20175_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6790 a_19931_4737# _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X6791 VGND tdc0.w_dly_sig[131] tdc0.w_dly_sig_n[131] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6792 VGND a_16826_14847# a_16784_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6793 tdc0.w_dly_sig[45] tdc0.w_dly_sig_n[44] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6794 VGND a_5475_8475# a_5433_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6795 a_2122_13103# a_1683_13109# a_2037_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6796 a_12526_9295# _087_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X6797 VGND a_27526_10116# a_27455_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6798 VGND tdc0.w_dly_sig[82] tdc0.w_dly_sig_n[83] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6799 tdc0.w_dly_sig[118] tdc0.w_dly_sig_n[117] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6800 VPWR a_25755_4917# a_25762_5217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6801 VPWR a_21380_14165# clknet_4_12_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6802 VGND tdc0.w_dly_sig_n[53] tdc0.w_dly_sig[55] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6803 a_27526_12292# a_27326_12137# a_27675_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6804 _088_ a_11251_4512# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6805 a_11141_14197# a_10975_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6806 a_10957_1679# a_10791_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6807 tdc0.w_dly_sig[9] tdc0.w_dly_sig_n[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6809 tdc0.o_result[97] a_9063_16341# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6810 a_25471_15797# a_25755_15797# a_25690_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6811 tdc0.w_dly_sig[8] tdc0.w_dly_sig_n[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6813 a_7423_14191# a_6559_14197# a_7166_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6814 VGND a_30166_7637# a_30124_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6815 a_6177_4399# tdc0.w_dly_sig[152] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6816 tdc0.w_dly_sig_n[12] tdc0.w_dly_sig[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6817 tdc0.o_result[97] a_9063_16341# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6818 tdc0.w_dly_sig[176] tdc0.w_dly_sig_n[175] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6819 a_23309_3855# _050_ a_23237_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6820 VGND a_7407_16341# a_7365_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6821 tdc0.w_dly_sig_n[50] tdc0.w_dly_sig[50] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6822 a_6687_13103# a_5823_13109# a_6430_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6824 VGND _145_ a_18059_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X6825 a_27307_9117# a_27087_9129# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6826 a_15143_10927# a_14361_10933# a_15059_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6827 tdc0.w_dly_sig_n[184] tdc0.w_dly_sig[184] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6828 a_11598_18543# a_11159_18549# a_11513_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6829 tdc0.o_result[150] a_3175_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6830 a_1696_7119# a_1297_7119# a_1570_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6832 VPWR tdc0.w_dly_sig[17] tdc0.w_dly_sig_n[17] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6833 VGND a_30711_6794# net24 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6834 a_7093_14191# a_6559_14197# a_6998_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6835 a_18935_3543# tdc0.o_result[176] a_19169_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6836 VGND a_17139_8759# _054_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X6837 VPWR clknet_4_8_0_clk a_16587_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6838 VGND tdc0.w_dly_sig_n[86] tdc0.w_dly_sig[88] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6839 tdc0.w_dly_sig_n[111] tdc0.w_dly_sig[110] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6841 VPWR a_8971_2197# a_8887_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6842 VPWR tdc0.w_dly_sig_n[183] tdc0.w_dly_sig[184] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6843 a_5510_9407# a_5342_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6844 VPWR clknet_4_0_0_clk a_5363_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6845 VPWR tdc0.w_dly_sig[171] tdc0.w_dly_sig_n[172] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6846 a_6357_13103# a_5823_13109# a_6262_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6847 VGND tdc0.w_dly_sig[176] tdc0.w_dly_sig_n[176] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6848 tdc0.w_dly_sig_n[115] tdc0.w_dly_sig[115] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6849 VGND tdc0.w_dly_sig[84] tdc0.w_dly_sig_n[84] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6850 VPWR clknet_0_clk a_26882_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6851 VGND a_9339_17429# a_9297_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6852 tdc0.w_dly_sig_n[189] tdc0.w_dly_sig[188] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6853 tdc0.w_dly_sig_n[92] tdc0.w_dly_sig[91] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6854 a_22971_957# a_22107_591# a_22714_703# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6855 a_11816_1513# a_11417_1141# a_11690_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6856 VPWR tdc0.o_result[188] a_19928_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X6857 a_26173_9661# a_25835_9447# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6858 a_17305_17999# a_17139_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6859 VGND tdc0.w_dly_sig[2] tdc0.w_dly_sig_n[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6860 VPWR a_27043_3829# a_27050_4129# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6861 VPWR tdc0.w_dly_sig[102] tdc0.w_dly_sig_n[102] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6862 VGND a_2547_11837# a_2715_11739# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6863 VGND tdc0.w_dly_sig[78] tdc0.w_dly_sig_n[78] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6864 VGND tdc0.w_dly_sig[4] tdc0.w_dly_sig_n[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6865 a_24823_4007# a_24919_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6866 VPWR tdc0.w_dly_sig[148] tdc0.w_dly_sig_n[149] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6867 VGND a_28078_2741# a_28007_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6868 tdc0.o_result[82] a_10903_13915# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6869 a_25375_12711# a_25471_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6870 tdc0.w_dly_sig_n[119] tdc0.w_dly_sig[119] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6871 VPWR tdc0.w_dly_sig_n[182] tdc0.w_dly_sig[184] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6872 VGND tdc0.w_dly_sig_n[74] tdc0.w_dly_sig[76] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6874 tdc0.w_dly_sig_n[15] tdc0.w_dly_sig[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6875 tdc0.w_dly_sig_n[8] tdc0.w_dly_sig[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6876 tdc0.w_dly_sig[83] tdc0.w_dly_sig_n[82] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6877 VGND tdc0.w_dly_sig[80] tdc0.w_dly_sig_n[81] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6878 a_17026_2223# a_16587_2229# a_16941_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6879 a_19579_5719# _011_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X6880 tdc0.w_dly_sig_n[45] tdc0.w_dly_sig[45] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6881 VGND tdc0.w_dly_sig_n[192] tdc0.w_dly_sig[193] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6883 VPWR tdc0.o_result[143] a_14931_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6884 a_20756_5193# _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X6886 VPWR tdc0.w_dly_sig[181] tdc0.w_dly_sig_n[182] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6887 a_15012_9071# tdc0.o_result[91] a_14437_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X6888 a_24283_18761# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6889 VPWR tdc0.w_dly_sig[183] a_26125_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6890 VGND tdc0.w_dly_sig[53] tdc0.w_dly_sig_n[54] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6891 VGND tdc0.w_dly_sig_n[37] tdc0.w_dly_sig[38] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6892 VGND tdc0.w_dly_sig_n[177] tdc0.w_dly_sig[179] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6893 VPWR tdc0.o_result[108] a_5261_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X6894 VPWR a_23075_4007# _052_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6895 a_13722_12559# tdc0.o_result[127] a_13641_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X6896 a_24469_12015# _170_ a_24197_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6897 VGND net26 a_27505_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6898 a_5491_15101# a_4627_14735# a_5234_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6899 tdc0.w_dly_sig[3] tdc0.w_dly_sig_n[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6900 VPWR a_14897_9813# _084_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X6901 VPWR tdc0.w_dly_sig_n[74] tdc0.w_dly_sig[75] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6902 VPWR tdc0.w_dly_sig_n[33] tdc0.w_dly_sig[34] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6903 VGND clknet_4_10_0_clk a_29559_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6904 clknet_4_2_0_clk a_11260_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6905 a_1570_5487# a_1131_5493# a_1485_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6906 a_3686_5487# a_3247_5493# a_3601_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6907 VGND a_26583_11445# a_26590_11745# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6908 _166_ a_12539_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X6910 a_17969_12559# _055_ a_17559_12711# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X6911 tdc0.o_result[142] a_11639_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6912 VPWR a_20945_13675# _055_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X6913 VGND clk a_16210_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6914 VPWR a_20379_15253# a_20295_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6915 VPWR tdc0.w_dly_sig[187] tdc0.w_dly_sig_n[188] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6916 a_11414_6575# a_11141_6581# a_11329_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6917 a_8565_8207# a_8399_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6918 a_17323_7663# net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6919 a_5161_15101# a_4627_14735# a_5066_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6920 VPWR clknet_0_clk a_6476_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6921 VGND a_24005_8725# _189_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X6922 tdc0.w_dly_sig[132] tdc0.w_dly_sig_n[130] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6923 _141_ a_13354_13423# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X6924 a_12778_5461# a_12610_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6926 a_22645_10383# tdc0.w_dly_sig[36] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6927 tdc0.w_dly_sig_n[11] tdc0.w_dly_sig[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6928 a_18823_6059# _030_ a_18737_6059# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X6929 VGND a_17467_10357# _034_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X6930 VGND a_29067_16585# a_29074_16489# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6931 a_24309_15279# _017_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X6932 a_13698_2197# a_13530_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6933 a_7442_2879# a_7274_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6935 VGND a_19487_6183# tdc0.o_result[25] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6936 VPWR clknet_4_0_0_clk a_3523_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6937 tdc0.w_dly_sig[184] tdc0.w_dly_sig_n[183] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6938 VPWR tdc0.w_dly_sig_n[145] tdc0.w_dly_sig[147] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6939 a_6687_5487# a_5989_5493# a_6430_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6940 VPWR a_4371_10901# a_4287_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6941 a_19202_4399# _202_ a_18888_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X6942 a_11785_2229# a_11619_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6944 VPWR a_12254_13103# clknet_4_6_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6945 tdc0.w_dly_sig_n[179] tdc0.w_dly_sig[178] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6946 a_7074_15253# a_6906_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6947 a_12426_11837# a_12153_11471# a_12341_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6948 tdc0.w_dly_sig[27] tdc0.w_dly_sig_n[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6949 tdc0.w_dly_sig_n[162] tdc0.w_dly_sig[161] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6950 a_26309_4943# a_25755_4917# a_25962_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6951 VPWR clknet_4_8_0_clk a_20175_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6953 VPWR tdc0.w_dly_sig_n[125] tdc0.w_dly_sig[126] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6954 a_25891_12559# a_25762_12833# a_25471_12533# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6955 a_15002_2223# a_14729_2229# a_14917_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6956 VPWR tdc0.w_dly_sig_n[8] tdc0.w_dly_sig[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6957 VPWR a_17383_5095# _040_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X6958 VGND tdc0.w_dly_sig[58] tdc0.w_dly_sig_n[58] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6959 tdc0.w_dly_sig_n[110] tdc0.w_dly_sig[110] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6961 tdc0.w_dly_sig[153] tdc0.w_dly_sig_n[151] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6962 VPWR _072_ a_18980_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X6963 VGND tdc0.w_dly_sig[101] tdc0.w_dly_sig_n[102] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6964 a_17409_8457# _105_ a_17313_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6965 tdc0.w_dly_sig[50] tdc0.w_dly_sig_n[48] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6967 VPWR a_7166_14165# a_7093_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6968 VGND clknet_4_2_0_clk a_9595_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6969 tdc0.o_result[91] a_14675_18517# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6970 VGND a_24186_16341# a_24144_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6972 VGND tdc0.w_dly_sig[16] tdc0.w_dly_sig_n[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6973 VPWR a_7331_15279# a_7499_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6974 _058_ a_18703_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6975 a_7005_10383# tdc0.w_dly_sig[129] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6976 VGND a_26939_12247# tdc0.o_result[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6977 a_4732_15657# a_4333_15285# a_4606_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6978 VGND a_1738_7231# a_1696_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6979 a_19885_14191# tdc0.w_dly_sig[69] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6980 VPWR tdc0.o_result[159] a_11527_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6981 a_11693_15285# a_11527_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6982 a_12759_9839# a_11895_9845# a_12502_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
R17 tt_um_hpretl_tt06_tdc_v1_16.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6983 a_3685_15657# a_2695_15285# a_3559_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6984 VGND a_16991_957# a_17159_859# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6985 VGND _110_ a_17415_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6987 VPWR tdc0.w_dly_sig[77] tdc0.w_dly_sig_n[78] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6988 VPWR tdc0.w_dly_sig_n[152] tdc0.w_dly_sig[153] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6989 a_16680_13103# tdc0.o_result[104] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X6990 tdc0.w_dly_sig[141] tdc0.w_dly_sig_n[139] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6991 VPWR a_29607_11159# tdc0.o_result[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6992 a_14287_3855# _007_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6993 _069_ a_19931_4737# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X6994 clknet_4_9_0_clk a_22852_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6995 a_10589_8207# a_10423_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6998 a_22457_10383# a_22291_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6999 _141_ a_13354_13423# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X7001 VGND tdc0.w_dly_sig_n[120] tdc0.w_dly_sig[122] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7002 tdc0.w_dly_sig[191] tdc0.w_dly_sig_n[189] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7005 a_29895_4617# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7006 tdc0.w_dly_sig_n[106] tdc0.w_dly_sig[105] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7007 a_17152_2601# a_16753_2229# a_17026_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7008 VPWR tdc0.o_result[161] a_14195_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7009 a_22303_2601# a_22167_2441# a_21883_2455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7010 VPWR tdc0.o_result[168] a_16311_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7011 tdc0.w_dly_sig[154] tdc0.w_dly_sig_n[152] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7012 VPWR a_25962_15797# a_25891_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X7013 a_22833_12015# _004_ a_22917_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7014 a_5823_10927# _023_ a_6001_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X7015 _130_ a_15115_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X7016 VPWR a_18751_5095# _142_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X7017 tdc0.w_dly_sig[170] tdc0.w_dly_sig_n[169] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7018 tdc0.w_dly_sig[143] tdc0.w_dly_sig_n[141] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7019 uo_out[7] a_20697_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7020 tdc0.w_dly_sig_n[172] tdc0.w_dly_sig[171] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7021 VPWR _065_ a_13552_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X7022 a_17773_14985# tdc0.o_result[125] a_17691_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7023 VPWR tdc0.w_dly_sig[125] tdc0.w_dly_sig_n[125] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7024 VPWR a_5307_6397# a_5475_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7025 a_24653_9545# tdc0.o_result[1] a_24843_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X7026 VPWR tdc0.w_dly_sig[24] tdc0.w_dly_sig_n[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7028 VPWR tdc0.o_result[166] a_12815_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7029 tdc0.w_dly_sig[94] tdc0.w_dly_sig_n[93] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7030 a_27503_5705# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7031 a_12115_1135# a_11417_1141# a_11858_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7033 VGND tdc0.w_dly_sig[60] a_17477_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7034 clknet_4_6_0_clk a_12254_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7036 tdc0.w_dly_sig[181] tdc0.w_dly_sig_n[179] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7037 a_3091_6575# a_2309_6581# a_3007_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7038 a_4333_7119# a_4167_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7039 VPWR a_5234_14847# a_5161_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7041 tdc0.o_result[28] a_22311_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7042 a_3812_5865# a_3413_5493# a_3686_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7043 a_1696_5865# a_1297_5493# a_1570_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7044 tdc0.w_dly_sig[26] tdc0.w_dly_sig_n[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7045 tdc0.w_dly_sig[164] tdc0.w_dly_sig_n[162] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7046 VGND a_30343_7284# net26 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7047 a_6817_10383# a_6651_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7048 VGND tdc0.w_dly_sig_n[173] tdc0.w_dly_sig[175] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7049 a_14591_18543# a_13809_18549# a_14507_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7050 tdc0.w_dly_sig_n[57] tdc0.w_dly_sig[56] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7051 a_8837_11247# tdc0.o_result[79] a_8491_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7052 VGND _051_ a_11681_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7053 VGND tdc0.w_dly_sig[120] tdc0.w_dly_sig_n[120] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7054 a_19727_7119# a_19598_7393# a_19307_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7055 VPWR tdc0.w_dly_sig_n[46] tdc0.w_dly_sig[47] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7056 a_19395_6807# tdc0.o_result[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7057 VPWR a_5291_8725# a_5207_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7059 tdc0.w_dly_sig[152] tdc0.w_dly_sig_n[150] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7060 a_26138_16189# a_25891_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7062 a_14313_10383# _054_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X7064 a_22461_15823# tdc0.w_dly_sig[63] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7065 VGND a_20039_13799# _118_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X7066 a_16679_10383# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7067 VGND net5 a_16355_7969# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7069 _025_ a_14011_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X7070 VPWR a_11490_9407# a_11417_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7071 tdc0.w_dly_sig[103] tdc0.w_dly_sig_n[101] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7072 VGND a_12778_5461# a_12736_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7073 tdc0.w_dly_sig[20] tdc0.w_dly_sig_n[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7074 VPWR clknet_4_7_0_clk a_9687_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7075 VGND tdc0.w_dly_sig_n[99] tdc0.w_dly_sig[100] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7076 a_4057_4399# a_3523_4405# a_3962_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7077 a_16393_3677# tdc0.o_result[168] a_16311_3424# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7078 a_14277_3677# tdc0.o_result[161] a_14195_3424# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7079 a_26966_7485# a_26719_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7080 a_14729_17999# a_14563_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7081 VGND a_26514_6575# clknet_4_11_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X7082 a_23009_8751# a_22475_8757# a_22914_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7083 tdc0.w_dly_sig_n[81] tdc0.w_dly_sig[81] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7084 VPWR tdc0.w_dly_sig_n[121] tdc0.w_dly_sig[122] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7085 a_16025_10633# _020_ a_16109_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7086 VPWR tdc0.w_dly_sig[151] tdc0.w_dly_sig_n[152] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7087 VPWR a_17691_7119# _010_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7088 VGND tdc0.w_dly_sig_n[38] tdc0.w_dly_sig[40] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7089 tdc0.w_dly_sig[121] tdc0.w_dly_sig_n[120] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7090 VPWR clknet_4_13_0_clk a_19531_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7091 clknet_4_14_0_clk a_26882_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7092 VGND tdc0.w_dly_sig_n[131] tdc0.w_dly_sig[133] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7093 a_22687_17277# a_21905_16911# a_22603_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7094 a_14193_13423# _039_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X7095 a_10034_4221# a_9595_3855# a_9949_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7096 VPWR a_9263_16189# a_9431_16091# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
R18 VGND uio_oe[3] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7097 a_4521_7119# tdc0.w_dly_sig[134] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
R19 VGND uio_oe[7] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7099 a_21399_13441# _001_ a_21313_13441# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X7101 VPWR clknet_4_8_0_clk a_20359_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7102 VPWR tdc0.w_dly_sig[111] tdc0.w_dly_sig_n[112] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7103 VGND clknet_4_7_0_clk a_9963_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7104 VGND a_24731_11623# tdc0.o_result[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7105 VPWR clknet_4_2_0_clk a_9595_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7106 a_4521_15279# tdc0.w_dly_sig[103] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7108 tdc0.w_dly_sig[2] tdc0.w_dly_sig_n[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7109 a_24113_16367# a_23579_16373# a_24018_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7110 a_4613_12015# tdc0.w_dly_sig[120] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7112 VPWR tdc0.w_dly_sig[117] tdc0.w_dly_sig_n[117] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7113 a_17578_18365# a_17305_17999# a_17493_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7114 VGND tdc0.w_dly_sig[36] tdc0.w_dly_sig_n[36] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7115 a_8638_3285# a_8470_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7116 a_22001_4399# tdc0.w_dly_sig[32] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7117 _187_ a_23855_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7118 tdc0.w_dly_sig[131] tdc0.w_dly_sig_n[130] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7119 a_19881_15279# a_19347_15285# a_19786_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7121 a_22530_15253# a_22362_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7122 VPWR tdc0.w_dly_sig_n[89] tdc0.w_dly_sig[91] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7123 VPWR a_4111_5487# a_4279_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7124 a_5989_10927# tdc0.o_result[100] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7125 a_15420_8457# _014_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7126 a_3225_8041# a_2235_7669# a_3099_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7127 tdc0.w_dly_sig[152] tdc0.w_dly_sig_n[151] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7129 tdc0.w_dly_sig[76] tdc0.w_dly_sig_n[75] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7130 VPWR tdc0.w_dly_sig[177] a_19685_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7131 a_26351_9295# a_26215_9269# a_25931_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7132 VGND tdc0.w_dly_sig_n[0] tdc0.w_dly_sig[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7133 VGND tdc0.w_dly_sig_n[10] tdc0.w_dly_sig[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7134 VPWR _065_ a_13552_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X7135 tdc0.w_dly_sig_n[184] tdc0.w_dly_sig[183] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7136 VPWR clknet_4_0_0_clk a_6559_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7137 tdc0.w_dly_sig_n[25] tdc0.w_dly_sig[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7138 VGND a_10570_18111# a_10528_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7139 VGND clknet_4_6_0_clk a_9871_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7140 tdc0.w_dly_sig_n[24] tdc0.w_dly_sig[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7142 tdc0.w_dly_sig[166] tdc0.w_dly_sig_n[164] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7143 a_25799_14735# a_25663_14709# a_25379_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7144 tdc0.w_dly_sig[176] tdc0.w_dly_sig_n[174] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7145 a_22362_15279# a_22089_15285# a_22277_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7146 a_12115_1135# a_11251_1141# a_11858_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7147 a_7458_10927# a_7019_10933# a_7373_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7149 a_15483_10383# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7150 a_22227_5487# a_21445_5493# a_22143_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7151 a_22971_13103# a_22107_13109# a_22714_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7152 VGND tdc0.w_dly_sig[76] tdc0.w_dly_sig_n[77] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7153 VGND net3 a_15530_6077# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X7154 VGND a_14989_8353# _101_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X7156 a_1849_13647# a_1683_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7157 a_1754_10927# a_1481_10933# a_1669_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7158 a_8197_3317# a_8031_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7160 VPWR tdc0.w_dly_sig_n[190] tdc0.w_dly_sig[192] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7161 VGND clknet_4_13_0_clk a_17139_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7162 tdc0.w_dly_sig[42] tdc0.w_dly_sig_n[41] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7163 a_4866_11989# a_4698_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7164 VPWR _008_ a_18888_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X7165 tdc0.w_dly_sig[41] tdc0.w_dly_sig_n[40] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7166 VGND clknet_4_0_0_clk a_1131_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7167 net4 a_17634_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7169 tdc0.w_dly_sig_n[126] tdc0.w_dly_sig[126] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7170 a_3785_11471# tdc0.w_dly_sig[119] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7171 VGND tdc0.w_dly_sig[4] tdc0.w_dly_sig_n[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7172 a_8481_10633# tdc0.o_result[112] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X7173 a_16109_9545# tdc0.o_result[75] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7174 a_22641_13103# a_22107_13109# a_22546_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7175 a_29939_5865# a_29803_5705# a_29519_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7176 VGND a_6476_6549# clknet_4_0_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7177 a_5069_9295# a_4903_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7178 a_20211_15279# a_19513_15285# a_19954_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7179 a_18751_5095# tdc0.o_result[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7180 VPWR a_19867_6005# a_19874_6305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7181 a_5767_9661# a_4903_9295# a_5510_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7182 a_24915_8359# a_25011_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7183 tdc0.w_dly_sig_n[154] tdc0.w_dly_sig[154] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7184 a_13997_15279# tdc0.w_dly_sig[87] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7185 _022_ a_16547_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7186 tdc0.w_dly_sig[82] tdc0.w_dly_sig_n[81] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7188 a_27135_7881# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7189 VGND a_17451_2223# a_17619_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7192 a_11923_7663# a_11141_7669# a_11839_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7193 VPWR _019_ a_15483_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X7195 a_10911_18365# a_10129_17999# a_10827_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7196 VPWR a_11582_6549# a_11509_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7197 a_2861_15285# a_2695_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7198 a_15112_13647# tdc0.o_result[86] a_14922_13897# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X7199 tdc0.o_result[129] a_9891_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7200 a_21223_2045# a_20359_1679# a_20966_1791# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7201 a_27066_15556# a_26866_15401# a_27215_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7202 tdc0.w_dly_sig_n[83] tdc0.w_dly_sig[83] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7203 VGND _072_ a_6261_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X7204 tdc0.w_dly_sig[177] tdc0.w_dly_sig_n[175] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7205 VGND a_3819_3285# a_3777_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7206 VGND a_10459_4221# a_10627_4123# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7207 VGND tdc0.w_dly_sig[20] a_27137_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7209 VGND a_29331_7284# net23 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7210 a_27307_8207# a_27087_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X7211 tdc0.w_dly_sig_n[141] tdc0.w_dly_sig[141] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7212 tdc0.w_dly_sig[144] tdc0.w_dly_sig_n[143] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7213 tdc0.w_dly_sig_n[79] tdc0.w_dly_sig[78] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7214 VGND tdc0.w_dly_sig_n[12] tdc0.w_dly_sig[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7215 a_10957_1679# a_10791_1679# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7216 VPWR tdc0.o_result[145] a_14379_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7217 a_14208_15657# a_13809_15285# a_14082_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7218 VGND tdc0.w_dly_sig_n[155] tdc0.w_dly_sig[157] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7219 VPWR tdc0.w_dly_sig[91] tdc0.w_dly_sig_n[91] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7220 a_14703_3543# _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X7221 VGND a_30591_3285# a_30549_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7222 VGND a_25375_15975# tdc0.o_result[48] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7223 _071_ a_20543_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X7224 VPWR tdc0.w_dly_sig[112] tdc0.w_dly_sig_n[113] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7225 a_18390_16341# a_18222_16367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7226 a_4111_5487# a_3413_5493# a_3854_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7227 a_17965_4719# _008_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X7228 tdc0.w_dly_sig[64] tdc0.w_dly_sig_n[62] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7229 tdc0.w_dly_sig[146] tdc0.w_dly_sig_n[144] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7230 a_18703_14985# _065_ a_18785_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7231 a_26966_11837# a_26719_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7232 a_22787_15279# a_22089_15285# a_22530_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7233 tdc0.w_dly_sig_n[148] tdc0.w_dly_sig[147] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7234 tdc0.w_dly_sig[147] tdc0.w_dly_sig_n[145] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7235 VPWR a_6550_12559# clknet_4_4_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7236 VGND tdc0.w_dly_sig[119] tdc0.w_dly_sig_n[120] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7237 VGND _134_ a_18703_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7238 a_17535_2223# a_16753_2229# a_17451_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7239 VGND net27 a_27689_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7240 a_22063_17821# a_21843_17833# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X7241 a_10310_12925# a_9871_12559# a_10225_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7243 VGND tdc0.w_dly_sig[128] tdc0.w_dly_sig_n[128] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7244 VGND a_22603_17277# a_22771_17179# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7245 _132_ a_5823_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X7246 a_10160_3855# a_9761_3855# a_10034_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7248 VPWR _037_ a_16837_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7249 VGND a_2731_9839# a_2899_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7250 tdc0.w_dly_sig[23] tdc0.w_dly_sig_n[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7251 VPWR tdc0.w_dly_sig_n[155] tdc0.w_dly_sig[156] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7252 VPWR a_24186_16341# a_24113_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7254 a_3877_4399# tdc0.w_dly_sig[149] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7255 a_3302_15253# a_3134_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7256 a_25375_13647# a_25155_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X7257 a_3597_11471# a_3431_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7258 a_23075_11159# a_23171_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7259 tdc0.w_dly_sig_n[39] tdc0.w_dly_sig[38] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7260 VPWR a_19954_15253# a_19881_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7261 tdc0.w_dly_sig[187] tdc0.w_dly_sig_n[185] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7262 VPWR clknet_4_5_0_clk a_6375_16373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7263 tdc0.w_dly_sig_n[125] tdc0.w_dly_sig[124] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7266 a_17076_12015# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7267 VPWR tdc0.w_dly_sig_n[113] tdc0.w_dly_sig[114] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7268 VPWR a_12927_9813# a_12843_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7269 a_17559_12711# _111_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X7270 a_22395_12559# a_22259_12533# a_21975_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7271 a_20782_2879# a_20614_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7272 VPWR _085_ a_16109_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7273 a_7699_3133# a_6835_2767# a_7442_2879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7274 VPWR a_28595_7284# net27 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7275 VPWR tdc0.w_dly_sig[158] tdc0.w_dly_sig_n[158] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7277 VPWR a_16713_8235# _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X7278 VPWR clknet_4_9_0_clk a_22475_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7279 VGND tdc0.w_dly_sig_n[191] tdc0.w_dly_sig[193] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7280 VGND tdc0.w_dly_sig[72] tdc0.w_dly_sig_n[73] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7281 tdc0.o_result[156] a_6395_3035# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7282 VPWR a_16916_4373# _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7283 tdc0.w_dly_sig[138] tdc0.w_dly_sig_n[136] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7284 tdc0.w_dly_sig[87] tdc0.w_dly_sig_n[85] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7285 VGND a_13149_6549# _165_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X7286 VPWR tdc0.w_dly_sig[30] tdc0.w_dly_sig_n[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7287 tdc0.w_dly_sig_n[76] tdc0.w_dly_sig[76] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R20 uio_oe[1] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7288 VPWR clknet_4_5_0_clk a_8307_17461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7289 a_1485_7119# tdc0.w_dly_sig[114] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7290 a_12977_14735# a_11987_14735# a_12851_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7291 VPWR tdc0.w_dly_sig[79] tdc0.w_dly_sig_n[79] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7292 a_25849_8207# a_25295_8181# a_25502_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7293 VGND a_2750_6549# a_2708_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7294 a_11839_14191# a_10975_14197# a_11582_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7295 VGND tdc0.w_dly_sig_n[114] tdc0.w_dly_sig[116] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7296 VPWR _060_ a_22790_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X7298 a_14821_15823# a_14655_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7299 a_30549_14569# a_29559_14197# a_30423_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7300 VGND a_12594_11583# a_12552_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7301 tdc0.o_result[76] a_15227_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7303 a_28783_16599# a_29067_16585# a_29002_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X7304 tdc0.w_dly_sig[131] tdc0.w_dly_sig_n[129] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7305 VGND tdc0.w_dly_sig[85] tdc0.w_dly_sig_n[86] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7306 a_7350_7231# a_7182_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7307 a_27965_13481# a_27411_13321# a_27618_13380# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7308 tdc0.w_dly_sig[112] tdc0.w_dly_sig_n[111] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7309 a_27250_4676# a_27050_4521# a_27399_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7310 VPWR a_22714_13077# a_22641_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7311 _134_ a_15943_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X7312 tdc0.w_dly_sig_n[142] tdc0.w_dly_sig[142] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7314 tdc0.w_dly_sig[59] tdc0.w_dly_sig_n[57] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7316 a_8565_8207# a_8399_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7317 tdc0.w_dly_sig_n[100] tdc0.w_dly_sig[99] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7318 VGND a_7378_13103# clknet_4_5_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X7320 a_26215_9269# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7321 tdc0.w_dly_sig[94] tdc0.w_dly_sig_n[92] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7322 _046_ a_13722_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X7323 a_13622_16367# a_13183_16373# a_13537_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7324 VGND tdc0.w_dly_sig_n[1] tdc0.w_dly_sig[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7325 a_24398_1412# a_24198_1257# a_24547_1501# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7326 VGND a_12134_15253# a_12092_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7327 VPWR a_15059_10927# a_15227_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7328 a_22090_10927# a_21843_11305# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7329 VGND a_8971_2197# a_8929_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7330 VPWR tdc0.w_dly_sig[22] a_25665_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7331 a_18647_16367# a_17949_16373# a_18390_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7332 _155_ a_13275_7776# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7333 VGND a_21313_13441# _004_ VGND sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X7334 a_20359_11721# _016_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7335 VGND a_20325_5089# _197_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X7336 tdc0.w_dly_sig_n[73] tdc0.w_dly_sig[73] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7339 VPWR tdc0.w_dly_sig[173] tdc0.w_dly_sig_n[173] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7340 _066_ a_18703_14985# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X7341 a_7553_12021# a_7387_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7342 a_8470_3311# a_8031_3317# a_8385_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7343 a_16749_2767# a_15759_2767# a_16623_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7344 a_19069_8207# _072_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X7345 VGND tdc0.w_dly_sig_n[32] tdc0.w_dly_sig[33] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7346 a_27871_2741# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7347 tdc0.o_result[141] a_10259_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7348 a_4111_5487# a_3247_5493# a_3854_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7349 a_7001_14735# a_6835_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7350 a_18383_8983# tdc0.o_result[58] a_18617_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7351 VPWR a_19225_11721# uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7352 VGND a_3727_15253# a_3685_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7353 a_27158_8181# a_26958_8481# a_27307_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7354 VPWR tdc0.w_dly_sig_n[156] tdc0.w_dly_sig[157] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7355 tdc0.o_result[80] a_10995_11739# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7357 VGND tdc0.w_dly_sig[157] tdc0.w_dly_sig_n[158] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7358 VGND tdc0.w_dly_sig[160] tdc0.w_dly_sig_n[161] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7359 a_21567_8207# a_21438_8481# a_21147_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7360 VPWR _002_ a_18703_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X7361 VGND a_16210_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X7362 VPWR tdc0.w_dly_sig[81] tdc0.w_dly_sig_n[82] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7363 a_20609_11721# _063_ a_20881_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7364 VPWR tdc0.w_dly_sig[65] tdc0.w_dly_sig_n[65] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7365 VPWR a_21707_17673# a_21714_17577# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7366 tdc0.w_dly_sig[60] tdc0.w_dly_sig_n[59] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7367 a_19867_11145# clknet_4_13_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7370 a_11414_14191# a_11141_14197# a_11329_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7372 VPWR a_21380_14165# clknet_4_12_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7373 VPWR tdc0.w_dly_sig[158] tdc0.w_dly_sig_n[159] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7374 a_30124_14569# a_29725_14197# a_29998_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7375 a_23138_13897# _147_ a_23058_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X7376 a_26719_11471# a_26583_11445# a_26299_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7377 a_12058_2223# a_11619_2229# a_11973_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7379 VPWR a_15795_12925# a_15963_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7380 a_5261_10927# _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X7381 VGND clknet_4_0_0_clk a_2051_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7382 a_7442_14847# a_7274_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7383 a_29423_5719# a_29519_5719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7384 a_27250_4676# a_27043_4617# a_27426_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7385 tdc0.w_dly_sig_n[30] tdc0.w_dly_sig[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7386 a_10589_8207# a_10423_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7387 VGND clknet_4_6_0_clk a_10975_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7388 tdc0.w_dly_sig[190] tdc0.w_dly_sig_n[188] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7389 a_24363_4007# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X7390 a_24639_13799# a_24735_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7391 a_12254_13103# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7393 VGND tdc0.w_dly_sig_n[17] tdc0.w_dly_sig[18] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7394 a_5161_15823# a_4995_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7395 VGND a_8051_10901# a_8009_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7396 a_24398_1412# a_24191_1353# a_24574_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7397 clknet_4_11_0_clk a_26514_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7398 a_13997_18543# tdc0.w_dly_sig[92] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7399 tdc0.w_dly_sig_n[41] tdc0.w_dly_sig[41] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7400 a_6388_13481# a_5989_13109# a_6262_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7401 a_16356_9071# _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X7402 tdc0.w_dly_sig[188] tdc0.w_dly_sig_n[187] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7403 a_15059_10927# a_14195_10933# a_14802_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7404 a_8837_8041# a_7847_7669# a_8711_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7405 a_13698_2197# a_13530_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7406 tdc0.o_result[170] a_17159_859# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7407 tdc0.w_dly_sig_n[139] tdc0.w_dly_sig[138] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7408 a_24131_9295# _071_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X7409 tdc0.w_dly_sig_n[162] tdc0.w_dly_sig[162] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7410 tdc0.w_dly_sig[88] tdc0.w_dly_sig_n[86] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7411 VPWR tdc0.w_dly_sig_n[87] tdc0.w_dly_sig[88] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7412 a_20051_10057# clknet_4_13_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7413 VPWR tdc0.w_dly_sig[55] a_22261_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7414 VGND a_29090_13380# a_29019_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X7416 a_4977_8573# a_4443_8207# a_4882_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7417 VPWR tdc0.w_dly_sig[176] tdc0.w_dly_sig_n[177] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7419 VGND a_21327_3543# _082_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X7420 VGND clknet_4_9_0_clk a_23027_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7421 VPWR net6 a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7422 VPWR a_12283_1109# a_12199_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7423 VPWR tdc0.o_result[187] a_23303_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7424 a_7515_10749# a_6817_10383# a_7258_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7425 VPWR tdc0.w_dly_sig_n[146] tdc0.w_dly_sig[148] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7426 clknet_4_2_0_clk a_11260_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X7427 tdc0.w_dly_sig_n[78] tdc0.w_dly_sig[78] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7428 VPWR tdc0.w_dly_sig_n[80] tdc0.w_dly_sig[81] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7429 VPWR a_25375_12711# tdc0.o_result[38] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7430 a_7507_3311# a_6725_3317# a_7423_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7431 a_16753_15101# a_16219_14735# a_16658_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7432 a_21914_11204# a_21707_11145# a_22090_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7433 a_27597_4777# a_27043_4617# a_27250_4676# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7434 VPWR a_30515_6397# a_30683_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7435 VGND tdc0.w_dly_sig[169] tdc0.w_dly_sig_n[169] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7436 VPWR tdc0.w_dly_sig[18] tdc0.w_dly_sig_n[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7437 VPWR tdc0.w_dly_sig[90] tdc0.w_dly_sig_n[90] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7438 a_22089_15285# a_21923_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7439 a_13257_2229# a_13091_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7440 VGND tdc0.w_dly_sig_n[102] tdc0.w_dly_sig[104] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7441 VPWR a_2547_12925# a_2715_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7442 tdc0.w_dly_sig_n[101] tdc0.w_dly_sig[100] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7443 VPWR _022_ a_15101_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7444 a_17814_8751# _033_ a_17565_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7446 tdc0.w_dly_sig_n[30] tdc0.w_dly_sig[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7447 a_3394_14165# a_3226_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7448 tdc0.w_dly_sig_n[186] tdc0.w_dly_sig[185] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7449 a_24745_1513# a_24191_1353# a_24398_1412# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7450 a_17503_7663# a_17323_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7451 a_20499_13799# tdc0.o_result[55] a_20733_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7454 VGND a_17691_7119# _010_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X7455 tdc0.w_dly_sig[38] tdc0.w_dly_sig_n[37] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7456 VPWR a_5935_9563# a_5851_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7457 VGND tdc0.w_dly_sig_n[173] tdc0.w_dly_sig[174] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7458 a_13552_6281# tdc0.o_result[136] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X7459 a_17010_17429# a_16842_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7461 a_8596_3689# a_8197_3317# a_8470_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7462 a_26719_7119# a_26590_7393# a_26299_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7463 VGND a_10506_7119# clknet_4_3_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7464 tdc0.w_dly_sig_n[135] tdc0.w_dly_sig[134] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7465 VPWR a_21391_1947# a_21307_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7466 tdc0.w_dly_sig_n[124] tdc0.w_dly_sig[123] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7468 a_17967_9839# _112_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7469 tdc0.w_dly_sig_n[42] tdc0.w_dly_sig[42] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7470 tdc0.w_dly_sig[99] tdc0.w_dly_sig_n[98] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7471 a_27505_8207# a_26951_8181# a_27158_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7472 a_8933_14013# a_8399_13647# a_8838_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7473 a_27871_2741# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7474 a_7001_14735# a_6835_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7475 VPWR tdc0.w_dly_sig[136] tdc0.w_dly_sig_n[136] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7476 VPWR tdc0.w_dly_sig_n[100] tdc0.w_dly_sig[101] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7478 a_23075_4007# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X7479 VGND _144_ a_18046_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X7480 VGND tdc0.w_dly_sig_n[61] tdc0.w_dly_sig[62] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7481 VPWR a_23139_16091# a_23055_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7482 VGND a_21886_5461# a_21844_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7483 a_23385_3677# tdc0.o_result[187] a_23303_3424# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7485 VGND a_2290_13759# a_2248_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7486 a_9025_8757# a_8859_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7487 a_14385_10383# _034_ a_14313_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7488 VGND clknet_4_8_0_clk a_20359_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7490 a_27426_4399# a_27179_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7491 a_24731_7271# a_24827_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7492 VPWR net1 tdc0.w_dly_sig_n[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7493 _034_ a_17467_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7494 VPWR tdc0.w_dly_sig[103] tdc0.w_dly_sig_n[104] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7495 VPWR _076_ a_12999_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X7497 VGND _096_ a_17565_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X7498 a_12184_2601# a_11785_2229# a_12058_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7499 VPWR a_25428_7637# clknet_4_10_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7501 a_24574_1135# a_24327_1513# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7502 VPWR tdc0.w_dly_sig[45] tdc0.w_dly_sig_n[46] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7503 VPWR tdc0.w_dly_sig_n[140] tdc0.w_dly_sig[141] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7504 _011_ net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7505 VGND tdc0.w_dly_sig[31] tdc0.w_dly_sig_n[31] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7506 VPWR clknet_4_7_0_clk a_13643_18549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7507 a_10961_4943# tdc0.w_dly_sig[143] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7508 a_17703_6895# net6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7509 a_22637_4777# a_21647_4405# a_22511_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7510 VGND a_18130_591# a_18236_591# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X7511 VGND _084_ a_14563_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X7512 VPWR a_12559_15253# a_12475_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7513 VPWR tdc0.w_dly_sig[172] tdc0.w_dly_sig_n[173] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7514 _064_ _001_ a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7515 uo_out[1] a_24653_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R21 uio_out[0] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7516 a_18489_9839# _064_ a_17967_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7518 tdc0.w_dly_sig[9] tdc0.w_dly_sig_n[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7519 a_20204_9545# _014_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7520 a_27526_10116# a_27319_10057# a_27702_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7521 a_10126_17277# a_9687_16911# a_10041_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7522 a_19544_18921# a_19145_18549# a_19418_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7523 VPWR tdc0.w_dly_sig[70] tdc0.w_dly_sig_n[70] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7524 tdc0.w_dly_sig[17] tdc0.w_dly_sig_n[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7525 VPWR a_14507_18543# a_14675_18517# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7526 tdc0.w_dly_sig_n[102] tdc0.w_dly_sig[101] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7527 a_4425_8757# a_4259_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7528 VPWR a_6687_4399# a_6855_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7530 tdc0.w_dly_sig[39] tdc0.w_dly_sig_n[38] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7531 a_27491_8029# a_27271_8041# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X7532 a_13722_8207# _033_ a_13968_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X7533 tdc0.w_dly_sig_n[63] tdc0.w_dly_sig[63] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7534 VPWR net4 a_17953_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X7535 VGND net4 _009_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7536 VGND a_14507_18543# a_14675_18517# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7537 VPWR tdc0.w_dly_sig[37] tdc0.w_dly_sig_n[37] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7538 VPWR a_10459_4221# a_10627_4123# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7539 tdc0.o_result[58] a_17435_17429# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7540 VGND _094_ a_17415_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7541 VGND tdc0.w_dly_sig[90] tdc0.w_dly_sig_n[91] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7542 VPWR a_7867_3035# a_7783_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7543 a_2631_14013# a_1849_13647# a_2547_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7544 VGND a_14255_6835# _035_ VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X7547 VGND a_5307_8573# a_5475_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7548 tdc0.w_dly_sig_n[155] tdc0.w_dly_sig[154] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7550 VGND _043_ a_12969_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7551 a_13997_17455# tdc0.w_dly_sig[91] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7552 VGND clknet_4_7_0_clk a_11527_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7553 a_9666_4399# a_9393_4405# a_9581_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7554 a_8491_10927# _027_ a_8573_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7555 a_11781_1679# a_10791_1679# a_11655_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7556 VGND tdc0.w_dly_sig_n[164] tdc0.w_dly_sig[165] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7557 VPWR a_11812_13621# clknet_4_7_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7558 VPWR _047_ a_16680_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X7559 VPWR a_16826_14847# a_16753_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7560 tdc0.w_dly_sig_n[6] tdc0.w_dly_sig[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7561 tdc0.w_dly_sig[119] tdc0.w_dly_sig_n[118] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7563 a_19415_11721# tdc0.o_result[4] a_19225_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X7564 VGND a_6476_7637# clknet_4_1_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7566 tdc0.w_dly_sig_n[74] tdc0.w_dly_sig[74] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7567 a_6262_5487# a_5823_5493# a_6177_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7568 tdc0.w_dly_sig_n[136] tdc0.w_dly_sig[136] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7569 a_11509_7663# a_10975_7669# a_11414_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7572 VPWR a_15333_4737# _039_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X7573 a_29817_6031# a_29651_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7574 tdc0.w_dly_sig_n[19] tdc0.w_dly_sig[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7575 a_10735_14013# a_10037_13647# a_10478_13759# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7576 _007_ a_14983_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7578 VGND _033_ a_14182_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X7579 a_20223_6031# a_20003_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X7581 a_2497_6575# tdc0.w_dly_sig[151] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7582 a_22917_12015# tdc0.o_result[37] a_22833_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7583 VGND clknet_4_0_0_clk a_8031_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7584 VGND tdc0.w_dly_sig[133] tdc0.w_dly_sig_n[134] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7585 tdc0.w_dly_sig_n[176] tdc0.w_dly_sig[176] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7587 clknet_4_6_0_clk a_12254_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7588 a_26125_1679# a_25571_1653# a_25778_1653# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7589 VGND a_20697_12809# uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7590 _028_ a_8399_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X7591 VPWR tdc0.w_dly_sig[23] tdc0.w_dly_sig_n[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7592 clknet_0_clk a_16210_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7593 a_13955_2223# a_13257_2229# a_13698_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7594 VGND a_25375_5095# tdc0.o_result[20] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7595 a_21327_17687# a_21423_17687# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7596 a_24469_12015# _064_ a_23947_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7597 a_13897_11471# tdc0.o_result[106] a_13551_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7598 VPWR tdc0.w_dly_sig[107] tdc0.w_dly_sig_n[108] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7599 VPWR a_2547_11837# a_2715_11739# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7600 a_26790_11445# a_26590_11745# a_26939_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7601 _011_ a_16495_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7602 VPWR a_2163_5461# a_2079_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7603 tdc0.w_dly_sig_n[32] tdc0.w_dly_sig[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7604 a_15128_17999# a_14729_17999# a_15002_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7605 VGND tdc0.w_dly_sig_n[66] tdc0.w_dly_sig[67] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7606 a_5993_3855# tdc0.w_dly_sig[158] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7607 _060_ a_16127_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X7608 VGND tdc0.w_dly_sig_n[122] tdc0.w_dly_sig[124] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7609 a_27158_8181# a_26951_8181# a_27334_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7612 a_18751_5095# _011_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X7613 a_14507_18543# a_13643_18549# a_14250_18517# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7614 tdc0.w_dly_sig[5] tdc0.w_dly_sig_n[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7615 tdc0.o_result[168] a_15595_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7617 tdc0.w_dly_sig[70] tdc0.w_dly_sig_n[68] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7618 tdc0.w_dly_sig_n[40] tdc0.w_dly_sig[39] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7619 a_7373_10927# tdc0.w_dly_sig[80] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7620 tdc0.w_dly_sig_n[120] tdc0.w_dly_sig[120] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7621 tdc0.o_result[173] a_16791_3035# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7622 VGND clknet_4_1_0_clk a_3707_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7623 VPWR tdc0.w_dly_sig[101] tdc0.w_dly_sig_n[101] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7624 tdc0.o_result[109] a_1979_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7625 a_22852_7093# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7628 tdc0.o_result[94] a_10995_18267# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7629 a_27702_9839# a_27455_10217# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7630 tdc0.w_dly_sig_n[96] tdc0.w_dly_sig[96] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7631 a_24843_9545# tdc0.o_result[1] a_24653_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X7632 a_14177_18543# a_13643_18549# a_14082_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7634 VPWR a_5050_6143# a_4977_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7635 a_18489_9839# tdc0.o_result[3] a_17967_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X7636 a_26790_7093# a_26590_7393# a_26939_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7637 tdc0.w_dly_sig[46] tdc0.w_dly_sig_n[44] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7639 VGND _051_ a_11865_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7641 VGND a_30591_14165# a_30549_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7642 tdc0.o_result[148] a_4555_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7643 VPWR a_6476_6549# clknet_4_0_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7644 a_29067_16585# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7645 VGND _035_ a_16833_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7646 a_18141_11721# _149_ a_18059_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X7647 _172_ a_5639_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X7648 _059_ a_16495_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7649 VPWR a_27319_12233# a_27326_12137# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7650 a_22730_10749# a_22291_10383# a_22645_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7651 tdc0.w_dly_sig[122] tdc0.w_dly_sig_n[121] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7652 a_16109_10633# tdc0.o_result[92] a_16025_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7653 a_6771_4399# a_5989_4405# a_6687_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7654 VGND net6 _013_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7655 VGND tdc0.w_dly_sig_n[66] tdc0.w_dly_sig[68] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7656 tdc0.w_dly_sig_n[119] tdc0.w_dly_sig[119] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7657 tdc0.o_result[122] a_6855_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7658 a_7741_12015# tdc0.w_dly_sig[128] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7659 tdc0.w_dly_sig[79] tdc0.w_dly_sig_n[77] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7660 tdc0.o_result[75] a_12927_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7661 VPWR clknet_4_7_0_clk a_13643_17461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7662 a_12935_16189# a_12153_15823# a_12851_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7663 VGND clknet_4_0_0_clk a_947_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7664 VGND tdc0.w_dly_sig_n[49] tdc0.w_dly_sig[50] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7665 VPWR a_2731_9839# a_2899_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7666 tdc0.o_result[139] a_12007_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7667 VPWR tdc0.w_dly_sig[128] tdc0.w_dly_sig_n[128] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7668 tdc0.w_dly_sig[65] tdc0.w_dly_sig_n[64] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7669 VGND tdc0.w_dly_sig_n[162] tdc0.w_dly_sig[163] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7670 VPWR tdc0.w_dly_sig_n[26] tdc0.w_dly_sig[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7671 a_22273_15823# a_22107_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7672 a_15921_12559# a_14931_12559# a_15795_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7673 VGND a_12483_2223# a_12651_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7674 VGND _026_ a_11589_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7675 tdc0.w_dly_sig_n[182] tdc0.w_dly_sig[181] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7678 a_3505_10933# a_3339_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7679 _000_ net6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7681 a_7649_4399# tdc0.w_dly_sig[144] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7682 a_14185_4943# tdc0.o_result[162] a_14103_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7683 clknet_4_3_0_clk a_10506_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7685 tdc0.w_dly_sig_n[167] tdc0.w_dly_sig[167] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7686 tdc0.w_dly_sig_n[170] tdc0.w_dly_sig[170] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7687 VPWR tdc0.w_dly_sig_n[22] tdc0.w_dly_sig[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7688 a_18479_6895# _001_ _064_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7689 VGND _017_ a_24385_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X7690 tdc0.o_result[144] a_13203_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7691 VPWR tdc0.w_dly_sig[99] tdc0.w_dly_sig_n[99] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7692 VPWR tdc0.w_dly_sig_n[20] tdc0.w_dly_sig[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7693 VPWR tdc0.w_dly_sig[19] tdc0.w_dly_sig_n[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7694 _036_ a_16679_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7695 VGND a_5031_15279# a_5199_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7696 _017_ a_19289_13441# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X7698 a_12618_7983# _123_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X7699 VPWR tdc0.w_dly_sig[84] tdc0.w_dly_sig_n[85] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7700 VPWR tdc0.w_dly_sig[108] tdc0.w_dly_sig_n[108] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7701 VGND tdc0.o_result[67] a_16684_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X7702 a_26111_15823# a_25891_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X7703 a_29987_11445# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7704 VPWR _030_ a_19855_8359# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X7705 a_22615_4007# tdc0.o_result[189] a_22849_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7706 a_6388_5865# a_5989_5493# a_6262_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7707 a_12999_8867# _161_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7708 tdc0.w_dly_sig_n[166] tdc0.w_dly_sig[165] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7709 tdc0.w_dly_sig_n[31] tdc0.w_dly_sig[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7710 VPWR a_25410_13103# clknet_4_15_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7711 tdc0.w_dly_sig[135] tdc0.w_dly_sig_n[133] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7712 a_8753_9295# tdc0.w_dly_sig[127] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7713 VGND a_16791_3035# a_16749_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7714 a_12567_2223# a_11785_2229# a_12483_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7715 a_20074_6005# a_19874_6305# a_20223_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7716 a_29423_6196# tdc0.w_dly_sig[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7717 VGND _197_ a_19255_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7719 VGND tdc0.w_dly_sig_n[166] tdc0.w_dly_sig[168] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7720 a_27334_8573# a_27087_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7721 a_22672_13481# a_22273_13109# a_22546_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7722 a_24419_2767# a_24290_3041# a_23999_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7723 VPWR tdc0.w_dly_sig_n[147] tdc0.w_dly_sig[148] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7724 VGND _085_ a_16381_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X7725 tdc0.w_dly_sig_n[84] tdc0.w_dly_sig[83] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7726 VPWR tdc0.o_result[129] a_11159_8864# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7727 VGND _019_ a_15637_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7728 VPWR a_12999_8867# _170_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7729 a_20881_11721# tdc0.o_result[0] a_20359_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X7730 _199_ a_12999_3424# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7731 a_11413_8207# a_10423_8207# a_11287_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7732 tdc0.w_dly_sig_n[106] tdc0.w_dly_sig[106] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7733 a_7189_14735# tdc0.w_dly_sig[126] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7734 a_8753_15823# tdc0.w_dly_sig[100] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7735 VGND tdc0.w_dly_sig[26] tdc0.w_dly_sig_n[27] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7737 VGND a_17323_6575# _030_ VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7738 a_19395_6807# tdc0.o_result[16] a_19629_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7739 a_22813_12559# a_22259_12533# a_22466_12533# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7740 a_14917_2223# tdc0.w_dly_sig[169] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7741 a_11398_1791# a_11230_2045# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7742 a_29913_8751# tdc0.w_dly_sig[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7743 VPWR clknet_4_1_0_clk a_4903_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7744 tdc0.w_dly_sig_n[185] tdc0.w_dly_sig[185] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7745 a_14922_13647# tdc0.o_result[94] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X7746 VGND _198_ a_13722_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X7747 VGND tdc0.w_dly_sig[179] tdc0.w_dly_sig_n[179] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7748 VPWR clknet_4_3_0_clk a_10975_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
R22 VGND uio_oe[6] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7749 VGND tdc0.w_dly_sig[50] tdc0.w_dly_sig_n[50] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7750 VPWR tdc0.o_result[183] a_23027_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X7751 VGND tdc0.w_dly_sig[162] tdc0.w_dly_sig_n[163] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7752 a_26759_3829# a_27050_4129# a_27001_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7753 tdc0.w_dly_sig_n[1] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7755 VGND tdc0.w_dly_sig[167] tdc0.w_dly_sig_n[168] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7756 tdc0.w_dly_sig_n[121] tdc0.w_dly_sig[121] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7757 a_12264_8457# tdc0.o_result[77] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X7759 a_11582_6549# a_11414_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7760 VGND a_11260_5461# clknet_4_2_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7761 a_5989_5493# a_5823_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7762 a_10827_18365# a_9963_17999# a_10570_18111# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7763 VPWR clknet_4_5_0_clk a_2695_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7764 a_7470_6005# a_7263_6005# a_7646_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7765 _035_ a_14255_6835# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X7766 a_8385_16367# tdc0.w_dly_sig[98] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7767 a_29913_14191# tdc0.w_dly_sig[45] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7768 a_7097_7119# tdc0.w_dly_sig[136] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7769 VPWR a_15262_15935# a_15189_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7770 VGND a_20881_11721# uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7771 VPWR tdc0.w_dly_sig[34] tdc0.w_dly_sig_n[34] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7772 VPWR tdc0.w_dly_sig_n[35] tdc0.w_dly_sig[37] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7773 a_27597_4777# a_27050_4521# a_27250_4676# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X7774 a_30090_6397# a_29817_6031# a_30005_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7775 VGND tdc0.w_dly_sig_n[160] tdc0.w_dly_sig[161] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7776 clknet_4_11_0_clk a_26514_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7777 a_15049_4765# _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X7778 tdc0.w_dly_sig_n[66] tdc0.w_dly_sig[65] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7779 a_21787_3543# tdc0.o_result[178] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7781 tdc0.o_result[73] a_11915_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7782 a_5031_15279# a_4167_15285# a_4774_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7783 tdc0.w_dly_sig[37] tdc0.w_dly_sig_n[36] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7784 a_27137_7119# a_26583_7093# a_26790_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7785 tdc0.o_result[115] a_3267_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7786 a_10497_18365# a_9963_17999# a_10402_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7787 tdc0.w_dly_sig[126] tdc0.w_dly_sig_n[124] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7788 a_1754_10927# a_1315_10933# a_1669_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7789 VPWR clknet_4_1_0_clk a_7847_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7790 a_24843_9545# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7791 a_24745_1513# a_24198_1257# a_24398_1412# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X7792 VPWR tdc0.w_dly_sig_n[129] tdc0.w_dly_sig[130] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7793 tdc0.w_dly_sig[172] tdc0.w_dly_sig_n[171] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7794 tdc0.w_dly_sig[44] tdc0.w_dly_sig_n[42] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7795 tdc0.w_dly_sig[175] tdc0.w_dly_sig_n[173] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7796 VPWR tdc0.w_dly_sig[61] tdc0.w_dly_sig_n[61] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7797 VPWR tdc0.w_dly_sig_n[152] tdc0.w_dly_sig[154] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7798 VGND a_13790_16341# a_13748_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7799 tdc0.w_dly_sig[173] tdc0.w_dly_sig_n[171] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7800 a_10217_4777# a_9227_4405# a_10091_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7801 a_21633_5487# tdc0.w_dly_sig[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7802 a_16739_7895# net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X7803 a_12149_18921# a_11159_18549# a_12023_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7804 VPWR tdc0.w_dly_sig_n[137] tdc0.w_dly_sig[139] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7805 a_3007_6575# a_2143_6581# a_2750_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7806 tdc0.w_dly_sig_n[62] tdc0.w_dly_sig[61] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7807 a_15879_12925# a_15097_12559# a_15795_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7808 a_22546_16189# a_22107_15823# a_22461_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7809 a_18703_11471# _132_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7810 VGND tdc0.w_dly_sig[70] tdc0.w_dly_sig_n[71] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7811 VPWR tdc0.w_dly_sig[110] tdc0.w_dly_sig_n[110] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7812 a_10570_18111# a_10402_18365# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7813 VPWR tdc0.w_dly_sig[174] tdc0.w_dly_sig_n[174] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7814 tdc0.w_dly_sig_n[128] tdc0.w_dly_sig[128] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7815 a_10317_11471# tdc0.w_dly_sig[81] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7816 a_23155_10749# a_22291_10383# a_22898_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7817 VGND tdc0.w_dly_sig_n[108] tdc0.w_dly_sig[110] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7819 a_23518_9839# _128_ a_23269_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7820 a_16938_16189# a_16691_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7821 VGND a_7423_14191# a_7591_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7822 VPWR _054_ a_12539_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X7824 tdc0.w_dly_sig_n[65] tdc0.w_dly_sig[65] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7826 VPWR tdc0.w_dly_sig_n[64] tdc0.w_dly_sig[66] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7827 VPWR tdc0.w_dly_sig_n[186] tdc0.w_dly_sig[187] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7828 a_15397_3677# _038_ a_15325_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7829 VPWR tdc0.w_dly_sig_n[103] tdc0.w_dly_sig[105] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7830 a_6001_11247# tdc0.o_result[116] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X7831 VGND a_11679_8983# _027_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X7832 VGND _007_ a_15085_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7833 tdc0.w_dly_sig_n[28] tdc0.w_dly_sig[27] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7834 VGND a_23075_11159# tdc0.o_result[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7836 tdc0.w_dly_sig_n[187] tdc0.w_dly_sig[187] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7837 VPWR a_16210_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7838 VPWR a_26479_15511# tdc0.o_result[47] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7839 VGND tdc0.w_dly_sig_n[110] tdc0.w_dly_sig[111] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7840 a_15511_2223# a_14729_2229# a_15427_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7841 a_24242_8457# _107_ a_24162_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X7842 a_17393_17833# a_16403_17461# a_17267_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7843 a_20893_14735# a_20727_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7845 VGND a_19735_859# a_19693_591# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7846 a_29090_12292# a_28890_12137# a_29239_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7847 a_20039_5719# tdc0.o_result[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7848 VPWR tdc0.w_dly_sig[130] tdc0.w_dly_sig_n[130] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7849 VPWR tdc0.o_result[56] a_17076_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X7850 VPWR a_9834_4373# a_9761_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7851 a_23027_5487# _031_ a_23110_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X7852 uo_out[2] a_17937_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7853 VPWR a_25410_3829# a_25339_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X7854 a_9006_8319# a_8838_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7855 VPWR tdc0.w_dly_sig[29] tdc0.w_dly_sig_n[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7856 VPWR a_7607_7485# a_7775_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7857 a_21787_3543# tdc0.o_result[178] a_22021_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7858 VGND _051_ a_11405_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7859 VPWR a_26882_12559# clknet_4_14_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7860 _135_ a_12999_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7861 a_11513_18543# tdc0.w_dly_sig[94] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7862 a_9006_8319# a_8838_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7863 a_16121_9295# tdc0.o_result[27] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X7864 a_7515_10749# a_6651_10383# a_7258_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7865 VGND tdc0.w_dly_sig[4] a_27873_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7867 VGND tdc0.w_dly_sig_n[180] tdc0.w_dly_sig[182] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7868 a_30343_11293# a_30123_11305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X7869 a_18505_2223# tdc0.w_dly_sig[176] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7870 VGND a_22852_7093# clknet_4_9_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7871 a_17746_18111# a_17578_18365# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7872 tdc0.w_dly_sig[77] tdc0.w_dly_sig_n[76] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7873 VPWR tdc0.w_dly_sig_n[100] tdc0.w_dly_sig[102] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7874 a_16555_15797# clknet_4_12_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7876 a_6982_16341# a_6814_16367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7877 VGND a_17083_15101# a_17251_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7878 a_20421_6031# a_19867_6005# a_20074_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7879 a_23947_12015# _154_ a_24197_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7880 a_24731_11623# a_24827_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7881 VGND a_15059_10927# a_15227_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7882 tdc0.w_dly_sig_n[86] tdc0.w_dly_sig[85] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7883 tdc0.w_dly_sig[29] tdc0.w_dly_sig_n[27] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7884 a_7185_10749# a_6651_10383# a_7090_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7885 tdc0.w_dly_sig[26] tdc0.w_dly_sig_n[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7886 clknet_4_0_0_clk a_6476_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7887 VGND tdc0.w_dly_sig_n[133] tdc0.w_dly_sig[134] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7888 a_2842_7637# a_2674_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7889 VGND a_24731_14423# _127_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X7891 clknet_4_7_0_clk a_11812_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X7893 a_17559_12711# tdc0.o_result[99] a_17685_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X7894 VGND clknet_4_2_0_clk a_13091_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7895 a_7646_6397# a_7399_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7896 VPWR clknet_4_5_0_clk a_8031_16373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7897 a_16513_16189# a_16175_15975# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X7898 VPWR tdc0.o_result[174] a_19899_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7899 a_20709_9545# tdc0.o_result[65] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7900 a_11839_14191# a_11141_14197# a_11582_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7901 a_29987_11145# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7902 a_8914_17429# a_8746_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7903 tdc0.w_dly_sig[114] tdc0.w_dly_sig_n[113] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7904 tdc0.o_result[78] a_10351_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7906 a_11414_14191# a_10975_14197# a_11329_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7907 a_20039_5719# tdc0.o_result[20] a_20273_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7909 VPWR tdc0.w_dly_sig_n[61] tdc0.w_dly_sig[63] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7910 tdc0.w_dly_sig[139] tdc0.w_dly_sig_n[138] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7911 VPWR clknet_4_4_0_clk a_7387_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7912 a_26939_12247# a_27035_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7913 VPWR clknet_4_0_0_clk a_5823_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7914 VPWR tdc0.w_dly_sig_n[90] tdc0.w_dly_sig[91] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7915 tdc0.w_dly_sig[187] tdc0.w_dly_sig_n[186] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7916 a_1301_6031# tdc0.w_dly_sig[110] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7917 VGND tdc0.w_dly_sig[115] tdc0.w_dly_sig_n[116] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7918 tdc0.w_dly_sig[33] tdc0.w_dly_sig_n[32] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7919 VPWR a_7499_15253# a_7415_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7920 VGND a_9263_14013# a_9431_13915# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7921 VGND tdc0.w_dly_sig_n[149] tdc0.w_dly_sig[151] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7922 VGND clknet_4_5_0_clk a_6835_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7923 a_23811_1367# a_23907_1367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7924 VPWR clknet_4_3_0_clk a_10975_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7925 a_3870_11837# a_3431_11471# a_3785_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7926 a_30166_15253# a_29998_15279# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7927 VPWR _072_ a_7645_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7928 a_19268_591# a_18869_591# a_19142_957# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7929 VGND a_20258_10116# a_20187_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X7930 VGND tdc0.w_dly_sig[188] tdc0.w_dly_sig_n[188] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7931 VPWR tdc0.w_dly_sig_n[185] tdc0.w_dly_sig[186] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7932 a_2631_13103# a_1849_13109# a_2547_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7933 clknet_4_3_0_clk a_10506_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7935 VPWR a_22955_15253# a_22871_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7936 VGND tdc0.w_dly_sig[107] tdc0.w_dly_sig_n[107] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7938 VGND _050_ a_18029_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7939 a_16175_15975# a_16271_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7940 a_27873_10217# a_27326_9961# a_27526_10116# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X7941 VPWR a_15170_18111# a_15097_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7942 VGND a_6550_12559# clknet_4_4_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7943 VGND a_15779_17179# a_15737_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7945 tdc0.o_result[167] a_12283_3035# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7947 tdc0.w_dly_sig_n[95] tdc0.w_dly_sig[94] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7948 VGND a_25410_13103# clknet_4_15_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7949 a_14151_10535# tdc0.o_result[89] a_14385_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7950 VGND a_10018_2197# a_9976_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7951 _114_ a_15943_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X7952 tdc0.w_dly_sig_n[82] tdc0.w_dly_sig[81] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7953 a_13968_6281# _044_ a_13866_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X7954 a_4606_7485# a_4333_7119# a_4521_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7955 VPWR tdc0.w_dly_sig[150] tdc0.w_dly_sig_n[151] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7956 VPWR a_25318_7093# a_25247_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X7957 a_11030_8319# a_10862_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7958 VPWR a_7378_13103# clknet_4_5_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7959 VPWR clknet_4_8_0_clk a_22107_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7960 a_25230_8207# a_24915_8359# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7961 tdc0.w_dly_sig_n[42] tdc0.w_dly_sig[41] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7962 VPWR tdc0.w_dly_sig[36] tdc0.w_dly_sig_n[37] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7963 a_25428_7637# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7964 VPWR tdc0.w_dly_sig[164] tdc0.w_dly_sig_n[164] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7965 tdc0.w_dly_sig_n[68] tdc0.w_dly_sig[67] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7966 a_1554_6143# a_1386_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7967 VGND a_24915_8359# tdc0.o_result[22] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7968 a_19077_13469# _003_ a_19005_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7969 VGND a_19890_13103# clknet_4_13_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X7970 a_22898_10495# a_22730_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7971 VGND tdc0.w_dly_sig_n[5] tdc0.w_dly_sig[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7973 VPWR _050_ a_17047_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X7974 a_23478_6852# a_23278_6697# a_23627_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7975 VGND a_27135_7881# a_27142_7785# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7977 a_22546_16189# a_22273_15823# a_22461_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7978 VGND tdc0.w_dly_sig[149] tdc0.w_dly_sig_n[149] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7979 a_19652_13897# _004_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7980 a_9761_4399# a_9227_4405# a_9666_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7981 a_13717_16367# a_13183_16373# a_13622_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7982 VGND clknet_4_12_0_clk a_21923_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7983 VPWR a_25019_3529# a_25026_3433# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7984 a_19981_3677# tdc0.o_result[174] a_19899_3424# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7985 VGND _117_ a_15115_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7986 tdc0.w_dly_sig[160] tdc0.w_dly_sig_n[158] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7987 VGND a_27618_13380# a_27547_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X7988 a_22787_3133# a_22089_2767# a_22530_2879# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7989 VGND tdc0.w_dly_sig[154] tdc0.w_dly_sig_n[154] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7990 a_7239_16367# a_6541_16373# a_6982_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7991 a_8638_16341# a_8470_16367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7992 VPWR tdc0.w_dly_sig_n[181] tdc0.w_dly_sig[183] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7993 VPWR tdc0.o_result[156] a_12171_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7994 tdc0.w_dly_sig[119] tdc0.w_dly_sig_n[117] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7996 VGND a_14802_10901# a_14760_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7997 tdc0.o_result[173] a_16791_3035# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7998 VGND clknet_4_5_0_clk a_4995_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7999 tdc0.w_dly_sig_n[26] tdc0.w_dly_sig[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8000 tdc0.w_dly_sig_n[22] tdc0.w_dly_sig[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8001 a_11966_15279# a_11693_15285# a_11881_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8002 a_20893_14735# a_20727_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8003 a_22273_13109# a_22107_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8004 VGND a_10995_18267# a_10953_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8005 a_8481_10383# tdc0.o_result[128] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8006 a_27346_13469# a_27031_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X8007 VGND tdc0.w_dly_sig_n[135] tdc0.w_dly_sig[137] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8008 VPWR a_18489_9839# uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8009 tdc0.w_dly_sig_n[13] tdc0.w_dly_sig[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8010 VGND tdc0.w_dly_sig_n[48] tdc0.w_dly_sig[49] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8012 tdc0.o_result[106] a_2715_13915# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8013 a_6177_13103# tdc0.w_dly_sig[123] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8014 tdc0.w_dly_sig[158] tdc0.w_dly_sig_n[157] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8015 tdc0.w_dly_sig_n[38] tdc0.w_dly_sig[37] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8016 tdc0.o_result[36] a_23139_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8017 tdc0.w_dly_sig[22] tdc0.w_dly_sig_n[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8018 VGND a_17923_5719# _019_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X8019 VGND a_28503_12247# tdc0.o_result[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8020 a_23125_14557# _003_ a_23053_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8021 VPWR _054_ a_13735_14304# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X8022 VPWR a_7258_10495# a_7185_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8023 VPWR tdc0.w_dly_sig[12] tdc0.w_dly_sig_n[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8024 tdc0.w_dly_sig[186] tdc0.w_dly_sig_n[185] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8025 VGND tdc0.w_dly_sig[89] tdc0.w_dly_sig_n[90] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8026 VPWR a_17130_16885# a_17059_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8028 VGND tdc0.w_dly_sig_n[45] tdc0.w_dly_sig[46] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8029 a_4697_8041# a_3707_7669# a_4571_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8030 tdc0.o_result[36] a_23139_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8032 a_11747_9661# a_11049_9295# a_11490_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8033 a_14563_10383# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8034 VPWR a_18815_16341# a_18731_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8035 VPWR _172_ a_19255_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8036 a_27505_8207# a_26958_8481# a_27158_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X8037 VPWR tdc0.w_dly_sig_n[183] tdc0.w_dly_sig[185] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8038 a_7461_4405# a_7295_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8041 a_15695_17277# a_14913_16911# a_15611_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8042 VPWR tdc0.w_dly_sig[51] tdc0.w_dly_sig_n[51] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8043 tdc0.w_dly_sig_n[160] tdc0.w_dly_sig[160] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8044 VGND tdc0.w_dly_sig[175] tdc0.w_dly_sig_n[176] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8046 VPWR a_27342_7940# a_27271_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8047 a_16446_9071# _026_ a_16356_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X8048 tdc0.w_dly_sig_n[40] tdc0.w_dly_sig[40] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8049 a_23240_13897# _146_ a_23138_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X8050 a_2547_12925# a_1849_12559# a_2290_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8051 a_4061_7663# tdc0.w_dly_sig[118] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8053 a_5529_16189# a_4995_15823# a_5434_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8054 VGND a_30039_5211# a_29997_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8055 a_4329_11305# a_3339_10933# a_4203_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8056 a_26663_4007# a_26759_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8057 a_12253_4765# tdc0.o_result[156] a_12171_4512# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8058 _050_ a_16916_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8059 a_10034_3133# a_9761_2767# a_9949_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8060 VGND a_19211_7271# tdc0.o_result[27] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8061 VGND tdc0.w_dly_sig_n[117] tdc0.w_dly_sig[118] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8062 VGND a_18171_18267# a_18129_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8063 VGND a_2347_10901# a_2305_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8064 VPWR tdc0.w_dly_sig[183] tdc0.w_dly_sig_n[183] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8065 a_19310_703# a_19142_957# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8067 tdc0.w_dly_sig_n[14] tdc0.w_dly_sig[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8068 a_19927_18543# a_19145_18549# a_19843_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8069 a_18953_11721# _150_ a_19225_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8070 VPWR tdc0.w_dly_sig_n[161] tdc0.w_dly_sig[162] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8071 a_16547_7093# _021_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X8072 VGND clknet_4_12_0_clk a_17783_16373# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8073 a_12341_14735# tdc0.w_dly_sig[72] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8074 a_19505_12809# _201_ a_19433_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X8075 VPWR _054_ a_14563_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X8076 a_6476_6549# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8077 VGND tdc0.w_dly_sig_n[13] tdc0.w_dly_sig[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8078 a_6357_4399# a_5823_4405# a_6262_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8079 VGND tdc0.w_dly_sig[147] tdc0.w_dly_sig_n[147] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8080 VPWR a_8711_7663# a_8879_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8082 VGND _007_ a_14533_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8083 VGND a_30166_3285# a_30124_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8084 tdc0.w_dly_sig_n[177] tdc0.w_dly_sig[177] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8086 VPWR net3 a_16665_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8087 tdc0.w_dly_sig[160] tdc0.w_dly_sig_n[159] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8088 a_4295_11837# a_3431_11471# a_4038_11583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8089 VPWR clknet_4_5_0_clk a_6835_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8090 a_11966_15279# a_11527_15285# a_11881_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8091 a_19255_12015# _174_ a_19505_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8092 tdc0.w_dly_sig[6] tdc0.w_dly_sig_n[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8093 uo_out[5] a_24469_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8094 tdc0.w_dly_sig[80] tdc0.w_dly_sig_n[78] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8095 VGND a_19131_2741# a_19138_3041# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8097 tdc0.w_dly_sig[28] tdc0.w_dly_sig_n[27] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8099 VGND ui_in[7] a_18151_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X8100 tdc0.w_dly_sig[58] tdc0.w_dly_sig_n[57] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8101 tdc0.w_dly_sig_n[104] tdc0.w_dly_sig[103] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8102 tdc0.w_dly_sig_n[122] tdc0.w_dly_sig[121] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8103 VGND a_23478_6852# a_23407_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X8104 VGND tdc0.w_dly_sig[159] tdc0.w_dly_sig_n[160] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8105 a_27179_4777# a_27050_4521# a_26759_4631# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X8106 VPWR tdc0.o_result[41] a_24309_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X8107 a_18935_3543# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X8109 VPWR tdc0.w_dly_sig_n[189] tdc0.w_dly_sig[190] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8110 a_3651_14191# a_2787_14197# a_3394_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8111 VPWR a_18390_16341# a_18317_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8112 VGND tdc0.w_dly_sig_n[47] tdc0.w_dly_sig[48] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8113 a_23825_6953# a_23271_6793# a_23478_6852# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X8114 a_30166_15253# a_29998_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8115 VPWR a_26951_8969# a_26958_8873# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8116 a_23055_13103# a_22273_13109# a_22971_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8117 VPWR _152_ a_23947_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8118 a_11711_4512# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8119 a_16109_9545# tdc0.o_result[27] a_16025_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8120 VPWR tdc0.w_dly_sig_n[31] tdc0.w_dly_sig[33] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8121 VPWR tdc0.w_dly_sig[38] tdc0.w_dly_sig_n[38] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8122 a_17231_8457# _109_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X8123 tdc0.w_dly_sig_n[158] tdc0.w_dly_sig[157] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8124 a_24490_4917# a_24283_4917# a_24666_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X8125 tdc0.w_dly_sig_n[171] tdc0.w_dly_sig[170] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8126 tdc0.w_dly_sig[169] tdc0.w_dly_sig_n[168] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8127 VPWR tdc0.w_dly_sig_n[128] tdc0.w_dly_sig[130] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8129 VGND tdc0.w_dly_sig[85] tdc0.w_dly_sig_n[85] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8130 tdc0.w_dly_sig[98] tdc0.w_dly_sig_n[97] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8131 VPWR a_25962_12533# a_25891_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8132 VGND a_19225_11721# uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8133 tdc0.o_result[140] a_12007_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8134 VPWR tdc0.w_dly_sig[66] tdc0.w_dly_sig_n[66] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8135 VGND a_26882_12559# clknet_4_14_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8137 a_9815_7485# a_8951_7119# a_9558_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8138 tdc0.w_dly_sig_n[70] tdc0.w_dly_sig[70] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8139 VGND tdc0.w_dly_sig[35] a_22261_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X8141 VPWR tdc0.w_dly_sig_n[17] tdc0.w_dly_sig[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8142 a_15328_9839# _081_ a_15226_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X8143 tdc0.w_dly_sig[182] tdc0.w_dly_sig_n[181] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8145 tdc0.w_dly_sig_n[112] tdc0.w_dly_sig[112] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8146 VPWR tdc0.w_dly_sig[62] tdc0.w_dly_sig_n[62] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8147 VPWR _003_ a_21313_13441# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X8148 tdc0.w_dly_sig_n[161] tdc0.w_dly_sig[161] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8149 tdc0.w_dly_sig_n[182] tdc0.w_dly_sig[182] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8151 tdc0.w_dly_sig[162] tdc0.w_dly_sig_n[160] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8152 a_6541_16373# a_6375_16373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8153 tdc0.w_dly_sig[128] tdc0.w_dly_sig_n[127] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8154 a_4513_4777# a_3523_4405# a_4387_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8155 _180_ a_13367_9952# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X8156 a_19333_18543# tdc0.w_dly_sig[56] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8157 tdc0.w_dly_sig_n[91] tdc0.w_dly_sig[90] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8158 a_21523_13799# _001_ a_21697_13675# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X8159 VGND a_29982_12671# a_29940_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8160 VGND a_4755_3133# a_4923_3035# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8161 VGND tdc0.w_dly_sig_n[69] tdc0.w_dly_sig[71] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8162 a_27087_8207# a_26958_8481# a_26667_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X8163 a_2547_14013# a_1683_13647# a_2290_13759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8164 tdc0.w_dly_sig_n[186] tdc0.w_dly_sig[186] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8165 tdc0.w_dly_sig[7] tdc0.w_dly_sig_n[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8166 _013_ a_15530_6077# a_15793_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X8168 a_9263_9661# a_8565_9295# a_9006_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8169 a_10570_11583# a_10402_11837# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8170 a_23097_591# a_22107_591# a_22971_957# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8171 a_26769_9295# a_26215_9269# a_26422_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X8172 VGND _191_ a_6191_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8173 a_23662_11204# a_23455_11145# a_23838_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X8174 a_20654_5193# _196_ a_20574_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X8175 VGND a_10827_11837# a_10995_11739# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8176 tdc0.w_dly_sig_n[109] tdc0.w_dly_sig[109] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8177 a_20746_4399# _183_ a_20666_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X8178 tdc0.o_result[134] a_9983_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8179 clknet_0_clk a_16210_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X8180 a_8979_16367# a_8197_16373# a_8895_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8181 a_14274_13423# tdc0.o_result[139] a_14193_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X8182 a_19395_7895# tdc0.o_result[13] a_19629_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8183 a_8473_17461# a_8307_17461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8185 VGND a_26571_8359# tdc0.o_result[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8186 a_16799_8235# _021_ a_16713_8235# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X8187 VGND a_19671_10071# tdc0.o_result[33] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8188 VGND tdc0.w_dly_sig_n[176] tdc0.w_dly_sig[177] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8189 tdc0.w_dly_sig[18] tdc0.w_dly_sig_n[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8190 a_10961_4943# tdc0.w_dly_sig[143] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8191 a_17194_14165# a_17026_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8192 a_10494_15101# a_10055_14735# a_10409_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8193 a_14878_11721# tdc0.o_result[82] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X8194 tdc0.w_dly_sig_n[36] tdc0.w_dly_sig[35] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8195 VGND a_15611_17277# a_15779_17179# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8196 VPWR tdc0.w_dly_sig_n[107] tdc0.w_dly_sig[109] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8197 VPWR tdc0.w_dly_sig[52] tdc0.w_dly_sig_n[53] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8198 a_20425_12809# _194_ a_20175_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8199 a_18703_11471# _134_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X8201 tdc0.w_dly_sig_n[100] tdc0.w_dly_sig[100] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8202 VGND a_5123_8751# a_5291_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8203 VGND a_21334_14847# a_21292_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8204 a_7817_6031# a_7270_6305# a_7470_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X8205 tdc0.o_result[61] a_22771_17179# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8206 a_5115_11159# tdc0.o_result[132] a_5261_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8207 VGND _078_ a_14805_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X8208 a_29982_9813# a_29814_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8209 VPWR a_16737_9441# _037_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X8210 a_7331_15279# a_6633_15285# a_7074_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8211 tdc0.w_dly_sig_n[0] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8212 VGND a_26514_6575# clknet_4_11_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8213 tdc0.w_dly_sig[78] tdc0.w_dly_sig_n[77] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8214 a_14255_6835# _013_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X8215 a_2547_11837# a_1849_11471# a_2290_11583# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8216 VGND a_21327_17687# tdc0.o_result[54] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8217 VGND tdc0.w_dly_sig[89] tdc0.w_dly_sig_n[89] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8218 a_7734_4399# a_7295_4405# a_7649_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8219 a_8795_7663# a_8013_7669# a_8711_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8221 a_10405_12925# a_9871_12559# a_10310_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8222 VPWR a_25288_10357# _638_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X8224 VPWR tdc0.w_dly_sig_n[43] tdc0.w_dly_sig[45] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8225 tdc0.w_dly_sig[155] tdc0.w_dly_sig_n[153] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8226 a_29614_5055# a_29446_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8227 VGND tdc0.w_dly_sig_n[11] tdc0.w_dly_sig[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8228 a_20051_10057# clknet_4_13_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8229 a_14922_13897# _020_ a_14922_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X8230 tdc0.w_dly_sig_n[46] tdc0.w_dly_sig[46] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8231 a_20359_11471# _064_ a_20881_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8232 tdc0.w_dly_sig[185] tdc0.w_dly_sig_n[183] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8233 tdc0.w_dly_sig_n[52] tdc0.w_dly_sig[51] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8234 VPWR tdc0.w_dly_sig[87] tdc0.w_dly_sig_n[87] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8236 VGND tdc0.w_dly_sig[16] tdc0.w_dly_sig_n[17] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8237 clknet_4_12_0_clk a_21380_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8238 VGND a_19579_5719# _202_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X8239 a_13866_8457# _155_ a_13552_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X8240 VGND a_19221_13793# _209_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X8241 a_4038_11583# a_3870_11837# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8242 a_17048_4105# tdc0.o_result[138] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X8244 a_2122_14013# a_1849_13647# a_2037_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8245 clknet_4_8_0_clk a_21104_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8247 a_30239_12925# a_29375_12559# a_29982_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8248 tdc0.w_dly_sig_n[69] tdc0.w_dly_sig[68] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8249 VPWR a_4038_11583# a_3965_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8250 tdc0.w_dly_sig_n[3] tdc0.w_dly_sig[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8251 VPWR tdc0.w_dly_sig[141] tdc0.w_dly_sig_n[141] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8252 VGND tdc0.w_dly_sig_n[50] tdc0.w_dly_sig[51] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8253 a_24666_5309# a_24419_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X8254 tdc0.w_dly_sig[164] tdc0.w_dly_sig_n[163] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8255 tdc0.w_dly_sig[17] tdc0.w_dly_sig_n[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8256 VPWR a_4774_7231# a_4701_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8257 tdc0.w_dly_sig_n[113] tdc0.w_dly_sig[113] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8258 a_15097_2223# a_14563_2229# a_15002_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8259 a_29803_5705# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8260 VPWR tdc0.w_dly_sig_n[157] tdc0.w_dly_sig[159] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8261 a_29002_16733# a_28687_16599# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X8262 a_7902_4373# a_7734_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8263 VPWR a_19131_2741# a_19138_3041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8264 tdc0.w_dly_sig_n[33] tdc0.w_dly_sig[32] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8265 a_17493_17999# tdc0.w_dly_sig[58] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8266 VGND tdc0.w_dly_sig[21] tdc0.w_dly_sig_n[21] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8267 VGND net1 tdc0.w_dly_sig_n[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8268 tdc0.w_dly_sig_n[151] tdc0.w_dly_sig[150] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8270 a_13889_4765# _007_ a_13817_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8271 VPWR clknet_4_12_0_clk a_18979_18549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8272 VPWR tdc0.w_dly_sig_n[35] tdc0.w_dly_sig[36] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8273 a_20223_11293# a_20003_11305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X8274 VGND a_6395_3035# a_6353_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8275 a_29173_4943# a_29007_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8276 a_13722_8207# tdc0.o_result[117] a_13641_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X8277 a_25011_8181# a_25295_8181# a_25230_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X8278 tdc0.o_result[70] a_17619_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8279 a_30166_14165# a_29998_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8280 a_13530_2223# a_13091_2229# a_13445_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8281 tdc0.w_dly_sig[68] tdc0.w_dly_sig_n[66] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8282 VGND a_12759_9839# a_12927_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8284 VPWR _043_ a_12539_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X8285 tdc0.w_dly_sig[20] tdc0.w_dly_sig_n[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8286 VPWR tdc0.w_dly_sig_n[123] tdc0.w_dly_sig[124] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8287 a_22829_8751# tdc0.w_dly_sig[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8288 a_24131_9295# _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8289 a_11582_6549# a_11414_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8290 a_24639_15823# a_24419_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X8291 tdc0.w_dly_sig[50] tdc0.w_dly_sig_n[49] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8292 VGND tdc0.w_dly_sig_n[43] tdc0.w_dly_sig[44] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8293 VPWR tdc0.w_dly_sig_n[6] tdc0.w_dly_sig[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8294 VGND ui_in[3] a_15575_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X8295 a_13161_5865# a_12171_5493# a_13035_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8296 a_18489_9839# tdc0.o_result[3] a_18679_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X8297 VGND clknet_4_4_0_clk a_9319_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8298 tdc0.w_dly_sig[100] tdc0.w_dly_sig_n[98] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8299 VPWR tdc0.w_dly_sig_n[151] tdc0.w_dly_sig[152] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8300 VPWR tdc0.w_dly_sig_n[18] tdc0.w_dly_sig[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8301 VPWR clknet_4_12_0_clk a_22107_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8302 VGND tdc0.w_dly_sig[7] tdc0.w_dly_sig_n[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8303 VPWR tdc0.w_dly_sig[100] tdc0.w_dly_sig_n[100] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8304 a_4655_17277# a_3873_16911# a_4571_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8305 a_13275_7776# _024_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8306 a_25375_12711# a_25471_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8309 VPWR net6 a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X8310 tdc0.o_result[167] a_12283_3035# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8311 tdc0.w_dly_sig_n[118] tdc0.w_dly_sig[118] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8312 tdc0.w_dly_sig[66] tdc0.w_dly_sig_n[64] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8313 VPWR a_25111_11445# a_25118_11745# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8314 a_9393_4405# a_9227_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8315 VGND tdc0.w_dly_sig_n[55] tdc0.w_dly_sig[57] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8316 VPWR tdc0.w_dly_sig_n[85] tdc0.w_dly_sig[86] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8317 VPWR tdc0.w_dly_sig[34] a_20605_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X8318 tdc0.w_dly_sig[48] tdc0.w_dly_sig_n[46] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8319 a_27965_13481# a_27418_13225# a_27618_13380# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X8320 tdc0.w_dly_sig_n[7] tdc0.w_dly_sig[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8321 a_14250_17429# a_14082_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8322 a_13354_13423# _140_ a_13600_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X8323 a_18309_11721# _141_ a_18237_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X8324 tdc0.w_dly_sig_n[85] tdc0.w_dly_sig[84] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8325 tdc0.w_dly_sig[154] tdc0.w_dly_sig_n[153] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8326 tdc0.w_dly_sig_n[10] tdc0.w_dly_sig[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8327 a_16198_3133# a_15759_2767# a_16113_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8328 tdc0.o_result[184] a_22955_3035# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8329 a_24363_4007# tdc0.o_result[186] a_24597_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8330 a_11251_4512# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8331 a_18977_4719# _008_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X8332 VGND a_22633_4917# _133_ VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8333 VGND a_1995_5487# a_2163_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8334 VGND a_4111_5487# a_4279_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8335 a_12578_8457# _166_ a_12264_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X8336 VPWR a_27618_13380# a_27547_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8338 a_17467_10357# _018_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X8340 a_15009_15823# tdc0.w_dly_sig[68] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8341 a_14082_17455# a_13809_17461# a_13997_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8342 a_5717_2767# tdc0.w_dly_sig[157] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8344 a_19255_12809# _201_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8345 VPWR a_10478_12671# a_10405_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8346 VPWR tdc0.w_dly_sig[140] tdc0.w_dly_sig_n[140] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8347 VPWR tdc0.w_dly_sig[142] tdc0.w_dly_sig_n[142] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8348 VGND tdc0.w_dly_sig_n[22] tdc0.w_dly_sig[24] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8349 tdc0.o_result[95] a_10719_17179# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8350 a_10543_4221# a_9761_3855# a_10459_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8351 tdc0.w_dly_sig[25] tdc0.w_dly_sig_n[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8352 a_17567_9447# _019_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X8353 a_18843_13335# tdc0.o_result[60] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8354 a_8979_3311# a_8197_3317# a_8895_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8355 VPWR a_22809_13793# _149_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X8356 a_29814_12925# a_29375_12559# a_29729_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8357 VPWR clknet_4_4_0_clk a_4259_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8358 a_23903_18775# a_23999_18775# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X8359 VPWR a_10202_2879# a_10129_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8360 tdc0.w_dly_sig[1] tdc0.w_dly_sig_n[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8361 a_6503_4221# a_5639_3855# a_6246_3967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8363 a_14151_10535# _054_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X8364 a_7860_4777# a_7461_4405# a_7734_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8365 VGND tdc0.w_dly_sig[19] tdc0.w_dly_sig_n[20] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8366 a_22461_13103# tdc0.w_dly_sig[37] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8367 a_12426_16189# a_12153_15823# a_12341_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8368 tdc0.w_dly_sig_n[93] tdc0.w_dly_sig[93] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8369 tdc0.w_dly_sig[97] tdc0.w_dly_sig_n[95] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8370 a_9466_8725# a_9298_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8371 a_9849_9129# a_8859_8757# a_9723_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8372 VGND tdc0.w_dly_sig[152] tdc0.w_dly_sig_n[152] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8373 a_4701_7485# a_4167_7119# a_4606_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8375 a_9021_16745# a_8031_16373# a_8895_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8376 VGND tdc0.w_dly_sig_n[149] tdc0.w_dly_sig[150] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8377 VPWR tdc0.w_dly_sig[190] tdc0.w_dly_sig_n[190] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8378 VPWR _042_ a_17231_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X8379 VPWR a_25835_9447# tdc0.o_result[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8380 a_13537_16367# tdc0.w_dly_sig[90] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8381 VPWR tdc0.w_dly_sig[182] tdc0.w_dly_sig_n[183] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8383 VPWR net1 tdc0.w_dly_sig_n[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8384 VPWR tdc0.w_dly_sig_n[34] tdc0.w_dly_sig[35] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8385 VGND tdc0.w_dly_sig[188] a_28425_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X8386 VPWR tdc0.w_dly_sig_n[161] tdc0.w_dly_sig[163] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8387 tdc0.w_dly_sig_n[114] tdc0.w_dly_sig[114] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8388 a_10129_3133# a_9595_2767# a_10034_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8390 a_25755_15797# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8391 VPWR tdc0.w_dly_sig_n[70] tdc0.w_dly_sig[72] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8392 a_11329_6575# tdc0.w_dly_sig[140] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8393 a_14989_8353# _100_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X8394 a_1669_10927# tdc0.w_dly_sig[111] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8396 VGND tdc0.w_dly_sig_n[13] tdc0.w_dly_sig[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8397 a_23384_13647# tdc0.o_result[36] a_22809_13793# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X8398 uo_out[0] a_20881_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8399 _190_ a_19163_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X8400 a_22374_2500# a_22167_2441# a_22550_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X8401 _011_ net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8403 a_17167_15101# a_16385_14735# a_17083_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8404 a_4330_3133# a_4057_2767# a_4245_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8405 a_30541_11471# a_29994_11745# a_30194_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X8406 tdc0.w_dly_sig_n[134] tdc0.w_dly_sig[133] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8407 a_2842_7637# a_2674_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8408 a_8565_15823# a_8399_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8409 a_28503_13335# a_28599_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X8410 a_7902_4373# a_7734_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8411 a_17681_13103# _020_ a_17765_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8412 a_6906_15279# a_6633_15285# a_6821_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8413 VPWR clknet_0_clk a_21380_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8414 a_22891_14423# tdc0.o_result[52] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8415 VGND a_12851_11837# a_13019_11739# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8416 a_23999_2741# a_24290_3041# a_24241_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8417 _193_ a_23110_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X8418 a_19395_6807# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X8419 a_8286_7663# a_7847_7669# a_8201_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8420 a_25713_16189# a_25375_15975# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X8422 VGND a_17691_6281# _033_ VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
X8423 a_10862_8573# a_10589_8207# a_10777_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8425 VGND tdc0.w_dly_sig[135] tdc0.w_dly_sig_n[136] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8426 tdc0.w_dly_sig[89] tdc0.w_dly_sig_n[87] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8427 tdc0.w_dly_sig_n[61] tdc0.w_dly_sig[61] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8428 tdc0.w_dly_sig[142] tdc0.w_dly_sig_n[141] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8429 tdc0.w_dly_sig_n[144] tdc0.w_dly_sig[143] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8430 VPWR _039_ a_13184_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X8431 a_18843_13335# tdc0.o_result[60] a_19077_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8433 a_14507_17455# a_13809_17461# a_14250_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8434 clknet_4_15_0_clk a_25410_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8435 tdc0.w_dly_sig[7] tdc0.w_dly_sig_n[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8436 a_3302_15253# a_3134_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8437 a_13656_2601# a_13257_2229# a_13530_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8438 tdc0.o_result[107] a_2715_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8439 VPWR a_9983_7387# a_9899_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8440 tdc0.w_dly_sig[110] tdc0.w_dly_sig_n[108] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8441 VPWR clknet_4_4_0_clk a_1683_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8443 tdc0.w_dly_sig[133] tdc0.w_dly_sig_n[131] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8444 tdc0.o_result[83] a_11087_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8445 VGND tdc0.w_dly_sig[123] tdc0.w_dly_sig_n[123] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8446 VPWR a_19798_7093# a_19727_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8447 tdc0.w_dly_sig[12] tdc0.w_dly_sig_n[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8448 tdc0.w_dly_sig_n[102] tdc0.w_dly_sig[102] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8449 tdc0.w_dly_sig[105] tdc0.w_dly_sig_n[103] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8450 a_10221_17277# a_9687_16911# a_10126_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8451 a_9347_14013# a_8565_13647# a_9263_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8452 a_3394_3285# a_3226_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8453 _191_ a_8491_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8454 VPWR a_10735_14013# a_10903_13915# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8455 VPWR tdc0.w_dly_sig[104] tdc0.w_dly_sig_n[105] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8456 VPWR a_2547_13103# a_2715_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8457 a_20529_2767# tdc0.w_dly_sig[178] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8458 VPWR a_9263_8573# a_9431_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8459 a_25375_15975# a_25471_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X8460 a_3134_15279# a_2861_15285# a_3049_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8461 a_30102_4676# a_29902_4521# a_30251_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X8462 VGND tdc0.w_dly_sig_n[2] tdc0.w_dly_sig[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8463 tdc0.w_dly_sig[19] tdc0.w_dly_sig_n[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8465 VGND a_4571_17277# a_4739_17179# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8466 a_5349_15823# tdc0.w_dly_sig[104] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8467 VGND clknet_4_13_0_clk a_20727_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8468 _070_ a_19982_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X8469 VPWR a_8159_4399# a_8327_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8470 VGND a_2547_13103# a_2715_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8471 VGND _047_ a_5341_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X8472 a_8159_4399# a_7461_4405# a_7902_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8473 VGND tdc0.w_dly_sig[143] tdc0.w_dly_sig_n[143] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8474 a_30166_3285# a_29998_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8475 VPWR a_26882_12559# clknet_4_14_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8476 a_23907_1367# a_24191_1353# a_24126_1501# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X8477 a_18703_13647# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8478 tdc0.w_dly_sig[173] tdc0.w_dly_sig_n[172] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8480 a_26978_4765# a_26663_4631# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X8481 VGND tdc0.w_dly_sig_n[65] tdc0.w_dly_sig[67] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8482 VGND _041_ a_13722_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X8483 VPWR a_25019_13621# a_25026_13921# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8484 tdc0.w_dly_sig_n[54] tdc0.w_dly_sig[53] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8485 a_20337_15657# a_19347_15285# a_20211_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8486 VPWR tdc0.w_dly_sig[93] tdc0.w_dly_sig_n[93] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8487 VGND tdc0.w_dly_sig_n[44] tdc0.w_dly_sig[45] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8488 VPWR a_24005_8725# _189_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X8489 a_16324_2767# a_15925_2767# a_16198_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8490 VPWR tdc0.w_dly_sig_n[114] tdc0.w_dly_sig[115] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8491 a_22891_14423# tdc0.o_result[52] a_23125_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8492 VPWR a_14011_5487# _025_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8494 VPWR _026_ a_12723_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X8496 a_9390_7485# a_8951_7119# a_9305_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8497 a_6476_7637# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8498 tdc0.w_dly_sig[102] tdc0.w_dly_sig_n[100] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8499 VPWR a_16555_15797# a_16562_16097# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8500 a_11839_6575# a_11141_6581# a_11582_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8501 VGND tdc0.w_dly_sig_n[191] tdc0.w_dly_sig[192] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R23 VGND uio_out[3] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X8502 a_3651_3311# a_2953_3317# a_3394_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8503 a_13722_12559# _200_ a_13968_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X8504 a_25471_12533# a_25755_12533# a_25690_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X8505 VPWR a_10719_17179# a_10635_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8506 VPWR a_7442_14847# a_7369_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8507 a_24197_12015# _154_ a_23947_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8508 tdc0.w_dly_sig[113] tdc0.w_dly_sig_n[111] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8509 VPWR tdc0.w_dly_sig[168] tdc0.w_dly_sig_n[168] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8510 a_14917_17999# tdc0.w_dly_sig[93] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8512 _064_ _001_ a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X8513 VGND a_26203_7271# tdc0.o_result[19] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8514 tdc0.w_dly_sig[21] tdc0.w_dly_sig_n[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8515 VPWR _054_ a_18703_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X8516 VPWR tdc0.w_dly_sig_n[127] tdc0.w_dly_sig[129] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8517 a_16845_10927# tdc0.o_result[42] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8518 VGND a_19497_5089# _137_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X8519 tdc0.w_dly_sig_n[55] tdc0.w_dly_sig[55] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8520 tdc0.o_result[113] a_2163_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8521 a_12621_10383# tdc0.o_result[93] a_12539_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8522 a_30423_3311# a_29725_3317# a_30166_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8524 tdc0.o_result[26] a_24059_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8525 _170_ a_12999_8867# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X8526 a_16911_15823# a_16691_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X8527 VGND a_30347_10357# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8528 VPWR tdc0.w_dly_sig_n[36] tdc0.w_dly_sig[38] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8530 VPWR tdc0.w_dly_sig_n[154] tdc0.w_dly_sig[155] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8531 VPWR a_4755_3133# a_4923_3035# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8532 VGND tdc0.w_dly_sig[187] a_25573_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X8533 a_22550_2223# a_22303_2601# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X8534 tdc0.w_dly_sig_n[130] tdc0.w_dly_sig[130] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8535 VPWR a_11087_15003# a_11003_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8536 tdc0.o_result[9] a_30591_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8537 a_15729_13647# _022_ a_15657_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8538 VPWR a_16210_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8539 VPWR clknet_4_7_0_clk a_14655_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8540 a_16850_13423# _049_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X8541 _198_ a_12999_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X8542 a_16945_4943# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
R24 tt_um_hpretl_tt06_tdc_v1_14.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X8543 tdc0.w_dly_sig[144] tdc0.w_dly_sig_n[142] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8544 a_27503_5705# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8545 VPWR tdc0.w_dly_sig[106] tdc0.w_dly_sig_n[107] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8546 tdc0.w_dly_sig_n[140] tdc0.w_dly_sig[139] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8548 a_22086_4399# a_21647_4405# a_22001_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8549 a_17691_14985# _065_ a_17773_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X8550 VGND clknet_4_14_0_clk a_22291_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8551 VGND tdc0.w_dly_sig[82] tdc0.w_dly_sig_n[82] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8552 VGND tdc0.w_dly_sig_n[39] tdc0.w_dly_sig[40] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8554 a_11435_7119# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8555 a_4609_8207# a_4443_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8556 a_9466_8725# a_9298_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8557 a_8838_16189# a_8399_15823# a_8753_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8558 a_3559_15279# a_2861_15285# a_3302_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8559 VPWR a_11287_8573# a_11455_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8560 tdc0.w_dly_sig[126] tdc0.w_dly_sig_n[125] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8561 tdc0.w_dly_sig_n[144] tdc0.w_dly_sig[144] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8562 a_3134_15279# a_2695_15285# a_3049_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8563 a_18869_591# a_18703_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8564 a_23903_4007# tdc0.o_result[179] a_24137_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8565 a_30102_4676# a_29895_4617# a_30278_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X8566 VPWR clknet_4_10_0_clk a_29651_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8567 a_24837_4943# a_24290_5217# a_24490_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X8568 VGND _007_ a_13429_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8569 VGND tdc0.w_dly_sig[38] a_22813_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X8570 _090_ a_14563_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X8571 a_2547_13103# a_1683_13109# a_2290_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8573 a_8251_12015# a_7553_12021# a_7994_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8574 VGND tdc0.w_dly_sig_n[88] tdc0.w_dly_sig[89] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8575 VPWR a_16175_15975# tdc0.o_result[64] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8576 a_26598_9661# a_26351_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X8578 a_16757_17455# tdc0.w_dly_sig[59] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8579 VGND tdc0.w_dly_sig[105] tdc0.w_dly_sig_n[105] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8580 _081_ a_15023_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X8581 a_29729_9839# tdc0.w_dly_sig[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8582 a_10225_13647# tdc0.w_dly_sig[83] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8583 VPWR a_25962_4917# a_25891_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8584 a_22987_6807# a_23278_6697# a_23229_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8585 VGND a_19890_13103# clknet_4_13_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8586 a_24735_3543# a_25019_3529# a_24954_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X8587 tdc0.w_dly_sig[84] tdc0.w_dly_sig_n[83] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8588 a_8412_8041# a_8013_7669# a_8286_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8589 tdc0.w_dly_sig_n[179] tdc0.w_dly_sig[179] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8590 tdc0.w_dly_sig[167] tdc0.w_dly_sig_n[165] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8591 a_18785_14985# tdc0.o_result[121] a_18703_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8592 a_7994_11989# a_7826_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8593 VPWR a_10570_11583# a_10497_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8594 net1 a_30347_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8595 a_8546_2197# a_8378_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8597 VPWR a_10294_17023# a_10221_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8598 VGND _059_ a_16645_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X8599 tdc0.w_dly_sig_n[4] tdc0.w_dly_sig[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8600 _122_ a_12539_6688# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X8602 VGND tdc0.w_dly_sig[137] tdc0.w_dly_sig_n[138] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8603 VPWR a_22852_7093# clknet_4_9_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8605 VGND clknet_4_13_0_clk a_19531_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8606 VPWR a_21104_6005# clknet_4_8_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8607 a_24977_14013# a_24639_13799# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X8609 _011_ a_16495_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8610 VGND tdc0.w_dly_sig[58] tdc0.w_dly_sig_n[59] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8611 tdc0.w_dly_sig_n[104] tdc0.w_dly_sig[104] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8612 tdc0.o_result[108] a_2715_11739# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8613 a_18292_4399# _143_ a_18190_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X8614 a_24009_11305# a_23455_11145# a_23662_11204# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X8615 VPWR a_4498_2879# a_4425_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8616 a_22891_6807# a_22987_6807# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X8617 a_23591_11305# a_23462_11049# a_23171_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X8618 VPWR _060_ a_21787_3543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X8619 VGND tdc0.w_dly_sig[48] tdc0.w_dly_sig_n[48] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8620 VPWR tdc0.w_dly_sig_n[178] tdc0.w_dly_sig[180] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8621 VPWR tdc0.o_result[96] a_16219_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8623 VPWR tdc0.w_dly_sig[21] a_26309_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X8624 a_22603_17277# a_21905_16911# a_22346_17023# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8625 _086_ a_11803_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X8626 VGND tdc0.w_dly_sig[9] tdc0.w_dly_sig_n[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8627 a_8838_9661# a_8565_9295# a_8753_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8628 _094_ a_16679_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X8630 VPWR clknet_4_13_0_clk a_20727_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8631 VPWR a_30039_5211# a_29955_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8632 a_27219_5719# a_27503_5705# a_27438_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X8633 VPWR clknet_4_13_0_clk a_22107_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8634 tdc0.w_dly_sig_n[66] tdc0.w_dly_sig[66] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8635 a_16941_14191# tdc0.w_dly_sig[71] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8636 VGND _204_ a_19058_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X8637 a_2290_13759# a_2122_14013# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8638 VGND tdc0.w_dly_sig_n[98] tdc0.w_dly_sig[99] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8639 VGND tdc0.w_dly_sig[140] tdc0.w_dly_sig_n[141] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8640 tdc0.w_dly_sig_n[125] tdc0.w_dly_sig[125] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8641 VGND a_10506_7119# clknet_4_3_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8642 VPWR clknet_0_clk a_11812_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8643 VGND a_16366_2879# a_16324_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8645 a_2122_13103# a_1849_13109# a_2037_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8646 tdc0.w_dly_sig_n[174] tdc0.w_dly_sig[174] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8647 a_20721_9295# tdc0.o_result[185] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X8648 tdc0.w_dly_sig_n[142] tdc0.w_dly_sig[141] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8649 VGND a_5491_15101# a_5659_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8650 VPWR a_22971_13103# a_23139_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8651 VPWR a_19015_2223# a_19183_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8653 tdc0.w_dly_sig[42] tdc0.w_dly_sig_n[40] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8654 tdc0.w_dly_sig_n[90] tdc0.w_dly_sig[89] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8655 VPWR clknet_4_4_0_clk a_6651_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8656 a_9516_7119# a_9117_7119# a_9390_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8657 tdc0.w_dly_sig_n[64] tdc0.w_dly_sig[64] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8658 tdc0.w_dly_sig[46] tdc0.w_dly_sig_n[45] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8659 VGND tdc0.w_dly_sig_n[70] tdc0.w_dly_sig[71] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8660 VGND tdc0.w_dly_sig_n[188] tdc0.w_dly_sig[189] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8662 a_16894_12015# _061_ a_16645_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X8663 a_3693_10927# tdc0.w_dly_sig[117] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8664 a_29423_6196# tdc0.w_dly_sig[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8665 a_18785_13647# tdc0.o_result[95] a_18703_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8666 a_20181_3855# _043_ a_20109_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8667 tdc0.o_result[62] a_23139_16091# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8668 a_11690_3133# a_11251_2767# a_11605_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8669 a_4054_4221# a_3615_3855# a_3969_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8670 a_19881_10633# tdc0.o_result[144] a_19797_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8671 VGND a_24283_15797# a_24290_16097# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8672 tdc0.w_dly_sig_n[130] tdc0.w_dly_sig[129] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8673 VPWR a_26755_7895# tdc0.o_result[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8674 VGND tdc0.w_dly_sig[54] tdc0.w_dly_sig_n[54] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8675 a_25379_14709# a_25663_14709# a_25598_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X8676 tdc0.o_result[86] a_14675_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8677 tdc0.w_dly_sig_n[110] tdc0.w_dly_sig[109] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8678 VGND tdc0.w_dly_sig_n[106] tdc0.w_dly_sig[107] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8679 a_12999_3424# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8680 VPWR a_6671_4123# a_6587_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8682 a_22362_3133# a_21923_2767# a_22277_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8683 uo_out[6] a_19777_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8684 tdc0.w_dly_sig[153] tdc0.w_dly_sig_n[152] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8685 VGND tdc0.w_dly_sig[139] tdc0.w_dly_sig_n[139] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8686 tdc0.w_dly_sig_n[108] tdc0.w_dly_sig[107] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8689 a_28007_2767# a_27878_3041# a_27587_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X8690 VGND a_24490_18820# a_24419_18921# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X8691 tdc0.w_dly_sig_n[26] tdc0.w_dly_sig[26] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8692 VPWR tdc0.w_dly_sig[189] a_27597_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X8693 VPWR a_24191_1353# a_24198_1257# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8694 a_7657_11471# tdc0.o_result[114] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X8695 a_7691_7485# a_6909_7119# a_7607_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8696 a_24488_8207# tdc0.o_result[26] a_23913_8353# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X8697 a_19163_9545# _181_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8698 VPWR clknet_4_13_0_clk a_16403_17461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8700 a_22212_4777# a_21813_4405# a_22086_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8701 VPWR a_25778_1653# a_25707_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8702 VPWR clknet_4_7_0_clk a_14563_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8703 a_15380_6895# tdc0.o_result[25] a_14805_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X8704 a_17704_17999# a_17305_17999# a_17578_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8705 a_2217_11837# a_1683_11471# a_2122_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8706 a_23455_11145# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8708 VGND a_20417_4373# _185_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X8709 tdc0.w_dly_sig[32] tdc0.w_dly_sig_n[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8710 VPWR tdc0.w_dly_sig[181] a_24745_1513# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X8711 VGND tdc0.w_dly_sig_n[138] tdc0.w_dly_sig[140] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8712 a_8838_16189# a_8565_15823# a_8753_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8713 tdc0.w_dly_sig_n[133] tdc0.w_dly_sig[132] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8714 a_12356_9545# tdc0.o_result[73] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X8715 a_2861_15285# a_2695_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8716 a_26583_7093# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8717 a_25253_8573# a_24915_8359# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X8718 tdc0.o_result[139] a_12007_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8719 a_29871_5309# a_29007_4943# a_29614_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8720 tdc0.w_dly_sig[36] tdc0.w_dly_sig_n[34] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8721 tdc0.w_dly_sig[61] tdc0.w_dly_sig_n[60] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8723 VGND a_14255_6835# _035_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8724 a_16465_3677# _038_ a_16393_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8725 a_14349_3677# _025_ a_14277_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8726 a_16401_6691# net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8727 VPWR a_17159_18517# a_17075_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8728 tdc0.w_dly_sig[11] tdc0.w_dly_sig_n[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8729 VPWR tdc0.w_dly_sig[73] tdc0.w_dly_sig_n[74] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8730 tdc0.o_result[16] a_30683_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8732 a_21349_1679# a_20359_1679# a_21223_2045# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8733 a_11322_9661# a_10883_9295# a_11237_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8734 VGND a_21380_14165# clknet_4_12_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8735 VPWR a_26514_6575# clknet_4_11_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8736 VPWR tdc0.w_dly_sig_n[1] tdc0.w_dly_sig[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8737 tdc0.w_dly_sig_n[52] tdc0.w_dly_sig[52] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8738 VPWR a_16991_957# a_17159_859# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8739 a_17577_2601# a_16587_2229# a_17451_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8741 VPWR a_15163_3543# _123_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X8742 _064_ net5 a_17703_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8743 VPWR tdc0.w_dly_sig[136] tdc0.w_dly_sig_n[137] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8744 VPWR a_7407_16341# a_7323_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8746 a_4425_3133# a_3891_2767# a_4330_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8747 a_15054_6575# _079_ a_14805_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X8748 VGND tdc0.w_dly_sig[33] tdc0.w_dly_sig_n[34] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8749 a_17464_4105# _103_ a_17362_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X8750 tdc0.w_dly_sig_n[188] tdc0.w_dly_sig[188] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8752 _171_ a_4995_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X8753 tdc0.w_dly_sig_n[38] tdc0.w_dly_sig[38] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8754 VPWR tdc0.w_dly_sig[77] tdc0.w_dly_sig_n[77] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8755 tdc0.w_dly_sig_n[175] tdc0.w_dly_sig[174] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8756 VPWR a_9063_3285# a_8979_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8757 a_21813_4405# a_21647_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8758 tdc0.w_dly_sig[59] tdc0.w_dly_sig_n[58] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8760 VPWR tdc0.w_dly_sig_n[16] tdc0.w_dly_sig[17] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8761 a_5602_15935# a_5434_16189# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8762 tdc0.w_dly_sig_n[85] tdc0.w_dly_sig[85] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8763 a_16293_591# a_16127_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8764 VGND a_30166_15253# a_30124_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8765 VPWR tdc0.w_dly_sig[106] tdc0.w_dly_sig_n[106] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8766 a_5721_11721# _023_ a_5805_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8768 a_14591_15279# a_13809_15285# a_14507_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8769 VPWR clknet_4_2_0_clk a_9227_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8770 tdc0.w_dly_sig[116] tdc0.w_dly_sig_n[114] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8771 tdc0.w_dly_sig[35] tdc0.w_dly_sig_n[33] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8772 a_25379_14709# a_25670_15009# a_25621_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8773 VPWR a_9339_17429# a_9255_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8774 a_29729_12559# tdc0.w_dly_sig[44] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8775 clknet_4_4_0_clk a_6550_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8776 a_19255_12809# _209_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X8777 VGND a_4479_4221# a_4647_4123# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8778 tdc0.w_dly_sig_n[16] tdc0.w_dly_sig[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8779 tdc0.w_dly_sig[129] tdc0.w_dly_sig_n[128] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8780 a_3651_14191# a_2953_14197# a_3394_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8781 tdc0.w_dly_sig_n[62] tdc0.w_dly_sig[62] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8782 a_21313_13441# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X8783 a_7185_10933# a_7019_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8784 a_4613_8751# tdc0.w_dly_sig[115] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8786 a_12610_5487# a_12337_5493# a_12525_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8787 VPWR a_18383_8983# _095_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X8788 VPWR tdc0.w_dly_sig_n[109] tdc0.w_dly_sig[111] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8789 VGND clknet_4_5_0_clk a_6375_16373# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8790 clknet_0_clk a_16210_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8792 a_21843_11305# a_21707_11145# a_21423_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X8793 a_21697_13675# _058_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X8795 VPWR _035_ a_23303_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X8796 tdc0.w_dly_sig[180] tdc0.w_dly_sig_n[179] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8797 tdc0.w_dly_sig[75] tdc0.w_dly_sig_n[74] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8798 tdc0.w_dly_sig[34] tdc0.w_dly_sig_n[33] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8799 VGND tdc0.w_dly_sig[168] tdc0.w_dly_sig_n[169] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8802 VGND tdc0.w_dly_sig_n[124] tdc0.w_dly_sig[125] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8803 a_7198_6031# a_6883_6183# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X8804 VPWR a_19591_7093# a_19598_7393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8805 VPWR tdc0.w_dly_sig[92] tdc0.w_dly_sig_n[92] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8806 tdc0.w_dly_sig_n[5] tdc0.w_dly_sig[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8807 tdc0.w_dly_sig[13] tdc0.w_dly_sig_n[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8809 VGND tdc0.w_dly_sig[157] tdc0.w_dly_sig_n[157] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8810 VGND a_2163_5461# a_2121_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8811 VPWR tdc0.w_dly_sig_n[104] tdc0.w_dly_sig[106] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8812 VGND clknet_4_5_0_clk a_8307_17461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8814 VGND a_9558_7231# a_9516_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8815 VGND net4 a_17953_591# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X8816 a_29614_5055# a_29446_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8817 VGND tdc0.w_dly_sig[134] tdc0.w_dly_sig_n[134] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8818 a_9723_8751# a_8859_8757# a_9466_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8819 VPWR clknet_0_clk a_19890_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8820 tdc0.w_dly_sig[31] tdc0.w_dly_sig_n[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8822 tdc0.w_dly_sig[96] tdc0.w_dly_sig_n[95] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8823 a_30541_11305# a_29994_11049# a_30194_11204# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X8825 a_4180_3855# a_3781_3855# a_4054_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8826 tdc0.w_dly_sig_n[132] tdc0.w_dly_sig[132] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8827 a_11816_2767# a_11417_2767# a_11690_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8828 _047_ a_15101_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.247 ps=2.06 w=0.65 l=0.15
X8829 a_23407_6953# a_23278_6697# a_22987_6807# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X8830 VGND clknet_4_4_0_clk a_3431_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8831 VPWR tdc0.o_result[33] a_15328_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X8832 a_27043_4617# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8833 VGND tdc0.w_dly_sig[53] a_23733_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X8834 a_23933_16367# tdc0.w_dly_sig[52] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8835 tdc0.w_dly_sig_n[53] tdc0.w_dly_sig[52] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8836 a_1386_6397# a_1113_6031# a_1301_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8837 VGND tdc0.w_dly_sig[12] tdc0.w_dly_sig_n[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8838 a_21883_2455# a_22174_2345# a_22125_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8840 a_11329_7663# tdc0.w_dly_sig[138] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8841 tdc0.w_dly_sig[55] tdc0.w_dly_sig_n[54] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8842 a_15381_12015# _004_ a_15465_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8844 VPWR a_20315_7895# _160_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X8846 VPWR a_27319_10057# a_27326_9961# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8847 a_22488_2767# a_22089_2767# a_22362_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8848 a_19245_9545# _189_ a_19163_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X8849 a_19005_13469# _054_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X8850 _154_ a_22751_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X8851 tdc0.w_dly_sig_n[91] tdc0.w_dly_sig[91] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8852 VPWR a_30194_11204# a_30123_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8853 VPWR a_6476_6549# clknet_4_0_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8854 tdc0.o_result[115] a_3267_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8855 a_10478_12671# a_10310_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8856 tdc0.o_result[87] a_13019_16091# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8857 a_24218_18909# a_23903_18775# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X8859 a_7216_10383# a_6817_10383# a_7090_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8860 tdc0.w_dly_sig_n[24] tdc0.w_dly_sig[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8861 tdc0.w_dly_sig_n[138] tdc0.w_dly_sig[138] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8862 _184_ a_19899_3424# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X8863 clknet_4_8_0_clk a_21104_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8864 a_27461_5487# a_27123_5719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X8865 VPWR tdc0.w_dly_sig[4] a_27873_10217# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X8866 a_24144_16745# a_23745_16373# a_24018_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8867 _638_.X a_25288_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8868 VGND clknet_4_2_0_clk a_14563_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8869 VGND clknet_4_11_0_clk a_29559_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8873 a_11414_6397# a_10975_6031# a_11329_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8874 a_9006_15935# a_8838_16189# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8876 VPWR tdc0.w_dly_sig[154] tdc0.w_dly_sig_n[155] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8877 a_18479_6895# _010_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8878 VGND a_15351_7093# _026_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X8879 tdc0.w_dly_sig[83] tdc0.w_dly_sig_n[81] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8880 tdc0.w_dly_sig_n[131] tdc0.w_dly_sig[130] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8881 tdc0.w_dly_sig_n[176] tdc0.w_dly_sig[175] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8882 tdc0.w_dly_sig_n[87] tdc0.w_dly_sig[87] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8883 VPWR tdc0.w_dly_sig_n[84] tdc0.w_dly_sig[85] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8884 tdc0.w_dly_sig[150] tdc0.w_dly_sig_n[148] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8886 a_17949_16373# a_17783_16373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8887 VPWR tdc0.o_result[71] a_13643_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8888 tdc0.w_dly_sig[145] tdc0.w_dly_sig_n[143] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8889 a_26138_12925# a_25891_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X8890 _179_ a_12815_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X8891 tdc0.w_dly_sig[183] tdc0.w_dly_sig_n[181] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8892 a_25375_3677# a_25155_3689# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X8893 a_10041_16911# tdc0.w_dly_sig[96] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8894 a_26769_9295# a_26222_9569# a_26422_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X8895 clknet_4_15_0_clk a_25410_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8896 a_18317_2229# a_18151_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8897 VGND a_20379_15253# a_20337_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8898 a_26150_9295# a_25835_9447# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X8899 a_17451_14191# a_16587_14197# a_17194_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8900 VGND a_29871_5309# a_30039_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8901 tdc0.w_dly_sig[32] tdc0.w_dly_sig_n[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8902 VGND tdc0.w_dly_sig_n[96] tdc0.w_dly_sig[97] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8903 a_12426_15101# a_11987_14735# a_12341_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8904 VPWR tdc0.w_dly_sig_n[123] tdc0.w_dly_sig[125] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8905 VGND tdc0.w_dly_sig_n[56] tdc0.w_dly_sig[58] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8906 tdc0.w_dly_sig[51] tdc0.w_dly_sig_n[50] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8907 a_21327_11159# a_21423_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X8908 a_26978_3855# a_26663_4007# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X8909 VGND a_25835_9447# tdc0.o_result[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8910 a_11448_9295# a_11049_9295# a_11322_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8911 VPWR tdc0.w_dly_sig_n[50] tdc0.w_dly_sig[52] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8912 a_10506_7119# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X8913 VGND _125_ a_15115_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8914 VPWR a_6550_12559# clknet_4_4_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8916 a_21591_15101# a_20727_14735# a_21334_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8917 tdc0.o_result[72] a_15963_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8918 VPWR a_25870_14709# a_25799_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8919 VGND tdc0.w_dly_sig_n[40] tdc0.w_dly_sig[41] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8920 a_24381_9545# _090_ a_24653_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8921 a_19671_10071# a_19767_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X8922 a_21975_12533# a_22266_12833# a_22217_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8923 a_24013_11445# _014_ a_24170_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X8925 VGND a_21707_17673# a_21714_17577# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8926 a_18479_6895# _010_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8927 VPWR tdc0.w_dly_sig[114] tdc0.w_dly_sig_n[114] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8928 tdc0.w_dly_sig[15] tdc0.w_dly_sig_n[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8929 a_23999_18775# a_24290_18665# a_24241_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8930 _085_ a_16205_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.247 ps=2.06 w=0.65 l=0.15
X8931 VPWR tdc0.w_dly_sig_n[166] tdc0.w_dly_sig[167] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8932 VPWR tdc0.w_dly_sig[88] tdc0.w_dly_sig_n[89] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8933 a_27127_13335# a_27411_13321# a_27346_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X8934 a_30166_3285# a_29998_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8935 VGND tdc0.w_dly_sig_n[170] tdc0.w_dly_sig[171] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8936 a_20709_9545# tdc0.o_result[185] a_20625_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8937 VGND a_18703_12559# _003_ VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8938 VPWR a_26790_7093# a_26719_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8939 VGND clknet_0_clk a_25428_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X8940 VPWR tdc0.w_dly_sig[49] tdc0.w_dly_sig_n[49] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8941 tdc0.w_dly_sig_n[73] tdc0.w_dly_sig[72] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8942 VGND tdc0.w_dly_sig[111] tdc0.w_dly_sig_n[111] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8943 a_22261_11305# a_21707_11145# a_21914_11204# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X8944 a_5115_7485# a_4333_7119# a_5031_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8945 a_21261_15101# a_20727_14735# a_21166_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8946 VGND a_25019_13621# a_25026_13921# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8947 VGND tdc0.w_dly_sig_n[105] tdc0.w_dly_sig[106] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8948 a_6430_13077# a_6262_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8949 a_12897_2767# tdc0.o_result[166] a_12815_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8950 a_29515_4631# a_29611_4631# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8951 a_14878_11721# tdc0.o_result[34] a_14721_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8955 VGND a_22955_15253# a_22913_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8956 tdc0.w_dly_sig[93] tdc0.w_dly_sig_n[92] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8957 a_15575_13647# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8959 a_22595_4399# a_21813_4405# a_22511_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8960 tdc0.w_dly_sig_n[53] tdc0.w_dly_sig[53] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8961 _023_ a_13997_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.247 ps=2.06 w=0.65 l=0.15
X8962 a_13722_9295# _179_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X8963 VGND tdc0.w_dly_sig[124] tdc0.w_dly_sig_n[124] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8964 VGND a_25375_12711# tdc0.o_result[38] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8965 tdc0.o_result[75] a_12927_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8966 a_28599_13335# a_28890_13225# a_28841_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8967 tdc0.w_dly_sig[24] tdc0.w_dly_sig_n[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8969 VPWR tdc0.w_dly_sig_n[167] tdc0.w_dly_sig[169] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8970 VGND tdc0.w_dly_sig[59] tdc0.w_dly_sig_n[60] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8973 VGND tdc0.w_dly_sig[126] tdc0.w_dly_sig_n[127] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8974 VPWR a_30194_11445# a_30123_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8975 VPWR tdc0.w_dly_sig_n[71] tdc0.w_dly_sig[72] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8976 a_4146_7663# a_3873_7669# a_4061_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8977 a_27411_13321# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8978 VPWR _016_ a_20359_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8979 VGND a_11260_5461# clknet_4_2_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8980 a_22672_591# a_22273_591# a_22546_957# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8981 VGND a_11858_2879# a_11816_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8982 tdc0.w_dly_sig_n[67] tdc0.w_dly_sig[66] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8983 a_21765_3855# _056_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X8984 a_19150_8207# _159_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X8985 a_18679_9839# tdc0.o_result[3] a_18489_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X8986 VGND tdc0.w_dly_sig_n[83] tdc0.w_dly_sig[85] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8988 a_29982_9813# a_29814_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8989 a_6725_14197# a_6559_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8990 clknet_4_11_0_clk a_26514_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8991 a_4609_8207# a_4443_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8992 a_16113_2767# tdc0.w_dly_sig[174] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8993 a_24033_14735# tdc0.o_result[63] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X8994 tdc0.w_dly_sig_n[6] tdc0.w_dly_sig[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8995 a_22799_17687# a_22895_17687# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X8996 a_10585_3855# a_9595_3855# a_10459_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8997 VPWR a_10827_11837# a_10995_11739# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8998 a_14989_8353# _098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X9000 a_3946_10901# a_3778_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9001 VGND a_22530_2879# a_22488_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9002 VGND tdc0.w_dly_sig_n[146] tdc0.w_dly_sig[147] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9003 tdc0.w_dly_sig[151] tdc0.w_dly_sig_n[149] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9004 a_11812_13621# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9005 a_5989_13109# a_5823_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9006 a_22089_15285# a_21923_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9007 a_12693_10383# _034_ a_12621_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9008 tdc0.o_result[123] a_7591_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9009 VGND tdc0.w_dly_sig[63] tdc0.w_dly_sig_n[64] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9011 a_4882_6397# a_4443_6031# a_4797_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9012 a_14884_11471# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X9013 a_19773_9441# _033_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9014 tdc0.o_result[171] a_14583_3035# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9016 tdc0.w_dly_sig_n[146] tdc0.w_dly_sig[146] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9017 a_21843_17833# a_21714_17577# a_21423_17687# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X9018 a_19701_15279# tdc0.w_dly_sig[66] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9019 VGND a_23082_8725# a_23040_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9020 a_11540_6031# a_11141_6031# a_11414_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9021 a_27150_17277# a_26903_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X9022 a_12115_3133# a_11417_2767# a_11858_2879# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9023 a_14103_4943# _024_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9024 VPWR tdc0.w_dly_sig[87] tdc0.w_dly_sig_n[88] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9025 a_20359_11721# _029_ a_20609_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9026 _124_ a_11435_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X9028 a_27526_10116# a_27326_9961# a_27675_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X9030 VGND a_7470_6005# a_7399_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X9031 a_11839_7663# a_10975_7669# a_11582_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9032 VPWR a_22466_12533# a_22395_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X9033 a_25431_8207# a_25295_8181# a_25011_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9034 tdc0.w_dly_sig[132] tdc0.w_dly_sig_n[131] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9035 a_26299_11445# a_26583_11445# a_26518_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X9037 VGND clknet_0_clk a_6476_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X9038 a_18140_9071# tdc0.o_result[122] a_17565_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X9039 a_24381_9545# _071_ a_24131_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9040 VPWR a_16210_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9041 VPWR a_29871_5309# a_30039_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9042 VGND a_18815_16341# a_18773_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9043 tdc0.w_dly_sig[72] tdc0.w_dly_sig_n[70] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9044 VPWR a_25755_15797# a_25762_16097# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9047 VGND a_3083_4373# a_3041_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9048 VGND tdc0.w_dly_sig[122] tdc0.w_dly_sig_n[123] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9049 tdc0.o_result[105] a_3819_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9050 tdc0.w_dly_sig_n[185] tdc0.w_dly_sig[184] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9051 VPWR tdc0.w_dly_sig_n[122] tdc0.w_dly_sig[123] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9052 tdc0.w_dly_sig[121] tdc0.w_dly_sig_n[119] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9053 a_10494_15101# a_10221_14735# a_10409_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9055 VGND a_11490_9407# a_11448_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9057 tdc0.w_dly_sig_n[191] tdc0.w_dly_sig[191] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9058 VGND _104_ a_17218_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X9059 VPWR a_28503_13335# tdc0.o_result[42] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9060 VPWR a_21334_14847# a_21261_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9061 clknet_4_15_0_clk a_25410_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9062 VPWR tdc0.w_dly_sig[163] tdc0.w_dly_sig_n[163] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9065 VPWR a_30166_8725# a_30093_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9066 VGND _093_ a_16679_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9067 a_7378_13103# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9069 a_8933_9661# a_8399_9295# a_8838_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9070 tdc0.w_dly_sig_n[143] tdc0.w_dly_sig[143] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9071 VGND _193_ a_23855_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9072 VPWR tdc0.w_dly_sig[6] a_27873_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9073 VGND clknet_4_7_0_clk a_13643_18549# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9075 VPWR _025_ a_11679_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X9076 VGND a_14703_3543# _073_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X9077 VPWR a_14123_2197# a_14039_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9078 VPWR tdc0.w_dly_sig[33] a_20421_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9080 clknet_4_13_0_clk a_19890_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9081 VPWR tdc0.w_dly_sig[22] tdc0.w_dly_sig_n[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9082 a_15709_6281# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X9083 tdc0.w_dly_sig_n[56] tdc0.w_dly_sig[55] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9084 VPWR a_10919_15101# a_11087_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9086 VGND a_6687_5487# a_6855_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9088 clknet_4_0_0_clk a_6476_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9089 VPWR a_17567_9447# _020_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X9090 VPWR a_18758_2197# a_18685_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9091 VPWR a_26882_12559# clknet_4_14_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9092 _192_ a_6191_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X9093 tdc0.w_dly_sig[81] tdc0.w_dly_sig_n[80] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9094 VGND tdc0.w_dly_sig[34] a_20605_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X9095 VGND tdc0.w_dly_sig[116] tdc0.w_dly_sig_n[116] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9096 VPWR tdc0.w_dly_sig_n[7] tdc0.w_dly_sig[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9097 VPWR a_25375_15975# tdc0.o_result[48] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9100 a_7507_14191# a_6725_14197# a_7423_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9103 VGND tdc0.w_dly_sig_n[145] tdc0.w_dly_sig[146] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9104 a_7221_6397# a_6883_6183# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X9106 VGND a_25283_14887# tdc0.o_result[41] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9107 a_24827_11445# a_25118_11745# a_25069_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9108 a_17317_6281# net2 a_17233_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9109 a_10317_11471# tdc0.w_dly_sig[81] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9110 VPWR tdc0.w_dly_sig_n[172] tdc0.w_dly_sig[173] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9111 VGND a_6227_3133# a_6395_3035# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9112 tdc0.w_dly_sig_n[35] tdc0.w_dly_sig[34] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9113 tdc0.o_result[141] a_10259_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9114 a_7277_7485# a_6743_7119# a_7182_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9115 tdc0.w_dly_sig_n[56] tdc0.w_dly_sig[56] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9116 _111_ a_17498_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X9117 a_17773_6281# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9119 a_2037_11471# tdc0.w_dly_sig[109] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9120 VPWR a_9891_8725# a_9807_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9121 VPWR tdc0.w_dly_sig[130] tdc0.w_dly_sig_n[131] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9123 tdc0.w_dly_sig_n[178] tdc0.w_dly_sig[177] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9124 a_5307_6397# a_4443_6031# a_5050_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9125 VGND net5 a_17593_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9126 VPWR a_27250_3829# a_27179_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X9127 VGND a_1979_6299# a_1937_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9128 a_2658_4373# a_2490_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9129 a_18857_13647# _058_ a_18785_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9130 VPWR a_1554_6143# a_1481_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9131 VGND tdc0.w_dly_sig[91] tdc0.w_dly_sig_n[92] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9132 _032_ a_15483_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X9133 a_19798_7093# a_19591_7093# a_19974_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X9134 clknet_4_7_0_clk a_11812_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9135 tdc0.o_result[71] a_13019_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9136 a_22790_5193# tdc0.o_result[180] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X9137 VPWR tdc0.w_dly_sig[60] a_17477_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9138 VGND tdc0.w_dly_sig[167] tdc0.w_dly_sig_n[167] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9139 VGND a_17507_1143# net5 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X9140 a_26583_7093# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9141 tdc0.w_dly_sig[184] tdc0.w_dly_sig_n[182] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9142 a_9305_7119# tdc0.w_dly_sig[135] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9143 VPWR a_2715_12827# a_2631_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9144 a_26974_16885# a_26767_16885# a_27150_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X9145 a_23634_7637# a_23466_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9146 a_20697_12809# _064_ a_20175_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9147 VPWR a_4479_4221# a_4647_4123# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9148 a_5008_6031# a_4609_6031# a_4882_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9149 a_16639_16885# a_16923_16885# a_16858_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X9150 VPWR tdc0.w_dly_sig_n[97] tdc0.w_dly_sig[98] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9151 a_7699_3133# a_7001_2767# a_7442_2879# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9152 a_8105_2229# a_7939_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9153 VPWR tdc0.w_dly_sig[187] tdc0.w_dly_sig_n[187] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9154 VGND _019_ a_17139_8759# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X9155 tdc0.w_dly_sig[57] tdc0.w_dly_sig_n[56] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9156 net1 a_30347_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9157 tdc0.w_dly_sig[38] tdc0.w_dly_sig_n[36] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9158 a_10294_17023# a_10126_17277# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9159 a_17059_16911# a_16930_17185# a_16639_16885# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X9160 VGND a_21391_1947# a_21349_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9161 clknet_4_11_0_clk a_26514_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9162 clknet_0_clk a_16210_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9163 tdc0.w_dly_sig_n[25] tdc0.w_dly_sig[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9164 tdc0.w_dly_sig_n[27] tdc0.w_dly_sig[26] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9166 tdc0.w_dly_sig[95] tdc0.w_dly_sig_n[93] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9167 a_17773_6281# _030_ a_17691_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9168 VGND a_9006_9407# a_8964_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9169 a_22461_15823# tdc0.w_dly_sig[63] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9171 a_23457_3677# _056_ a_23385_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9172 _110_ a_17231_8457# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X9173 a_30093_8751# a_29559_8757# a_29998_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9174 tdc0.w_dly_sig_n[84] tdc0.w_dly_sig[84] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9175 a_5575_15101# a_4793_14735# a_5491_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9176 a_11605_1135# tdc0.w_dly_sig[167] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9177 a_15609_4971# _005_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X9178 VPWR a_30239_9839# a_30407_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9179 a_10129_11471# a_9963_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9180 tdc0.w_dly_sig[157] tdc0.w_dly_sig_n[156] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9181 VGND clknet_4_3_0_clk a_10607_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9182 VGND a_19890_13103# clknet_4_13_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9183 a_19773_9441# _175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X9184 a_2248_13481# a_1849_13109# a_2122_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9185 VPWR _040_ a_15391_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9186 VGND a_30591_8725# a_30549_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9187 a_23351_14423# _003_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X9188 a_10202_3967# a_10034_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9189 VPWR clknet_4_9_0_clk a_21647_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9190 VPWR a_14675_17429# a_14591_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9191 a_10275_2223# a_9411_2229# a_10018_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9192 a_17023_5487# net6 a_16665_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9193 VPWR a_17559_12711# _112_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X9194 a_27873_12393# a_27319_12233# a_27526_12292# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X9195 a_16991_957# a_16293_591# a_16734_703# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9196 a_16734_18517# a_16566_18543# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9197 VGND a_23662_11204# a_23591_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X9198 a_11881_15279# tdc0.w_dly_sig[86] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9199 a_3226_3311# a_2787_3317# a_3141_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9201 VPWR a_30423_3311# a_30591_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9202 a_12526_9295# tdc0.o_result[73] a_12445_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X9203 a_18685_2223# a_18151_2229# a_18590_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9204 VGND _007_ a_15695_4971# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X9205 a_25295_8181# clknet_4_11_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9206 tdc0.w_dly_sig_n[159] tdc0.w_dly_sig[158] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9207 a_22895_17687# a_23186_17577# a_23137_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9208 tdc0.o_result[88] a_15779_17179# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9209 VGND a_21039_3133# a_21207_3035# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9210 a_17026_2223# a_16753_2229# a_16941_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9211 a_6813_4777# a_5823_4405# a_6687_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9212 a_29067_16585# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9213 VGND a_30347_10357# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9215 _031_ a_18737_6059# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X9216 _042_ a_16401_6691# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X9218 VPWR a_13019_15003# a_12935_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9219 tdc0.w_dly_sig[31] tdc0.w_dly_sig_n[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9220 tdc0.w_dly_sig_n[93] tdc0.w_dly_sig[92] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9221 a_16566_18543# a_16293_18549# a_16481_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9222 VGND a_7378_13103# clknet_4_5_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9224 VGND a_19591_7093# a_19598_7393# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9225 VPWR a_2290_12671# a_2217_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9226 a_6979_6005# a_7263_6005# a_7198_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X9228 VPWR a_25375_8983# _106_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X9229 a_12092_15657# a_11693_15285# a_11966_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9230 a_11724_18921# a_11325_18549# a_11598_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9231 a_20713_1679# tdc0.w_dly_sig[179] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9232 VGND clknet_4_7_0_clk a_13643_17461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9233 a_13081_8867# _169_ a_12999_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9234 a_14437_8725# _115_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X9235 VPWR a_5602_15935# a_5529_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9236 tdc0.w_dly_sig_n[77] tdc0.w_dly_sig[77] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9237 VGND tdc0.w_dly_sig_n[179] tdc0.w_dly_sig[181] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9238 VPWR a_20074_11204# a_20003_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X9239 VPWR tdc0.o_result[165] a_12999_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X9240 VGND tdc0.w_dly_sig_n[148] tdc0.w_dly_sig[149] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9241 tdc0.w_dly_sig_n[48] tdc0.w_dly_sig[48] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9242 a_11045_14735# a_10055_14735# a_10919_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9243 a_18847_2741# a_19138_3041# a_19089_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9244 a_23811_1367# a_23907_1367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9245 a_13449_10205# tdc0.o_result[78] a_13367_9952# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9246 VPWR tdc0.w_dly_sig_n[48] tdc0.w_dly_sig[50] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9248 VGND net24 a_30357_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X9249 tdc0.w_dly_sig_n[9] tdc0.w_dly_sig[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9250 a_22833_12015# _153_ a_22751_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9251 VGND a_18703_10383# _058_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X9252 a_1481_6397# a_947_6031# a_1386_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9253 VPWR a_10903_13915# a_10819_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9254 a_12851_16189# a_12153_15823# a_12594_15935# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9256 VPWR a_4314_7637# a_4241_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9257 a_13613_3677# _025_ a_13541_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9259 a_28599_12247# a_28883_12233# a_28818_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X9260 a_23947_12335# _064_ a_24469_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9261 VPWR tdc0.w_dly_sig[3] tdc0.w_dly_sig_n[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9262 VGND a_9063_3285# a_9021_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9263 _144_ a_17875_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X9264 VGND a_16193_8725# _113_ VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X9265 a_8746_17455# a_8473_17461# a_8661_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9266 a_20039_5719# _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X9267 VGND a_16210_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9268 a_16850_13423# tdc0.o_result[104] a_16769_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X9269 a_17383_5095# net3 a_17557_4971# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X9270 a_30423_15279# a_29725_15285# a_30166_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9271 a_22714_13077# a_22546_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9272 VGND tdc0.w_dly_sig_n[180] tdc0.w_dly_sig[181] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9273 tdc0.w_dly_sig[67] tdc0.w_dly_sig_n[66] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9274 a_12609_2601# a_11619_2229# a_12483_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9275 VGND tdc0.w_dly_sig[159] tdc0.w_dly_sig_n[159] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9276 VPWR tdc0.w_dly_sig_n[28] tdc0.w_dly_sig[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9277 tdc0.w_dly_sig[115] tdc0.w_dly_sig_n[114] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9278 tdc0.w_dly_sig[124] tdc0.w_dly_sig_n[122] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9279 a_20697_12809# tdc0.o_result[7] a_20175_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X9280 a_29607_11159# a_29703_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9281 VGND tdc0.w_dly_sig_n[135] tdc0.w_dly_sig[136] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9282 a_16381_10383# tdc0.o_result[76] a_15943_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9283 VPWR a_14507_15279# a_14675_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9284 VPWR a_19855_8359# _159_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X9286 a_15351_7093# _006_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X9287 VPWR a_22971_16189# a_23139_16091# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9288 VGND a_30102_4676# a_30031_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X9289 VGND a_20395_14191# a_20563_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9290 a_19797_10633# _015_ a_19715_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9291 tdc0.w_dly_sig_n[157] tdc0.w_dly_sig[156] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9292 VPWR tdc0.w_dly_sig[129] tdc0.w_dly_sig_n[130] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9293 tdc0.w_dly_sig_n[3] tdc0.w_dly_sig[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9294 VGND a_14507_15279# a_14675_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9295 VGND tdc0.w_dly_sig_n[37] tdc0.w_dly_sig[39] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9296 a_11417_1141# a_11251_1141# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9297 VPWR tdc0.w_dly_sig_n[11] tdc0.w_dly_sig[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9298 VPWR a_3727_15253# a_3643_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9299 a_11605_2767# tdc0.w_dly_sig[168] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9300 VGND tdc0.w_dly_sig_n[113] tdc0.w_dly_sig[115] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9303 VPWR tdc0.w_dly_sig_n[170] tdc0.w_dly_sig[172] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9305 a_15795_12925# a_15097_12559# a_15538_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9306 tdc0.w_dly_sig_n[96] tdc0.w_dly_sig[95] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9307 VPWR tdc0.o_result[164] a_12999_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9308 VPWR _064_ a_18679_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9309 a_16566_18543# a_16127_18549# a_16481_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9310 a_30031_4777# a_29902_4521# a_29611_4631# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X9311 VGND tdc0.w_dly_sig[21] a_26309_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X9312 VPWR a_19487_6183# tdc0.o_result[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9313 a_17083_15101# a_16385_14735# a_16826_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9314 tdc0.w_dly_sig[45] tdc0.w_dly_sig_n[43] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9315 tdc0.w_dly_sig[161] tdc0.w_dly_sig_n[159] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9316 tdc0.w_dly_sig[163] tdc0.w_dly_sig_n[162] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9317 VPWR tdc0.w_dly_sig_n[98] tdc0.w_dly_sig[100] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9318 VGND a_20697_12809# uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9319 a_29982_12671# a_29814_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9320 a_10953_11471# a_9963_11471# a_10827_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9321 a_22277_2767# tdc0.w_dly_sig[185] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9322 a_8803_2223# a_8105_2229# a_8546_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9323 VPWR a_21523_13799# _068_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X9324 a_17691_14985# _065_ a_17773_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9325 tdc0.w_dly_sig[191] tdc0.w_dly_sig_n[190] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9326 tdc0.w_dly_sig[136] tdc0.w_dly_sig_n[134] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9327 tdc0.w_dly_sig[8] tdc0.w_dly_sig_n[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9328 VPWR tdc0.w_dly_sig_n[93] tdc0.w_dly_sig[94] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9329 a_4866_11989# a_4698_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9330 VPWR a_23455_11145# a_23462_11049# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9331 a_30423_3311# a_29559_3317# a_30166_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9332 a_12999_4399# _039_ a_13082_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X9334 a_6814_16367# a_6375_16373# a_6729_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9335 VPWR _197_ a_19505_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X9336 a_29725_3317# a_29559_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9337 VPWR tdc0.w_dly_sig[28] tdc0.w_dly_sig_n[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9338 VPWR tdc0.w_dly_sig_n[116] tdc0.w_dly_sig[117] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9339 a_25111_11445# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9341 VGND clknet_4_5_0_clk a_2695_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9342 VGND a_21380_14165# clknet_4_12_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9343 a_17415_10927# _092_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9344 VPWR tdc0.w_dly_sig[42] a_26217_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9345 tdc0.w_dly_sig[122] tdc0.w_dly_sig_n[120] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9346 tdc0.w_dly_sig_n[9] tdc0.w_dly_sig[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9347 VPWR tdc0.w_dly_sig[56] tdc0.w_dly_sig_n[57] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9349 a_4698_12015# a_4425_12021# a_4613_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9350 tdc0.w_dly_sig_n[14] tdc0.w_dly_sig[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9351 tdc0.w_dly_sig_n[74] tdc0.w_dly_sig[73] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9352 a_3352_3689# a_2953_3317# a_3226_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9353 a_8746_17455# a_8307_17461# a_8661_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9355 a_11555_5309# a_10773_4943# a_11471_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9356 a_17010_17429# a_16842_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9357 a_9263_14013# a_8565_13647# a_9006_13759# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9358 VPWR tdc0.w_dly_sig[169] tdc0.w_dly_sig_n[170] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9360 tdc0.w_dly_sig[69] tdc0.w_dly_sig_n[68] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9361 VGND clknet_4_8_0_clk a_21923_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9362 VGND a_25203_3829# a_25210_4129# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9363 VGND _004_ a_20153_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X9364 a_11237_9295# tdc0.w_dly_sig[74] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9365 VPWR tdc0.w_dly_sig_n[119] tdc0.w_dly_sig[120] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9366 VGND tdc0.w_dly_sig_n[14] tdc0.w_dly_sig[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9368 a_27587_2741# a_27878_3041# a_27829_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9369 tdc0.w_dly_sig[113] tdc0.w_dly_sig_n[112] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9370 tdc0.o_result[171] a_14583_3035# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9371 tdc0.w_dly_sig[52] tdc0.w_dly_sig_n[50] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9372 clknet_4_4_0_clk a_6550_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9373 VPWR a_23271_6793# a_23278_6697# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9374 a_1485_5487# tdc0.w_dly_sig[150] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9376 a_3601_5487# tdc0.w_dly_sig[148] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9377 tdc0.w_dly_sig_n[149] tdc0.w_dly_sig[149] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9378 VPWR a_29987_11445# a_29994_11745# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9379 a_6883_6183# a_6979_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9380 a_11371_8573# a_10589_8207# a_11287_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9381 a_12670_9545# _086_ a_12356_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X9382 VPWR tdc0.w_dly_sig[47] a_29621_16745# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9384 VGND tdc0.w_dly_sig_n[0] tdc0.w_dly_sig[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9385 a_30166_7637# a_29998_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9386 VGND tdc0.w_dly_sig_n[91] tdc0.w_dly_sig[92] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9387 a_14507_15279# a_13643_15285# a_14250_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9388 VGND tdc0.w_dly_sig[160] tdc0.w_dly_sig_n[160] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9389 a_4241_7663# a_3707_7669# a_4146_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9391 VGND tdc0.w_dly_sig_n[82] tdc0.w_dly_sig[83] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9392 VPWR tdc0.w_dly_sig_n[120] tdc0.w_dly_sig[121] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9393 tdc0.w_dly_sig_n[168] tdc0.w_dly_sig[168] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9394 VGND tdc0.w_dly_sig[135] tdc0.w_dly_sig_n[135] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9395 VGND clknet_4_9_0_clk a_22475_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9396 a_19697_14197# a_19531_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9397 VPWR tdc0.o_result[170] a_17047_3424# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9398 a_14257_4943# _024_ a_14185_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9399 VPWR _007_ a_14379_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9400 tdc0.w_dly_sig_n[89] tdc0.w_dly_sig[88] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9401 tdc0.w_dly_sig[11] tdc0.w_dly_sig_n[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9402 a_6729_16367# tdc0.w_dly_sig[99] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9403 a_11329_6031# tdc0.w_dly_sig[141] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9404 tdc0.o_result[99] a_9431_16091# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9405 VPWR tdc0.w_dly_sig[142] tdc0.w_dly_sig_n[143] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9406 a_24527_16367# a_23745_16373# a_24443_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9407 VGND _009_ a_17691_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X9409 tdc0.w_dly_sig_n[72] tdc0.w_dly_sig[71] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9410 tdc0.w_dly_sig[111] tdc0.w_dly_sig_n[109] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9411 tdc0.w_dly_sig_n[168] tdc0.w_dly_sig[167] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9412 VPWR tdc0.w_dly_sig[153] tdc0.w_dly_sig_n[153] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9413 VPWR _007_ a_14931_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9414 a_21423_11159# a_21714_11049# a_21665_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9415 a_18151_10383# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9416 VPWR clknet_4_8_0_clk a_18151_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9417 a_14177_15279# a_13643_15285# a_14082_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9418 _016_ a_19715_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X9419 VGND a_10627_4123# a_10585_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9420 a_24731_11623# a_24827_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9421 VGND tdc0.w_dly_sig_n[115] tdc0.w_dly_sig[117] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9422 tdc0.o_result[120] a_5935_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9423 a_2953_3317# a_2787_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9424 a_22346_17023# a_22178_17277# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9425 VGND clknet_4_3_0_clk a_10883_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9426 tdc0.w_dly_sig[114] tdc0.w_dly_sig_n[112] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9427 VPWR tdc0.w_dly_sig_n[0] tdc0.w_dly_sig[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9428 tdc0.w_dly_sig_n[117] tdc0.w_dly_sig[117] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9429 a_9298_8751# a_8859_8757# a_9213_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9430 tdc0.w_dly_sig_n[92] tdc0.w_dly_sig[92] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9431 tdc0.w_dly_sig[161] tdc0.w_dly_sig_n[160] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9432 VGND tdc0.w_dly_sig_n[184] tdc0.w_dly_sig[186] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9433 VPWR a_5475_6299# a_5391_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9434 VPWR a_9063_16341# a_8979_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9435 a_24283_2741# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9436 VPWR clknet_4_8_0_clk a_18703_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9437 VPWR a_23913_8353# _109_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X9438 tdc0.w_dly_sig_n[187] tdc0.w_dly_sig[186] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9440 VGND clknet_4_5_0_clk a_8399_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9441 a_22796_4943# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X9443 VGND tdc0.w_dly_sig_n[117] tdc0.w_dly_sig[119] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9445 VPWR tdc0.w_dly_sig_n[75] tdc0.w_dly_sig[76] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9446 VPWR a_18737_6059# _031_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X9447 tdc0.w_dly_sig[40] tdc0.w_dly_sig_n[38] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9448 a_5050_6143# a_4882_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9449 VPWR tdc0.w_dly_sig_n[102] tdc0.w_dly_sig[103] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9450 VPWR a_8419_11989# a_8335_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9451 a_24827_7093# a_25118_7393# a_25069_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9452 VGND clknet_0_clk a_6476_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X9453 VPWR _018_ a_18151_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9455 a_3965_11837# a_3431_11471# a_3870_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9456 a_15163_3543# tdc0.o_result[171] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9457 VPWR tdc0.w_dly_sig_n[71] tdc0.w_dly_sig[73] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9458 a_19395_3543# tdc0.o_result[175] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9459 a_22714_15935# a_22546_16189# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9460 a_17231_8457# _101_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9461 VGND _054_ a_12693_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9462 a_17129_3677# tdc0.o_result[170] a_17047_3424# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9463 VPWR tdc0.w_dly_sig[24] a_24837_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9464 tdc0.w_dly_sig[193] tdc0.w_dly_sig_n[191] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9466 VGND clknet_4_5_0_clk a_8031_16373# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9467 a_17267_17455# a_16569_17461# a_17010_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9468 VPWR clknet_4_4_0_clk a_1683_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9469 a_1481_10933# a_1315_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9470 tdc0.w_dly_sig_n[15] tdc0.w_dly_sig[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9471 a_17305_17999# a_17139_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9472 VGND a_25318_7093# a_25247_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X9473 _048_ a_16219_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X9474 VPWR a_19221_13793# _209_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X9475 tdc0.w_dly_sig[189] tdc0.w_dly_sig_n[188] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9476 VPWR a_13149_6549# _165_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X9477 VPWR tdc0.w_dly_sig_n[68] tdc0.w_dly_sig[69] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9479 tdc0.o_result[111] a_2715_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9481 VGND tdc0.w_dly_sig[126] tdc0.w_dly_sig_n[126] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9482 tdc0.o_result[100] a_4739_17179# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9483 _173_ a_14922_13897# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X9484 tdc0.w_dly_sig[127] tdc0.w_dly_sig_n[125] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9485 VPWR a_6227_3133# a_6395_3035# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9486 a_26111_12559# a_25891_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X9487 a_10202_2879# a_10034_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9488 VPWR tdc0.w_dly_sig[189] tdc0.w_dly_sig_n[189] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9490 tdc0.w_dly_sig_n[147] tdc0.w_dly_sig[147] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9491 a_24915_8359# a_25011_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9492 a_18383_8983# tdc0.o_result[58] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9493 _001_ a_18059_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X9494 VGND tdc0.w_dly_sig_n[81] tdc0.w_dly_sig[82] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9495 VGND a_23323_10651# a_23281_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9496 VGND clknet_4_3_0_clk a_10975_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9497 tdc0.w_dly_sig[180] tdc0.w_dly_sig_n[178] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9499 VGND tdc0.w_dly_sig_n[136] tdc0.w_dly_sig[138] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9500 tdc0.w_dly_sig[56] tdc0.w_dly_sig_n[55] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9502 VPWR a_10443_2197# a_10359_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9503 tdc0.w_dly_sig_n[153] tdc0.w_dly_sig[153] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9504 a_3413_5493# a_3247_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9505 a_1297_5493# a_1131_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9506 VPWR tdc0.w_dly_sig[146] tdc0.w_dly_sig_n[146] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9507 tdc0.w_dly_sig_n[80] tdc0.w_dly_sig[80] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9508 tdc0.w_dly_sig[58] tdc0.w_dly_sig_n[56] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9509 tdc0.w_dly_sig_n[156] tdc0.w_dly_sig[156] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9510 VPWR net5 a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9511 _099_ a_14379_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X9512 tdc0.o_result[144] a_13203_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9513 VPWR tdc0.w_dly_sig[152] tdc0.w_dly_sig_n[153] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9514 a_29998_3311# a_29559_3317# a_29913_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9515 VPWR a_22891_14423# _147_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X9516 _011_ net6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9517 VPWR tdc0.w_dly_sig_n[131] tdc0.w_dly_sig[132] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9518 a_15837_8181# _013_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X9520 a_15163_3543# tdc0.o_result[171] a_15397_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9521 VPWR a_11655_2045# a_11823_1947# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9522 a_19395_3543# tdc0.o_result[175] a_19629_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9523 VPWR tdc0.w_dly_sig_n[141] tdc0.w_dly_sig[142] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9524 VGND tdc0.w_dly_sig_n[150] tdc0.w_dly_sig[151] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9525 a_17967_9839# _114_ a_18217_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9526 VPWR tdc0.w_dly_sig_n[62] tdc0.w_dly_sig[64] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9527 a_17451_14191# a_16753_14197# a_17194_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9528 tdc0.w_dly_sig_n[111] tdc0.w_dly_sig[111] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9529 VPWR clknet_4_8_0_clk a_21923_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9530 VPWR a_25203_3829# a_25210_4129# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9531 a_17168_9545# _032_ a_17066_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X9532 tdc0.w_dly_sig[171] tdc0.w_dly_sig_n[169] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9533 VGND net28 a_28057_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X9534 VPWR a_29982_12671# a_29909_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9535 tdc0.w_dly_sig[106] tdc0.w_dly_sig_n[105] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9537 a_18751_2919# a_18847_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9538 VGND tdc0.w_dly_sig_n[21] tdc0.w_dly_sig[22] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9539 VGND _004_ a_23384_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X9540 VGND clknet_4_1_0_clk a_8399_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9541 tdc0.w_dly_sig_n[39] tdc0.w_dly_sig[39] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9542 VPWR tdc0.o_result[111] a_15575_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9543 a_5341_10383# tdc0.o_result[110] a_4995_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X9544 a_12762_7663# _122_ a_12448_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X9545 VGND tdc0.w_dly_sig[185] tdc0.w_dly_sig_n[185] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9547 _157_ a_13722_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X9548 tdc0.w_dly_sig_n[115] tdc0.w_dly_sig[114] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9549 a_9006_13759# a_8838_14013# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9550 VPWR a_29274_16644# a_29203_16745# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X9551 a_15370_12925# a_15097_12559# a_15285_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9552 a_6357_12015# tdc0.o_result[103] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9553 a_20145_7119# a_19598_7393# a_19798_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X9554 a_12502_9813# a_12334_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9555 a_7457_15657# a_6467_15285# a_7331_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9556 a_13551_11721# _085_ a_13633_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9557 VGND a_22167_2441# a_22174_2345# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9559 tdc0.o_result[26] a_24059_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9560 _087_ a_11159_8864# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X9561 a_15943_9295# _031_ a_16121_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9562 tdc0.w_dly_sig_n[124] tdc0.w_dly_sig[124] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9564 a_22714_703# a_22546_957# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9565 a_30515_6397# a_29651_6031# a_30258_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9566 VPWR _043_ a_12815_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9568 a_5050_8319# a_4882_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9571 VGND _058_ a_16649_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9572 a_7584_11305# a_7185_10933# a_7458_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9573 a_9424_9129# a_9025_8757# a_9298_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9574 VPWR tdc0.w_dly_sig_n[41] tdc0.w_dly_sig[43] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9575 clknet_4_14_0_clk a_26882_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9576 a_23891_7663# a_23027_7669# a_23634_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9577 VGND a_29987_11145# a_29994_11049# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9578 VGND a_14123_2197# a_14081_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9579 tdc0.w_dly_sig_n[158] tdc0.w_dly_sig[158] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9580 VGND a_16543_17063# tdc0.o_result[59] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9581 tdc0.w_dly_sig_n[189] tdc0.w_dly_sig[189] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9582 VPWR tdc0.w_dly_sig[69] tdc0.w_dly_sig_n[70] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9584 clknet_4_3_0_clk a_10506_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9585 VPWR a_21039_3133# a_21207_3035# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9586 a_9347_9661# a_8565_9295# a_9263_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9587 a_30159_5853# a_29939_5865# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X9588 VPWR a_30343_7284# net26 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9589 VGND a_21914_17732# a_21843_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X9590 VPWR tdc0.w_dly_sig[5] a_27137_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9591 a_20003_11305# a_19867_11145# a_19583_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9592 a_7263_6005# clknet_4_3_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9593 VPWR _137_ a_18309_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X9594 VGND tdc0.w_dly_sig[33] tdc0.w_dly_sig_n[33] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9595 tdc0.w_dly_sig[91] tdc0.w_dly_sig_n[90] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9596 VPWR tdc0.w_dly_sig_n[139] tdc0.w_dly_sig[140] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9597 VPWR a_9006_8319# a_8933_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9598 VPWR tdc0.w_dly_sig[76] tdc0.w_dly_sig_n[76] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9599 a_24283_2741# clknet_4_10_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9601 a_4057_2767# a_3891_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9602 VPWR tdc0.w_dly_sig_n[105] tdc0.w_dly_sig[107] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9603 VGND tdc0.w_dly_sig[11] tdc0.w_dly_sig_n[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9604 tdc0.w_dly_sig_n[107] tdc0.w_dly_sig[107] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9605 tdc0.w_dly_sig_n[153] tdc0.w_dly_sig[152] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9606 VGND tdc0.w_dly_sig[17] tdc0.w_dly_sig_n[17] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9607 tdc0.w_dly_sig[12] tdc0.w_dly_sig_n[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9608 VPWR tdc0.w_dly_sig_n[79] tdc0.w_dly_sig[81] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9609 _092_ a_7479_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X9610 VGND a_27123_5719# tdc0.o_result[17] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9611 VPWR tdc0.w_dly_sig_n[147] tdc0.w_dly_sig[149] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9612 VPWR tdc0.w_dly_sig[145] tdc0.w_dly_sig_n[146] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9613 VGND a_13997_7637# _023_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X9614 VPWR tdc0.w_dly_sig_n[111] tdc0.w_dly_sig[112] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9615 tdc0.w_dly_sig_n[157] tdc0.w_dly_sig[157] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9616 VGND tdc0.w_dly_sig[45] tdc0.w_dly_sig_n[45] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9617 tdc0.w_dly_sig_n[67] tdc0.w_dly_sig[67] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9618 a_26046_15101# a_25799_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X9619 a_6821_15279# tdc0.w_dly_sig[102] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9620 VPWR tdc0.w_dly_sig[104] tdc0.w_dly_sig_n[104] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9621 a_27413_15657# a_26859_15497# a_27066_15556# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X9622 VGND tdc0.w_dly_sig[99] tdc0.w_dly_sig_n[100] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9624 VPWR a_22771_17179# a_22687_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9625 VGND tdc0.w_dly_sig[115] tdc0.w_dly_sig_n[115] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9626 VGND tdc0.w_dly_sig_n[92] tdc0.w_dly_sig[94] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9627 VPWR tdc0.w_dly_sig[57] tdc0.w_dly_sig_n[57] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9628 a_19221_13793# _208_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9629 VPWR tdc0.w_dly_sig[139] tdc0.w_dly_sig_n[140] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9630 a_9025_8757# a_8859_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9631 VGND tdc0.w_dly_sig[148] tdc0.w_dly_sig_n[149] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9632 VGND tdc0.w_dly_sig_n[23] tdc0.w_dly_sig[24] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9633 a_4797_6031# tdc0.w_dly_sig[147] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9634 VPWR a_30591_3285# a_30507_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9635 a_25295_8181# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9636 VPWR a_21879_12711# tdc0.o_result[37] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9638 VGND a_14151_10535# _074_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X9639 a_18751_2919# a_18847_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9640 a_19693_591# a_18703_591# a_19567_957# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9641 _169_ a_12434_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9642 a_20609_11721# _029_ a_20359_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9643 a_13367_9952# _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9644 VGND tdc0.w_dly_sig_n[187] tdc0.w_dly_sig[188] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9645 tdc0.w_dly_sig_n[173] tdc0.w_dly_sig[173] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9646 a_20089_8207# _030_ a_20017_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9647 tdc0.w_dly_sig_n[49] tdc0.w_dly_sig[48] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9648 a_26111_4943# a_25891_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X9649 a_23027_5487# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X9650 VGND a_23139_16091# a_23097_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9651 a_24490_18820# a_24290_18665# a_24639_18909# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X9652 VPWR tdc0.w_dly_sig_n[163] tdc0.w_dly_sig[165] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9653 a_5767_9661# a_5069_9295# a_5510_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9654 VGND tdc0.w_dly_sig[191] tdc0.w_dly_sig_n[192] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9655 _164_ a_12723_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X9656 a_16707_3133# a_15925_2767# a_16623_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9657 VPWR a_3651_14191# a_3819_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9658 tdc0.w_dly_sig[123] tdc0.w_dly_sig_n[122] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9659 a_25410_13103# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X9660 a_10436_12559# a_10037_12559# a_10310_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9661 VGND _024_ a_14011_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X9662 tdc0.w_dly_sig_n[99] tdc0.w_dly_sig[99] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9664 a_6077_11471# tdc0.o_result[102] a_5639_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9665 VGND tdc0.w_dly_sig[150] tdc0.w_dly_sig_n[150] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9666 VGND a_9983_7387# a_9941_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9667 tdc0.w_dly_sig[93] tdc0.w_dly_sig_n[91] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9668 clknet_4_13_0_clk a_19890_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9669 a_22914_8751# a_22641_8757# a_22829_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9670 a_25226_13621# a_25026_13921# a_25375_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X9671 VGND tdc0.w_dly_sig_n[15] tdc0.w_dly_sig[17] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9672 a_4698_8751# a_4425_8757# a_4613_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9676 a_21707_17673# clknet_4_12_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9677 VGND tdc0.w_dly_sig[23] a_25849_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X9678 VGND a_19015_2223# a_19183_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9679 a_19487_11159# a_19583_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9680 a_29519_5719# a_29803_5705# a_29738_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X9681 a_19225_11721# _064_ a_18703_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9682 a_5897_3133# a_5363_2767# a_5802_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9683 VGND a_20359_3855# _051_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X9684 VPWR ui_in[6] a_17507_1143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X9686 tdc0.o_result[72] a_15963_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9687 VGND tdc0.w_dly_sig_n[126] tdc0.w_dly_sig[128] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9689 VPWR tdc0.o_result[90] a_14563_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9690 VPWR a_20499_13799# _207_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X9691 a_13641_12559# _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X9692 a_15013_5487# net2 _024_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9693 a_24013_11445# tdc0.o_result[8] a_24266_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X9694 _064_ _010_ a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9695 a_28883_13321# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9696 VPWR _009_ a_17323_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X9697 a_14729_17999# a_14563_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9698 tdc0.w_dly_sig_n[51] tdc0.w_dly_sig[51] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9699 _200_ a_13643_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X9700 VGND tdc0.w_dly_sig[134] tdc0.w_dly_sig_n[135] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9701 a_28503_13335# a_28599_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9702 a_13990_3133# a_13551_2767# a_13905_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9703 VGND tdc0.w_dly_sig_n[96] tdc0.w_dly_sig[98] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9704 VPWR a_16210_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9705 VPWR tdc0.w_dly_sig[43] tdc0.w_dly_sig_n[44] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9708 VPWR _043_ a_19947_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X9709 a_23999_18775# a_24283_18761# a_24218_18909# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X9710 VGND tdc0.w_dly_sig[41] tdc0.w_dly_sig_n[41] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R25 VPWR tt_um_hpretl_tt06_tdc_v1_15.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X9711 VGND a_17383_5095# _040_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X9712 a_19099_2223# a_18317_2229# a_19015_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9713 tdc0.w_dly_sig[25] tdc0.w_dly_sig_n[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9714 a_16679_10927# _008_ a_16857_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9716 a_19843_18543# a_18979_18549# a_19586_18517# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9717 a_14064_7093# _013_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X9718 VPWR tdc0.w_dly_sig[141] tdc0.w_dly_sig_n[142] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9719 clknet_4_7_0_clk a_11812_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9720 VPWR tdc0.w_dly_sig[182] a_22721_2601# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9721 VGND a_11655_2045# a_11823_1947# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9722 VPWR clknet_4_0_0_clk a_4443_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9723 tdc0.w_dly_sig_n[88] tdc0.w_dly_sig[88] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9724 a_19150_8207# _160_ a_19396_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X9725 tdc0.w_dly_sig[165] tdc0.w_dly_sig_n[163] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9727 tdc0.w_dly_sig_n[155] tdc0.w_dly_sig[155] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9728 tdc0.w_dly_sig_n[172] tdc0.w_dly_sig[172] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9729 a_21638_8181# a_21431_8181# a_21814_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X9730 VGND a_27491_2919# tdc0.o_result[187] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9731 a_13748_16745# a_13349_16373# a_13622_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9733 a_25870_14709# a_25663_14709# a_26046_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X9735 VGND tdc0.w_dly_sig[23] tdc0.w_dly_sig_n[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9736 VPWR a_12851_15101# a_13019_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9737 VPWR a_21223_2045# a_21391_1947# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9738 VPWR tdc0.w_dly_sig_n[165] tdc0.w_dly_sig[166] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9739 a_18751_5095# tdc0.o_result[12] a_18985_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9740 VPWR a_29331_7284# net23 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9741 a_4057_2767# a_3891_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9742 tdc0.w_dly_sig[134] tdc0.w_dly_sig_n[133] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9743 a_9853_16911# a_9687_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9744 VPWR a_7883_10927# a_8051_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9745 VGND a_4463_11739# a_4421_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9746 VPWR tdc0.w_dly_sig_n[178] tdc0.w_dly_sig[179] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9747 a_18479_6895# _001_ _064_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9748 tdc0.o_result[130] a_9431_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9749 clknet_0_clk a_16210_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9750 VPWR _017_ a_16845_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X9751 a_19304_4399# _203_ a_19202_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X9752 a_9926_9813# a_9758_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9753 a_25155_3689# a_25019_3529# a_24735_3543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9754 clknet_4_0_0_clk a_6476_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9755 a_14250_18517# a_14082_18543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9756 VGND tdc0.w_dly_sig[100] tdc0.w_dly_sig_n[101] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9757 a_19550_13897# _207_ a_19470_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X9758 VPWR a_24490_2741# a_24419_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X9759 tdc0.w_dly_sig_n[20] tdc0.w_dly_sig[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9760 VPWR a_21104_6005# clknet_4_8_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9761 a_2673_13647# a_1683_13647# a_2547_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9763 a_30515_6397# a_29817_6031# a_30258_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9764 a_3099_7663# a_2235_7669# a_2842_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9765 a_6633_15285# a_6467_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9766 clknet_4_6_0_clk a_12254_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9767 a_20709_3133# a_20175_2767# a_20614_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9768 a_29266_13103# a_29019_13481# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X9769 a_25962_4917# a_25762_5217# a_26111_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X9770 a_25283_14887# a_25379_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9772 uo_out[4] a_19225_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9773 VPWR clknet_4_3_0_clk a_8951_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9774 VPWR tdc0.w_dly_sig[123] tdc0.w_dly_sig_n[124] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9775 VGND tdc0.w_dly_sig[97] tdc0.w_dly_sig_n[97] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9777 VGND a_18751_5095# _142_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X9778 tdc0.w_dly_sig[143] tdc0.w_dly_sig_n[141] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9779 a_4237_5865# a_3247_5493# a_4111_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9780 a_30166_7637# a_29998_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9781 a_24021_14985# tdc0.o_result[47] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9782 VGND tdc0.w_dly_sig[42] tdc0.w_dly_sig_n[42] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9784 tdc0.w_dly_sig_n[132] tdc0.w_dly_sig[131] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9786 tdc0.w_dly_sig_n[145] tdc0.w_dly_sig[144] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9788 VPWR a_10506_7119# clknet_4_3_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9789 tdc0.w_dly_sig[169] tdc0.w_dly_sig_n[167] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9790 VGND clknet_0_clk a_10506_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9791 a_4498_2879# a_4330_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9792 a_2037_13103# tdc0.w_dly_sig[112] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9793 tdc0.w_dly_sig[47] tdc0.w_dly_sig_n[45] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9794 a_24731_7271# a_24827_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9795 a_10183_9839# a_9485_9845# a_9926_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9797 tdc0.w_dly_sig_n[136] tdc0.w_dly_sig[135] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9798 VGND clknet_4_12_0_clk a_18979_18549# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9799 a_13580_6575# _162_ a_13478_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X9800 a_10459_3133# a_9595_2767# a_10202_2879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9801 VPWR a_27491_2919# tdc0.o_result[187] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9802 a_14418_13103# _118_ a_14104_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X9804 VPWR clknet_4_0_0_clk a_2787_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9805 a_13809_18549# a_13643_18549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9806 VPWR tdc0.w_dly_sig[88] tdc0.w_dly_sig_n[88] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9808 a_2217_4405# a_2051_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9810 tdc0.w_dly_sig[166] tdc0.w_dly_sig_n[165] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9811 a_24735_13621# a_25026_13921# a_24977_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9812 tdc0.w_dly_sig_n[173] tdc0.w_dly_sig[172] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9813 VGND a_24653_9545# uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9814 a_21603_4007# tdc0.o_result[182] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9815 VPWR clknet_4_2_0_clk a_12171_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9816 tdc0.w_dly_sig[71] tdc0.w_dly_sig_n[70] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9817 VGND tdc0.w_dly_sig_n[21] tdc0.w_dly_sig[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9818 tdc0.o_result[91] a_14675_18517# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9819 a_20175_12809# _192_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9820 VGND tdc0.w_dly_sig[137] tdc0.w_dly_sig_n[137] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9821 a_11513_18543# tdc0.w_dly_sig[94] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9822 a_21814_8573# a_21567_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X9823 VPWR tdc0.w_dly_sig[63] tdc0.w_dly_sig_n[63] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9824 VGND a_15687_16091# a_15645_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9825 VPWR a_30683_6299# a_30599_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9826 VGND _031_ a_24488_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X9827 a_28883_12233# clknet_4_14_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9828 a_5261_10927# _027_ a_5115_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X9829 VGND tdc0.w_dly_sig[184] tdc0.w_dly_sig_n[185] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9830 _035_ a_14255_6835# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9831 VGND _031_ a_15380_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X9832 VGND a_16210_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9833 a_17415_11247# _094_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X9834 VGND a_8914_17429# a_8872_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9835 VPWR tdc0.w_dly_sig_n[59] tdc0.w_dly_sig[61] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9836 VPWR tdc0.w_dly_sig[192] a_30449_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9837 _139_ a_12723_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X9838 tdc0.w_dly_sig_n[154] tdc0.w_dly_sig[153] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9839 a_30258_6143# a_30090_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9840 VGND a_6550_12559# clknet_4_4_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9841 a_6191_12015# _023_ a_6369_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9842 tdc0.w_dly_sig[134] tdc0.w_dly_sig_n[132] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9843 VPWR a_24283_18761# a_24290_18665# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9844 a_23385_8207# tdc0.o_result[22] a_23303_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9845 a_4571_17277# a_3873_16911# a_4314_17023# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9846 a_28078_2741# a_27871_2741# a_28254_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X9847 VPWR tdc0.w_dly_sig[165] tdc0.w_dly_sig_n[165] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9848 a_29761_5487# a_29423_5719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X9849 a_8753_15823# tdc0.w_dly_sig[100] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9850 VPWR tdc0.w_dly_sig_n[136] tdc0.w_dly_sig[137] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9851 a_15146_9839# _083_ a_14897_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X9852 a_8638_16341# a_8470_16367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9853 a_10402_11837# a_9963_11471# a_10317_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9854 tdc0.w_dly_sig_n[86] tdc0.w_dly_sig[86] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9855 VPWR tdc0.w_dly_sig[44] tdc0.w_dly_sig_n[45] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9856 VGND tdc0.w_dly_sig[74] tdc0.w_dly_sig_n[74] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9857 tdc0.w_dly_sig[185] tdc0.w_dly_sig_n[184] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9858 a_8377_12393# a_7387_12021# a_8251_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9859 VGND a_27526_12292# a_27455_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X9863 VGND clknet_4_3_0_clk a_10975_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9864 VPWR a_26514_6575# clknet_4_11_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9865 tdc0.o_result[89] a_14215_16341# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9866 VPWR tdc0.o_result[149] a_12723_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9867 a_27087_9129# a_26951_8969# a_26667_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9868 tdc0.w_dly_sig_n[163] tdc0.w_dly_sig[163] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9869 a_8470_16367# a_8197_16373# a_8385_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9870 a_16193_8725# tdc0.o_result[155] a_16446_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X9872 _001_ a_18059_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9873 a_2750_6549# a_2582_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9874 tdc0.w_dly_sig[145] tdc0.w_dly_sig_n[144] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9876 VPWR _067_ a_24131_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9877 VPWR a_20074_6005# a_20003_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X9878 a_22891_6807# a_22987_6807# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9880 VGND tdc0.w_dly_sig[163] tdc0.w_dly_sig_n[164] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9881 tdc0.w_dly_sig_n[146] tdc0.w_dly_sig[145] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9882 tdc0.w_dly_sig[149] tdc0.w_dly_sig_n[147] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9883 _033_ a_17691_6281# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.157 ps=1.32 w=1 l=0.15
X9884 a_29090_13380# a_28883_13321# a_29266_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X9885 VPWR tdc0.w_dly_sig[147] tdc0.w_dly_sig_n[148] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9887 a_19307_7093# a_19598_7393# a_19549_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9889 VPWR a_28883_13321# a_28890_13225# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9890 VGND tdc0.w_dly_sig[180] tdc0.w_dly_sig_n[180] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9891 VGND tdc0.w_dly_sig_n[14] tdc0.w_dly_sig[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9892 a_23947_12335# tdc0.o_result[5] a_24469_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X9893 VGND net6 a_18045_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X9894 tdc0.w_dly_sig[36] tdc0.w_dly_sig_n[35] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9895 VGND clknet_4_1_0_clk a_7847_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9896 VGND a_7499_15253# a_7457_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9897 VPWR a_12115_1135# a_12283_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9898 net5 a_17507_1143# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X9899 a_29019_13481# a_28883_13321# a_28599_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9900 a_24823_4007# a_24919_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9901 a_24504_11471# _014_ a_24013_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X9902 VGND _142_ a_18046_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X9903 VPWR net2 a_17923_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X9904 a_23386_17732# a_23186_17577# a_23535_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X9905 _057_ a_16311_3424# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X9906 _079_ a_14195_3424# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X9907 clknet_0_clk a_16210_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9908 VPWR tdc0.w_dly_sig[103] tdc0.w_dly_sig_n[103] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9909 VPWR _092_ a_17415_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9911 VGND tdc0.w_dly_sig_n[3] tdc0.w_dly_sig[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9912 VGND tdc0.w_dly_sig[7] tdc0.w_dly_sig_n[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9913 VPWR tdc0.w_dly_sig_n[68] tdc0.w_dly_sig[70] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9914 VPWR tdc0.w_dly_sig[39] tdc0.w_dly_sig_n[40] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9915 a_16566_957# a_16127_591# a_16481_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9916 VPWR tdc0.w_dly_sig[177] tdc0.w_dly_sig_n[178] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9917 VGND tdc0.w_dly_sig_n[92] tdc0.w_dly_sig[93] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9918 a_15603_16189# a_14821_15823# a_15519_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9919 tdc0.o_result[31] a_22679_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9920 VPWR a_4130_4373# a_4057_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9921 VGND tdc0.w_dly_sig[20] tdc0.w_dly_sig_n[21] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9922 VGND tdc0.w_dly_sig_n[137] tdc0.w_dly_sig[138] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9923 VPWR a_12007_6549# a_11923_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9924 a_22729_16911# a_21739_16911# a_22603_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9925 VPWR tdc0.w_dly_sig_n[158] tdc0.w_dly_sig[159] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9926 VGND a_21223_2045# a_21391_1947# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9928 a_4563_4221# a_3781_3855# a_4479_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9929 a_23110_5487# tdc0.o_result[31] a_23027_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9930 tdc0.w_dly_sig[49] tdc0.w_dly_sig_n[48] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9931 VGND a_26755_7895# tdc0.o_result[18] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9932 a_10252_16911# a_9853_16911# a_10126_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9933 VGND a_2547_14013# a_2715_13915# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9934 VPWR a_4866_8725# a_4793_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9935 VGND a_19867_11145# a_19874_11049# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9936 VPWR tdc0.w_dly_sig[189] tdc0.w_dly_sig_n[190] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9937 VPWR tdc0.w_dly_sig_n[72] tdc0.w_dly_sig[74] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9939 VPWR tdc0.w_dly_sig[96] tdc0.w_dly_sig_n[96] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9940 VPWR tdc0.w_dly_sig_n[29] tdc0.w_dly_sig[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9942 VPWR tdc0.w_dly_sig_n[82] tdc0.w_dly_sig[84] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9943 tdc0.w_dly_sig[86] tdc0.w_dly_sig_n[85] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9944 a_11230_2045# a_10957_1679# a_11145_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9945 tdc0.w_dly_sig_n[94] tdc0.w_dly_sig[93] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9946 VPWR tdc0.w_dly_sig_n[44] tdc0.w_dly_sig[46] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9947 tdc0.w_dly_sig[120] tdc0.w_dly_sig_n[119] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9948 tdc0.w_dly_sig_n[28] tdc0.w_dly_sig[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9949 a_10037_12559# a_9871_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9951 tdc0.w_dly_sig[130] tdc0.w_dly_sig_n[128] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9952 a_17937_10927# _110_ a_17665_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9953 tdc0.w_dly_sig[22] tdc0.w_dly_sig_n[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9954 tdc0.w_dly_sig_n[138] tdc0.w_dly_sig[137] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9955 VGND tdc0.w_dly_sig[30] a_21985_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X9956 a_27319_12233# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9957 VGND a_14675_18517# a_14633_18921# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9958 tdc0.w_dly_sig[92] tdc0.w_dly_sig_n[91] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9959 a_14131_16367# a_13349_16373# a_14047_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9960 VGND a_10443_2197# a_10401_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9961 a_16661_957# a_16127_591# a_16566_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9963 a_8895_16367# a_8197_16373# a_8638_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9964 a_24125_14511# tdc0.o_result[53] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X9965 tdc0.w_dly_sig_n[188] tdc0.w_dly_sig[187] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9966 a_8378_2223# a_7939_2229# a_8293_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9967 VGND a_15731_7271# _006_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X9968 tdc0.w_dly_sig[76] tdc0.w_dly_sig_n[74] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9969 VPWR tdc0.w_dly_sig_n[77] tdc0.w_dly_sig[79] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9970 a_25651_8207# a_25431_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X9971 a_13809_17461# a_13643_17461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9972 a_25799_14735# a_25670_15009# a_25379_14709# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X9973 VPWR tdc0.w_dly_sig_n[9] tdc0.w_dly_sig[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9974 tdc0.w_dly_sig_n[81] tdc0.w_dly_sig[80] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9975 VPWR a_6476_6549# clknet_4_0_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9976 VGND tdc0.w_dly_sig[38] tdc0.w_dly_sig_n[39] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9977 VGND _005_ a_16127_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X9978 VPWR clknet_4_6_0_clk a_9871_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9979 VGND _205_ a_19255_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X9980 a_28254_3133# a_28007_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X9981 tdc0.w_dly_sig[146] tdc0.w_dly_sig_n[144] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9983 VPWR tdc0.w_dly_sig_n[64] tdc0.w_dly_sig[65] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9984 a_17937_10927# _064_ a_17415_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9985 clknet_4_8_0_clk a_21104_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9986 VPWR _035_ a_16679_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9987 a_2490_4399# a_2051_4405# a_2405_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9988 _150_ a_18059_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X9989 a_7561_11721# _091_ a_7479_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9990 a_29025_16367# a_28687_16599# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X9991 tdc0.o_result[43] a_30407_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9992 tdc0.o_result[172] a_17619_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9993 tdc0.w_dly_sig_n[129] tdc0.w_dly_sig[128] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9994 a_4882_8573# a_4609_8207# a_4797_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9995 VGND _138_ a_13354_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X9996 a_12594_15935# a_12426_16189# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9998 tdc0.o_result[142] a_11639_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9999 tdc0.w_dly_sig[27] tdc0.w_dly_sig_n[26] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10000 tdc0.w_dly_sig[135] tdc0.w_dly_sig_n[134] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10001 a_26667_8181# a_26958_8481# a_26909_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X10002 VPWR tdc0.w_dly_sig_n[126] tdc0.w_dly_sig[127] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10003 VGND tdc0.w_dly_sig_n[168] tdc0.w_dly_sig[170] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10004 tdc0.w_dly_sig[35] tdc0.w_dly_sig_n[34] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10005 _100_ a_14563_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X10006 a_12115_3133# a_11251_2767# a_11858_2879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10007 VGND tdc0.w_dly_sig_n[171] tdc0.w_dly_sig[172] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10008 net3 a_16219_1143# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X10009 VGND net3 _024_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10010 a_14415_3133# a_13717_2767# a_14158_2879# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10011 VPWR tdc0.w_dly_sig_n[142] tdc0.w_dly_sig[143] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10012 a_27137_11471# a_26583_11445# a_26790_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X10013 tdc0.w_dly_sig[103] tdc0.w_dly_sig_n[102] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10014 VPWR _085_ a_8573_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X10015 VGND tdc0.w_dly_sig_n[156] tdc0.w_dly_sig[158] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10016 VGND a_15170_18111# a_15128_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10017 a_7166_14165# a_6998_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10018 tdc0.w_dly_sig[78] tdc0.w_dly_sig_n[76] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10019 a_5491_15101# a_4793_14735# a_5234_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10020 _065_ a_16713_8235# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X10021 VGND tdc0.w_dly_sig[55] tdc0.w_dly_sig_n[56] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10022 tdc0.w_dly_sig[87] tdc0.w_dly_sig_n[85] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10023 a_26583_11445# clknet_4_14_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10024 tdc0.w_dly_sig[34] tdc0.w_dly_sig_n[32] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10025 a_26995_15657# a_26859_15497# a_26575_15511# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X10026 VPWR tdc0.w_dly_sig[83] tdc0.w_dly_sig_n[84] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10027 VPWR clknet_4_1_0_clk a_2143_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10028 a_26903_16911# a_26774_17185# a_26483_16885# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X10029 VGND a_25755_4917# a_25762_5217# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10030 VGND a_25428_7637# clknet_4_10_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R26 tt_um_hpretl_tt06_tdc_v1_19.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10031 VGND clknet_4_4_0_clk a_1315_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10032 VGND _151_ a_23947_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10033 a_2033_9845# a_1867_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10034 tdc0.w_dly_sig[136] tdc0.w_dly_sig_n[135] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10035 VPWR a_3267_7637# a_3183_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10036 VGND tdc0.w_dly_sig_n[12] tdc0.w_dly_sig[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10038 a_9577_2229# a_9411_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10039 a_22886_4943# _060_ a_22796_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X10041 tdc0.w_dly_sig[109] tdc0.w_dly_sig_n[107] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10042 a_17023_5487# net6 a_16665_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10043 tdc0.w_dly_sig_n[29] tdc0.w_dly_sig[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10045 VGND a_30166_8725# a_30124_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10046 VGND clknet_4_8_0_clk a_16127_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10047 tdc0.w_dly_sig[109] tdc0.w_dly_sig_n[108] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10049 a_4793_8751# a_4259_8757# a_4698_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10050 a_14563_9545# _089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X10051 VPWR _039_ a_17048_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X10052 a_6177_5487# tdc0.w_dly_sig[146] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10053 VPWR a_28883_12233# a_28890_12137# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10054 tdc0.w_dly_sig_n[20] tdc0.w_dly_sig[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10055 tdc0.w_dly_sig[140] tdc0.w_dly_sig_n[138] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10057 VPWR a_30423_7663# a_30591_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10058 tdc0.w_dly_sig[68] tdc0.w_dly_sig_n[67] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10059 a_3777_14569# a_2787_14197# a_3651_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10060 a_22856_10383# a_22457_10383# a_22730_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10062 VPWR tdc0.w_dly_sig_n[154] tdc0.w_dly_sig[156] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10063 a_17075_957# a_16293_591# a_16991_957# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10064 VPWR a_15101_7637# _047_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X10065 tdc0.w_dly_sig_n[55] tdc0.w_dly_sig[54] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10066 a_20798_2045# a_20525_1679# a_20713_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10067 a_22777_3855# _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10070 VPWR a_3651_3311# a_3819_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10071 a_15511_18365# a_14729_17999# a_15427_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10072 VPWR tdc0.w_dly_sig[47] tdc0.w_dly_sig_n[47] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10073 VGND tdc0.w_dly_sig[74] tdc0.w_dly_sig_n[75] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10074 _030_ a_17323_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X10075 tdc0.w_dly_sig_n[190] tdc0.w_dly_sig[190] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10076 clknet_4_5_0_clk a_7378_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10078 VGND a_24915_8983# _186_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X10079 VPWR tdc0.w_dly_sig_n[112] tdc0.w_dly_sig[114] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10080 VPWR tdc0.w_dly_sig_n[36] tdc0.w_dly_sig[37] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10081 uo_out[2] a_17937_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10082 a_24131_9295# _064_ a_24653_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10083 VGND tdc0.w_dly_sig_n[124] tdc0.w_dly_sig[126] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10084 tdc0.w_dly_sig_n[32] tdc0.w_dly_sig[32] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10086 VPWR _005_ a_14887_4631# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X10087 VGND a_7442_2879# a_7400_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10088 VGND tdc0.w_dly_sig[24] a_24837_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X10089 tdc0.w_dly_sig[130] tdc0.w_dly_sig_n[129] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10090 VPWR a_10627_3035# a_10543_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10091 a_18037_13423# tdc0.o_result[40] a_17599_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10092 VPWR net3 a_16665_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10093 VPWR a_1995_5487# a_2163_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10094 tdc0.w_dly_sig[45] tdc0.w_dly_sig_n[44] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10095 VGND tdc0.w_dly_sig_n[42] tdc0.w_dly_sig[44] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10096 a_14441_3855# _007_ a_14369_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10097 VPWR a_6982_16341# a_6909_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10099 VGND tdc0.w_dly_sig[61] tdc0.w_dly_sig_n[62] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10100 VGND _054_ a_24009_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10102 a_26514_6575# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10103 VGND a_21787_3543# _103_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X10105 VPWR a_5307_8573# a_5475_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10106 tdc0.o_result[9] a_30591_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10107 a_22362_15279# a_21923_15285# a_22277_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10108 a_8504_2601# a_8105_2229# a_8378_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10110 VGND tdc0.w_dly_sig_n[190] tdc0.w_dly_sig[191] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10111 a_23239_10749# a_22457_10383# a_23155_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10112 a_25502_8181# a_25302_8481# a_25651_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X10113 a_14361_10933# a_14195_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10114 a_19557_6941# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10115 VPWR tdc0.w_dly_sig_n[15] tdc0.w_dly_sig[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10116 VGND tdc0.w_dly_sig[65] tdc0.w_dly_sig_n[65] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10120 VPWR tdc0.w_dly_sig[7] a_29437_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X10121 a_21985_8207# a_21438_8481# a_21638_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X10122 VGND a_14675_17429# a_14633_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10124 VGND a_26479_15511# tdc0.o_result[47] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10125 VGND tdc0.w_dly_sig_n[157] tdc0.w_dly_sig[158] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10126 a_25962_15797# a_25762_16097# a_26111_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X10127 a_16941_2223# tdc0.w_dly_sig[173] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10128 VPWR _019_ a_16713_8235# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X10129 a_2616_4777# a_2217_4405# a_2490_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10130 a_26479_15511# a_26575_15511# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X10131 a_4755_3133# a_3891_2767# a_4498_2879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10132 VGND a_8327_4373# a_8285_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10133 a_12618_7983# tdc0.o_result[115] a_12537_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X10135 a_4606_7485# a_4167_7119# a_4521_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10136 _138_ a_11711_13216# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X10137 VPWR a_11398_1791# a_11325_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10138 VGND a_17937_10927# uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10139 tdc0.w_dly_sig_n[135] tdc0.w_dly_sig[135] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10140 a_10183_9839# a_9319_9845# a_9926_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10141 tdc0.w_dly_sig_n[68] tdc0.w_dly_sig[68] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10142 tdc0.w_dly_sig_n[70] tdc0.w_dly_sig[69] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10143 VPWR a_25226_3588# a_25155_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X10144 a_11414_7663# a_11141_7669# a_11329_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10145 a_8565_9295# a_8399_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10146 VGND a_25778_1653# a_25707_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X10147 VGND a_29982_9813# a_29940_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10148 VPWR tdc0.o_result[22] a_23303_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10149 VGND tdc0.w_dly_sig_n[101] tdc0.w_dly_sig[102] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10150 a_14461_7119# tdc0.o_result[113] a_14379_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10152 VPWR a_17435_17429# a_17351_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10153 a_7599_10749# a_6817_10383# a_7515_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10154 VPWR tdc0.w_dly_sig_n[67] tdc0.w_dly_sig[69] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10155 tdc0.w_dly_sig[107] tdc0.w_dly_sig_n[105] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10156 a_11313_9117# _025_ a_11241_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10157 a_20258_10116# a_20058_9961# a_20407_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X10158 VGND tdc0.w_dly_sig_n[76] tdc0.w_dly_sig[77] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10159 a_12778_5461# a_12610_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10160 VPWR tdc0.w_dly_sig[60] tdc0.w_dly_sig_n[60] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10161 tdc0.o_result[69] a_17251_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10162 a_2037_12559# tdc0.w_dly_sig[108] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10163 tdc0.w_dly_sig_n[95] tdc0.w_dly_sig[95] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10164 tdc0.w_dly_sig_n[15] tdc0.w_dly_sig[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10165 VGND clknet_4_3_0_clk a_8951_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10166 tdc0.w_dly_sig_n[13] tdc0.w_dly_sig[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10167 tdc0.w_dly_sig[81] tdc0.w_dly_sig_n[79] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10168 tdc0.w_dly_sig[186] tdc0.w_dly_sig_n[184] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10169 tdc0.w_dly_sig_n[170] tdc0.w_dly_sig[169] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10170 a_30423_7663# a_29559_7669# a_30166_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10172 tdc0.w_dly_sig_n[45] tdc0.w_dly_sig[45] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10173 VGND a_30423_3311# a_30591_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10174 VPWR a_30010_5764# a_29939_5865# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X10175 a_29725_7669# a_29559_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10176 a_23171_11159# a_23455_11145# a_23390_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X10177 a_16986_9545# _036_ a_16737_9441# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X10178 a_27547_13481# a_27418_13225# a_27127_13335# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X10179 VGND tdc0.w_dly_sig[30] tdc0.w_dly_sig_n[31] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10180 VPWR a_26951_8181# a_26958_8481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10181 a_8197_16373# a_8031_16373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10182 VGND a_24191_1353# a_24198_1257# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10184 tdc0.w_dly_sig_n[57] tdc0.w_dly_sig[57] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10185 a_29725_14197# a_29559_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10186 VGND tdc0.w_dly_sig_n[146] tdc0.w_dly_sig[148] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10187 tdc0.w_dly_sig_n[150] tdc0.w_dly_sig[149] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10188 tdc0.w_dly_sig[150] tdc0.w_dly_sig_n[149] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10189 VGND clknet_4_13_0_clk a_16403_17461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10190 a_27873_12393# a_27326_12137# a_27526_12292# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X10191 tdc0.w_dly_sig_n[150] tdc0.w_dly_sig[150] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10192 tdc0.w_dly_sig[124] tdc0.w_dly_sig_n[123] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10193 tdc0.w_dly_sig_n[183] tdc0.w_dly_sig[182] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10194 a_23999_15797# a_24290_16097# a_24241_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X10195 VPWR _010_ a_24170_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10196 tdc0.w_dly_sig[163] tdc0.w_dly_sig_n[161] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10197 tdc0.w_dly_sig[65] tdc0.w_dly_sig_n[63] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10198 a_1880_11305# a_1481_10933# a_1754_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10199 a_18222_16367# a_17783_16373# a_18137_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10200 tdc0.o_result[158] a_7591_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10201 tdc0.w_dly_sig[18] tdc0.w_dly_sig_n[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10202 VGND a_20945_13675# _055_ VGND sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X10203 a_3735_3311# a_2953_3317# a_3651_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10204 a_17967_10159# _130_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10205 a_25288_10357# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X10206 VGND a_26951_8969# a_26958_8873# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10207 a_16547_4373# _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X10208 tdc0.o_result[124] a_9431_13915# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10209 VPWR a_27526_12292# a_27455_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X10210 a_22672_15823# a_22273_15823# a_22546_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10211 a_3686_5487# a_3413_5493# a_3601_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10213 a_25713_12925# a_25375_12711# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X10214 tdc0.w_dly_sig[132] tdc0.w_dly_sig_n[130] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10215 a_6503_4221# a_5805_3855# a_6246_3967# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10216 tdc0.w_dly_sig_n[36] tdc0.w_dly_sig[36] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10217 a_21642_17821# a_21327_17687# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X10218 a_16490_15823# a_16175_15975# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X10220 VPWR tdc0.w_dly_sig_n[176] tdc0.w_dly_sig[178] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10222 VGND tdc0.w_dly_sig[94] tdc0.w_dly_sig_n[95] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10223 VGND a_8419_11989# a_8377_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10224 a_18489_9839# _130_ a_18217_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10226 tdc0.w_dly_sig[99] tdc0.w_dly_sig_n[98] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10227 VGND tdc0.w_dly_sig_n[4] tdc0.w_dly_sig[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10228 tdc0.w_dly_sig_n[164] tdc0.w_dly_sig[164] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10229 VPWR clknet_4_1_0_clk a_4259_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10230 VGND tdc0.w_dly_sig[41] tdc0.w_dly_sig_n[42] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10231 a_30347_10357# ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10232 VPWR tdc0.w_dly_sig[67] tdc0.w_dly_sig_n[68] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10233 a_24954_13647# a_24639_13799# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X10234 VPWR tdc0.w_dly_sig[40] tdc0.w_dly_sig_n[41] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10235 a_29437_12393# a_28883_12233# a_29090_12292# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X10236 VPWR clknet_4_9_0_clk a_21279_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10237 VGND a_4314_7637# a_4272_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10238 a_18703_11471# _064_ a_19225_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10239 VPWR a_24915_8359# tdc0.o_result[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10240 VGND tdc0.w_dly_sig_n[125] tdc0.w_dly_sig[126] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10241 VGND a_19395_6807# _045_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X10242 clknet_4_5_0_clk a_7378_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10243 VPWR a_10551_17277# a_10719_17179# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10244 a_11325_2045# a_10791_1679# a_11230_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10245 a_7350_7231# a_7182_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10246 tdc0.w_dly_sig[128] tdc0.w_dly_sig_n[126] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10247 VPWR tdc0.w_dly_sig[118] tdc0.w_dly_sig_n[119] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10248 a_28425_2767# a_27878_3041# a_28078_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X10249 VGND tdc0.w_dly_sig[103] tdc0.w_dly_sig_n[104] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10250 tdc0.w_dly_sig_n[77] tdc0.w_dly_sig[76] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10251 a_12525_5487# tdc0.w_dly_sig[145] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10252 VPWR a_23903_18775# tdc0.o_result[53] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10254 a_17477_16911# a_16930_17185# a_17130_16885# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X10255 tdc0.w_dly_sig_n[54] tdc0.w_dly_sig[54] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10256 VPWR tdc0.o_result[147] a_12539_6688# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10257 a_20543_9295# _069_ a_20721_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X10258 VGND tdc0.w_dly_sig_n[54] tdc0.w_dly_sig[56] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10260 a_13641_9295# _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X10261 tdc0.w_dly_sig_n[80] tdc0.w_dly_sig[79] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10262 VGND _171_ a_5639_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10263 a_3778_10927# a_3505_10933# a_3693_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10264 VGND tdc0.w_dly_sig_n[140] tdc0.w_dly_sig[141] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10265 VGND clknet_4_4_0_clk a_3339_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10266 a_5342_9661# a_4903_9295# a_5257_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10268 tdc0.w_dly_sig[112] tdc0.w_dly_sig_n[110] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10269 a_4732_7119# a_4333_7119# a_4606_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10270 tdc0.w_dly_sig_n[44] tdc0.w_dly_sig[43] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10271 VPWR _040_ a_14287_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X10272 a_2953_14197# a_2787_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10274 a_19947_4007# tdc0.o_result[190] a_20181_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10275 a_17023_5487# a_16495_5487# _011_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10276 VPWR a_27158_9028# a_27087_9129# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X10277 VGND tdc0.w_dly_sig_n[51] tdc0.w_dly_sig[53] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10279 a_13905_2767# tdc0.w_dly_sig[172] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10280 VGND a_10903_12827# a_10861_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10281 tdc0.w_dly_sig_n[148] tdc0.w_dly_sig[148] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10282 a_19395_7895# tdc0.o_result[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10283 VGND a_7883_10927# a_8051_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10285 a_10409_14735# tdc0.w_dly_sig[84] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10286 a_26719_11471# a_26590_11745# a_26299_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X10287 VPWR a_12283_3035# a_12199_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10288 tdc0.w_dly_sig[183] tdc0.w_dly_sig_n[182] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10289 tdc0.w_dly_sig_n[129] tdc0.w_dly_sig[129] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10290 VPWR a_21380_14165# clknet_4_12_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10291 a_19337_12809# _209_ a_19255_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
R27 VPWR tt_um_hpretl_tt06_tdc_v1_12.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10292 clknet_0_clk a_16210_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10293 a_24731_14423# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X10294 VGND tdc0.w_dly_sig[37] tdc0.w_dly_sig_n[38] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10295 VPWR tdc0.w_dly_sig_n[63] tdc0.w_dly_sig[65] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10296 a_17498_12015# tdc0.o_result[107] a_17415_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10297 tdc0.w_dly_sig[156] tdc0.w_dly_sig_n[155] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10298 tdc0.w_dly_sig_n[16] tdc0.w_dly_sig[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10299 VGND a_14897_9813# _084_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X10300 VPWR a_25571_1653# a_25578_1953# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10301 a_23855_13647# _003_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10302 VPWR clknet_4_2_0_clk a_11619_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10303 clknet_0_clk a_16210_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10304 a_14461_6031# tdc0.o_result[145] a_14379_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10305 a_8201_7663# tdc0.w_dly_sig[132] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10306 VGND a_9431_16091# a_9389_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10307 a_11540_14569# a_11141_14197# a_11414_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10308 a_27093_7663# a_26755_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X10309 VGND tdc0.w_dly_sig[166] tdc0.w_dly_sig_n[166] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10310 VPWR a_11858_1109# a_11785_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10312 VGND tdc0.w_dly_sig_n[168] tdc0.w_dly_sig[169] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10313 VGND clknet_4_7_0_clk a_9687_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10314 a_15333_4737# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X10315 tdc0.w_dly_sig[178] tdc0.w_dly_sig_n[176] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10316 VPWR clknet_0_clk a_21104_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10317 VPWR tdc0.w_dly_sig_n[132] tdc0.w_dly_sig[134] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10318 VGND clknet_4_2_0_clk a_11251_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10319 a_26299_7093# a_26590_7393# a_26541_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X10320 a_25713_5309# a_25375_5095# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X10321 a_17565_8725# _095_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X10322 VPWR a_13019_11739# a_12935_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10325 a_4149_4221# a_3615_3855# a_4054_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10326 VGND tdc0.w_dly_sig[40] tdc0.w_dly_sig_n[40] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10327 VPWR a_15963_12827# a_15879_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10328 a_2037_11471# tdc0.w_dly_sig[109] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10329 clknet_4_6_0_clk a_12254_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10330 a_3996_11471# a_3597_11471# a_3870_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10331 VGND a_24398_1412# a_24327_1513# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X10332 a_8887_2223# a_8105_2229# a_8803_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10333 VGND tdc0.w_dly_sig[178] tdc0.w_dly_sig_n[178] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10334 a_1113_6031# a_947_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10335 _029_ a_17599_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X10336 uo_out[6] a_19777_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10337 VGND tdc0.w_dly_sig_n[181] tdc0.w_dly_sig[182] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10338 VGND tdc0.w_dly_sig[161] tdc0.w_dly_sig_n[161] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10339 a_17773_14735# tdc0.o_result[125] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X10340 VGND tdc0.w_dly_sig[125] tdc0.w_dly_sig_n[125] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10341 a_6913_3311# tdc0.w_dly_sig[159] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10342 _107_ a_21923_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X10343 VPWR tdc0.w_dly_sig_n[90] tdc0.w_dly_sig[92] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10344 VGND tdc0.w_dly_sig[57] tdc0.w_dly_sig_n[58] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10345 VGND a_9063_16341# a_9021_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10346 tdc0.w_dly_sig_n[183] tdc0.w_dly_sig[183] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10347 _126_ a_23303_3424# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X10348 a_27710_5764# a_27510_5609# a_27859_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X10349 _076_ a_14064_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X10350 VGND tdc0.w_dly_sig[71] tdc0.w_dly_sig_n[72] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10351 tdc0.w_dly_sig[162] tdc0.w_dly_sig_n[161] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10352 VGND _056_ a_16465_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10353 VPWR a_19211_7271# tdc0.o_result[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10354 a_16481_18543# tdc0.w_dly_sig[57] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10355 VPWR clknet_4_5_0_clk a_6467_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10356 VPWR a_11260_5461# clknet_4_2_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10357 VPWR tdc0.o_result[109] a_13580_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10358 a_15354_17023# a_15186_17277# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10360 a_2999_4399# a_2217_4405# a_2915_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10361 VPWR a_25283_14887# tdc0.o_result[41] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10362 _011_ net6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X10363 a_17949_16373# a_17783_16373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10364 a_10037_12559# a_9871_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10365 _038_ a_16733_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10366 a_14897_9813# _083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X10367 VGND clknet_0_clk a_21380_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X10368 a_25288_10357# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X10369 tdc0.w_dly_sig[8] tdc0.w_dly_sig_n[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10370 VGND tdc0.o_result[48] a_24504_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X10371 a_25339_3855# a_25203_3829# a_24919_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X10372 VPWR a_20966_1791# a_20893_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10373 a_13997_7637# _022_ a_14243_8001# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X10374 a_17887_12809# tdc0.o_result[59] a_17685_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10375 a_4379_11837# a_3597_11471# a_4295_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10376 tdc0.w_dly_sig_n[107] tdc0.w_dly_sig[106] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10377 VPWR tdc0.w_dly_sig_n[4] tdc0.w_dly_sig[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10378 VGND tdc0.w_dly_sig_n[62] tdc0.w_dly_sig[63] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10379 VGND a_24469_12015# uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10380 VPWR tdc0.w_dly_sig_n[78] tdc0.w_dly_sig[80] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10381 a_5993_3855# tdc0.w_dly_sig[158] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10382 a_29515_4631# a_29611_4631# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X10383 _060_ a_16127_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X10384 a_2750_6549# a_2582_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10385 VGND clknet_4_6_0_clk a_9871_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10386 a_27001_4221# a_26663_4007# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X10388 VGND tdc0.w_dly_sig_n[57] tdc0.w_dly_sig[58] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10389 VGND tdc0.w_dly_sig[121] tdc0.w_dly_sig_n[122] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10390 VPWR _005_ a_16127_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X10391 VPWR clknet_4_12_0_clk a_21739_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10393 VPWR tdc0.w_dly_sig[28] a_20145_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X10394 tdc0.w_dly_sig[116] tdc0.w_dly_sig_n[115] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10395 VPWR a_9723_8751# a_9891_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10396 a_8661_17455# tdc0.w_dly_sig[97] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10397 a_27369_13103# a_27031_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X10399 a_3735_14191# a_2953_14197# a_3651_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10401 a_30365_12559# a_29375_12559# a_30239_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10402 tdc0.w_dly_sig_n[118] tdc0.w_dly_sig[117] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10403 VPWR tdc0.w_dly_sig[171] tdc0.w_dly_sig_n[171] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10404 tdc0.w_dly_sig_n[31] tdc0.w_dly_sig[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10405 tdc0.w_dly_sig[106] tdc0.w_dly_sig_n[104] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10406 VPWR tdc0.w_dly_sig[172] tdc0.w_dly_sig_n[172] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10407 _157_ a_13722_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X10408 tdc0.w_dly_sig[33] tdc0.w_dly_sig_n[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10410 VGND a_7626_10901# a_7584_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10411 VPWR tdc0.o_result[105] a_15023_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10412 a_14766_8751# _116_ a_14686_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X10413 a_23947_14191# _014_ a_24125_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X10414 a_7189_2767# tdc0.w_dly_sig[160] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10415 a_24639_4943# a_24419_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X10416 VGND clknet_4_3_0_clk a_10975_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10417 a_8838_8573# a_8399_8207# a_8753_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10419 a_19767_10071# a_20058_9961# a_20009_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X10420 VGND a_20499_5719# _196_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X10422 VPWR tdc0.w_dly_sig_n[125] tdc0.w_dly_sig[127] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10423 VPWR _192_ a_20175_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10424 a_25678_8573# a_25431_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X10426 VPWR tdc0.w_dly_sig[28] tdc0.w_dly_sig_n[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10427 VPWR a_4923_3035# a_4839_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10428 a_16488_6935# a_16301_6575# a_16401_6691# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X10429 VPWR a_24469_12015# uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10430 a_5468_9295# a_5069_9295# a_5342_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10431 a_19255_12335# _172_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10432 tdc0.w_dly_sig_n[151] tdc0.w_dly_sig[151] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10433 VGND a_4774_7231# a_4732_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10434 a_12521_15101# a_11987_14735# a_12426_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10435 VGND a_25226_13621# a_25155_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X10436 VGND a_16734_703# a_16692_591# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10437 VPWR tdc0.w_dly_sig_n[127] tdc0.w_dly_sig[128] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10438 tdc0.w_dly_sig[3] tdc0.w_dly_sig_n[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10439 a_27710_5764# a_27503_5705# a_27886_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X10441 _044_ a_13459_3424# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X10442 VGND a_12254_13103# clknet_4_6_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10443 tdc0.o_result[30] a_23507_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10444 VPWR _068_ a_17773_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X10445 VPWR a_10351_9813# a_10267_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10446 VPWR tdc0.w_dly_sig_n[6] tdc0.w_dly_sig[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10447 tdc0.w_dly_sig[61] tdc0.w_dly_sig_n[59] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10448 VGND a_3819_14165# a_3777_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10449 _187_ a_23855_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X10450 VGND tdc0.w_dly_sig[179] tdc0.w_dly_sig_n[180] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10451 a_11785_1135# a_11251_1141# a_11690_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10452 VPWR a_11582_7637# a_11509_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10453 a_15885_7369# net4 a_15801_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10454 VGND tdc0.w_dly_sig_n[163] tdc0.w_dly_sig[164] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10455 VGND tdc0.w_dly_sig_n[58] tdc0.w_dly_sig[60] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10456 a_20661_13647# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10458 VGND tdc0.w_dly_sig[137] a_7817_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X10459 a_24254_8751# _188_ a_24005_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X10460 a_12594_14847# a_12426_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10461 a_8385_3311# tdc0.w_dly_sig[161] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10462 VGND a_15595_2197# a_15553_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10463 tdc0.w_dly_sig_n[181] tdc0.w_dly_sig[181] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10464 VGND tdc0.w_dly_sig[1] tdc0.w_dly_sig_n[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10465 VPWR tdc0.o_result[113] a_14379_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10466 _167_ a_11711_4512# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X10467 VGND clknet_4_0_0_clk a_6835_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10468 VPWR a_26571_8359# tdc0.o_result[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10469 a_19671_10071# a_19767_10071# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10470 tdc0.w_dly_sig_n[45] tdc0.w_dly_sig[44] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10471 VPWR a_14047_16367# a_14215_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10472 a_15185_11305# a_14195_10933# a_15059_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10473 a_9941_7119# a_8951_7119# a_9815_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10474 a_6725_14197# a_6559_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10475 VPWR _010_ a_19119_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X10476 VPWR a_25375_5095# tdc0.o_result[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10478 a_30423_8751# a_29725_8757# a_30166_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10479 VPWR a_30591_7637# a_30507_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10480 VGND a_14047_16367# a_14215_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10481 VGND tdc0.w_dly_sig[99] tdc0.w_dly_sig_n[99] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10482 a_4613_12015# tdc0.w_dly_sig[120] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10483 a_9761_2767# a_9595_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10484 a_20175_12809# _194_ a_20425_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10485 a_10819_12925# a_10037_12559# a_10735_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10486 VGND tdc0.w_dly_sig_n[19] tdc0.w_dly_sig[20] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10487 a_26215_9269# clknet_4_11_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10488 a_10310_14013# a_9871_13647# a_10225_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10489 tdc0.w_dly_sig_n[22] tdc0.w_dly_sig[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10490 VPWR clknet_4_2_0_clk a_11251_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10491 VPWR tdc0.w_dly_sig_n[26] tdc0.w_dly_sig[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10492 a_14182_10159# _033_ a_14428_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X10493 a_14520_13103# _119_ a_14418_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X10494 VPWR tdc0.w_dly_sig_n[24] tdc0.w_dly_sig[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10495 tdc0.w_dly_sig[41] tdc0.w_dly_sig_n[40] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10496 VPWR tdc0.w_dly_sig_n[134] tdc0.w_dly_sig[135] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10498 _182_ a_14287_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X10499 a_20893_2045# a_20359_1679# a_20798_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10500 _072_ a_14045_12353# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X10502 VPWR a_2163_7387# a_2079_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10503 a_10862_8573# a_10423_8207# a_10777_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10504 VPWR tdc0.w_dly_sig_n[73] tdc0.w_dly_sig[75] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10505 VGND clknet_4_2_0_clk a_9411_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10506 VGND tdc0.w_dly_sig[113] tdc0.w_dly_sig_n[114] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10508 VPWR tdc0.w_dly_sig_n[85] tdc0.w_dly_sig[87] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10509 a_17349_13647# _034_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10510 VGND _187_ a_24005_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X10511 a_25467_11471# a_25247_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X10512 VPWR tdc0.w_dly_sig_n[89] tdc0.w_dly_sig[90] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10513 a_16366_2879# a_16198_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10514 tdc0.o_result[165] a_12651_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10515 VGND tdc0.w_dly_sig_n[147] tdc0.w_dly_sig[148] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10516 VPWR a_26583_7093# a_26590_7393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10517 VGND tdc0.w_dly_sig_n[140] tdc0.w_dly_sig[142] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10518 a_20881_11721# _064_ a_20359_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10519 VPWR tdc0.w_dly_sig[51] tdc0.w_dly_sig_n[52] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10520 VGND tdc0.w_dly_sig_n[186] tdc0.w_dly_sig[188] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10521 VPWR a_3854_5461# a_3781_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10522 VPWR a_1738_5461# a_1665_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10523 VGND _040_ a_15545_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10524 VGND tdc0.w_dly_sig[51] a_27321_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X10525 tdc0.w_dly_sig_n[7] tdc0.w_dly_sig[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10526 a_4605_3855# a_3615_3855# a_4479_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10527 a_19557_8029# _011_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10529 a_15519_16189# a_14655_15823# a_15262_15935# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10530 VGND a_15262_15935# a_15220_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10531 VGND tdc0.w_dly_sig[68] tdc0.w_dly_sig_n[69] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10532 VGND tdc0.w_dly_sig[2] a_26769_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X10533 a_8573_10927# tdc0.o_result[79] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X10534 VPWR a_19338_2741# a_19267_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X10535 a_20499_5719# tdc0.o_result[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10536 VPWR tdc0.w_dly_sig[29] tdc0.w_dly_sig_n[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10537 VPWR tdc0.w_dly_sig_n[116] tdc0.w_dly_sig[118] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R28 uio_oe[2] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10538 VGND clknet_0_clk a_11260_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X10539 VPWR tdc0.w_dly_sig_n[38] tdc0.w_dly_sig[39] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10540 a_19375_13441# _011_ a_19289_13441# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X10541 a_12977_15823# a_11987_15823# a_12851_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10542 tdc0.w_dly_sig_n[152] tdc0.w_dly_sig[152] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10543 a_17703_6895# net6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10544 tdc0.w_dly_sig[74] tdc0.w_dly_sig_n[72] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10545 a_12969_2767# _025_ a_12897_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10546 VPWR tdc0.o_result[154] a_15391_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10547 a_29019_12393# a_28890_12137# a_28599_12247# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X10548 tdc0.w_dly_sig_n[109] tdc0.w_dly_sig[108] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10549 a_16739_7895# net5 a_16913_8001# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X10550 VGND tdc0.w_dly_sig[32] tdc0.w_dly_sig_n[33] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10551 tdc0.w_dly_sig[84] tdc0.w_dly_sig_n[82] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10552 a_15189_16189# a_14655_15823# a_15094_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10553 VGND tdc0.w_dly_sig[180] tdc0.w_dly_sig_n[181] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10554 a_30549_15657# a_29559_15285# a_30423_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10556 clknet_4_14_0_clk a_26882_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10557 tdc0.w_dly_sig[113] tdc0.w_dly_sig_n[111] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10558 a_27886_5487# a_27639_5865# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X10560 a_16734_703# a_16566_957# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10561 VGND _180_ a_13722_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X10562 a_21423_17687# a_21707_17673# a_21642_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X10564 a_19145_18549# a_18979_18549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10565 a_23423_8751# a_22641_8757# a_23339_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10566 a_5207_8751# a_4425_8757# a_5123_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10567 a_14047_16367# a_13183_16373# a_13790_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10568 VGND tdc0.w_dly_sig[153] tdc0.w_dly_sig_n[154] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10569 VPWR a_12594_14847# a_12521_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10572 a_24490_4917# a_24290_5217# a_24639_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X10573 a_13552_8457# tdc0.o_result[117] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X10574 a_8964_8207# a_8565_8207# a_8838_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10576 VPWR clknet_4_5_0_clk a_6559_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10577 VGND tdc0.w_dly_sig[41] a_27965_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X10578 VGND a_7442_14847# a_7400_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10579 a_19855_7895# tdc0.o_result[19] a_20089_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10580 VPWR a_22799_17687# tdc0.o_result[52] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10581 tdc0.w_dly_sig_n[39] tdc0.w_dly_sig[38] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10582 a_4061_7663# tdc0.w_dly_sig[118] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10583 VGND tdc0.w_dly_sig_n[179] tdc0.w_dly_sig[180] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10584 VGND tdc0.w_dly_sig[61] tdc0.w_dly_sig_n[61] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10585 VGND a_5510_9407# a_5468_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10586 VGND tdc0.w_dly_sig_n[42] tdc0.w_dly_sig[43] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10587 a_9485_9845# a_9319_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10588 a_17415_11247# _064_ a_17937_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10589 VPWR a_7423_14191# a_7591_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10590 a_3007_6575# a_2309_6581# a_2750_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10591 a_10620_14735# a_10221_14735# a_10494_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10592 VGND a_30239_12925# a_30407_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10593 a_21837_3855# _060_ a_21765_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10594 a_17209_14735# a_16219_14735# a_17083_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10595 VPWR tdc0.w_dly_sig[24] tdc0.w_dly_sig_n[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10596 tdc0.w_dly_sig_n[10] tdc0.w_dly_sig[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10597 VGND a_16713_8235# _065_ VGND sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X10598 VGND a_29423_5719# tdc0.o_result[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10599 VPWR tdc0.w_dly_sig_n[138] tdc0.w_dly_sig[139] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10600 VPWR a_5031_15279# a_5199_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10601 VGND tdc0.w_dly_sig_n[64] tdc0.w_dly_sig[66] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10602 a_23700_9839# _004_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X10603 VPWR tdc0.w_dly_sig_n[94] tdc0.w_dly_sig[96] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10604 VGND tdc0.w_dly_sig_n[103] tdc0.w_dly_sig[105] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10605 a_20499_5719# tdc0.o_result[23] a_20733_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10606 VGND a_26951_8181# a_26958_8481# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10607 VPWR tdc0.w_dly_sig_n[46] tdc0.w_dly_sig[48] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10608 VPWR tdc0.w_dly_sig[6] tdc0.w_dly_sig_n[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10609 VPWR tdc0.w_dly_sig_n[94] tdc0.w_dly_sig[95] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10610 VGND a_10719_17179# a_10677_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10611 VGND tdc0.w_dly_sig_n[175] tdc0.w_dly_sig[176] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10612 tdc0.w_dly_sig[127] tdc0.w_dly_sig_n[126] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10614 a_4314_17023# a_4146_17277# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10615 VGND a_22530_15253# a_22488_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10616 tdc0.w_dly_sig_n[191] tdc0.w_dly_sig[190] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10617 a_27271_8041# a_27135_7881# a_26851_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X10618 VGND tdc0.w_dly_sig[184] tdc0.w_dly_sig_n[184] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10619 VGND a_20211_15279# a_20379_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10620 VPWR clknet_4_0_0_clk a_6835_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10621 a_25891_4943# a_25755_4917# a_25471_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X10622 a_17593_8029# a_17323_7663# a_17503_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X10623 _089_ a_12526_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X10624 VPWR tdc0.w_dly_sig[8] tdc0.w_dly_sig_n[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10625 tdc0.o_result[179] a_23139_859# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10626 a_7783_15101# a_7001_14735# a_7699_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10627 tdc0.w_dly_sig_n[58] tdc0.w_dly_sig[58] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10628 a_30124_15657# a_29725_15285# a_29998_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10629 tdc0.w_dly_sig_n[69] tdc0.w_dly_sig[69] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10630 VGND a_20039_5719# _136_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X10631 VPWR clknet_4_4_0_clk a_9319_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10633 a_19881_10633# tdc0.o_result[32] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X10634 a_30423_7663# a_29725_7669# a_30166_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10635 VGND a_21591_15101# a_21759_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10636 a_9389_13647# a_8399_13647# a_9263_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10637 a_9761_2767# a_9595_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10638 tdc0.w_dly_sig[10] tdc0.w_dly_sig_n[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10639 VGND a_13019_15003# a_12977_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10640 a_3781_5487# a_3247_5493# a_3686_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10641 a_1665_5487# a_1131_5493# a_1570_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10642 VPWR a_16547_7093# _022_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X10643 a_7561_11721# _023_ a_7645_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10644 VGND tdc0.w_dly_sig[188] tdc0.w_dly_sig_n[189] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10645 _152_ a_23947_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X10646 a_16842_17455# a_16569_17461# a_16757_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10647 a_19928_5193# _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X10648 a_11973_2223# tdc0.w_dly_sig[166] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10649 _104_ a_17047_3424# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X10650 a_2290_13077# a_2122_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10651 a_6262_4399# a_5989_4405# a_6177_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10652 a_10988_8207# a_10589_8207# a_10862_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10653 tdc0.w_dly_sig[57] tdc0.w_dly_sig_n[55] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10655 clknet_4_9_0_clk a_22852_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10656 a_7921_12015# a_7387_12021# a_7826_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10657 a_16761_10383# tdc0.o_result[80] a_16679_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10658 VPWR a_15575_591# net2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10659 VGND tdc0.w_dly_sig_n[95] tdc0.w_dly_sig[97] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10660 clknet_4_8_0_clk a_21104_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10661 a_5905_10927# _131_ a_5823_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10662 tdc0.w_dly_sig[192] tdc0.w_dly_sig_n[191] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10663 VPWR a_21603_4007# _183_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10664 VPWR clk a_16210_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10665 a_22395_12559# a_22266_12833# a_21975_12533# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X10666 VPWR tdc0.w_dly_sig_n[97] tdc0.w_dly_sig[99] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10667 tdc0.w_dly_sig[189] tdc0.w_dly_sig_n[187] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10668 VPWR a_18935_3543# _061_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10669 a_9558_7231# a_9390_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10670 a_24344_8457# _106_ a_24242_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X10671 VGND tdc0.w_dly_sig[35] tdc0.w_dly_sig_n[35] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10672 VPWR tdc0.w_dly_sig[186] tdc0.w_dly_sig_n[187] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10673 a_13354_13423# _139_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X10674 a_14158_2879# a_13990_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10675 VGND tdc0.w_dly_sig_n[159] tdc0.w_dly_sig[161] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10676 VPWR tdc0.w_dly_sig[43] tdc0.w_dly_sig_n[43] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10677 tdc0.w_dly_sig[15] tdc0.w_dly_sig_n[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10678 a_15427_18365# a_14563_17999# a_15170_18111# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10680 tdc0.w_dly_sig_n[47] tdc0.w_dly_sig[47] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10681 tdc0.w_dly_sig_n[75] tdc0.w_dly_sig[74] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10682 a_26851_7895# a_27135_7881# a_27070_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X10684 a_24490_15797# a_24290_16097# a_24639_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X10685 tdc0.w_dly_sig[167] tdc0.w_dly_sig_n[166] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10686 tdc0.o_result[140] a_12007_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10687 clknet_4_3_0_clk a_10506_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10688 VPWR tdc0.w_dly_sig[128] tdc0.w_dly_sig_n[129] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10689 VPWR tdc0.w_dly_sig[146] tdc0.w_dly_sig_n[147] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10690 a_16999_4917# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0767 ps=0.785 w=0.42 l=0.15
X10691 tdc0.o_result[74] a_13019_11739# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10692 a_10911_11837# a_10129_11471# a_10827_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10693 tdc0.w_dly_sig_n[165] tdc0.w_dly_sig[165] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10694 VPWR _072_ a_14012_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X10695 VGND _147_ a_22809_13793# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X10696 VPWR tdc0.w_dly_sig_n[87] tdc0.w_dly_sig[89] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10697 tdc0.w_dly_sig_n[156] tdc0.w_dly_sig[155] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10698 a_15097_18365# a_14563_17999# a_15002_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10699 a_13184_13103# tdc0.o_result[140] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X10700 VGND a_27710_5764# a_27639_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X10701 a_27137_11471# a_26590_11745# a_26790_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X10702 VPWR a_7166_3285# a_7093_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10703 VPWR _050_ a_24363_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X10704 a_20211_15279# a_19347_15285# a_19954_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10705 VGND tdc0.w_dly_sig[46] tdc0.w_dly_sig_n[47] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10706 VPWR tdc0.w_dly_sig_n[5] tdc0.w_dly_sig[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10707 a_24837_4943# a_24283_4917# a_24490_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X10708 a_11965_6031# a_10975_6031# a_11839_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10709 VGND tdc0.w_dly_sig[116] tdc0.w_dly_sig_n[117] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10710 VGND a_18390_16341# a_18348_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10711 a_12058_2223# a_11785_2229# a_11973_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10713 a_2815_9839# a_2033_9845# a_2731_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10714 VPWR tdc0.w_dly_sig[10] tdc0.w_dly_sig_n[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10715 VGND _019_ a_18823_6059# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X10716 a_9389_9295# a_8399_9295# a_9263_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10717 a_1849_13109# a_1683_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10718 tdc0.w_dly_sig_n[114] tdc0.w_dly_sig[113] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10719 VPWR clknet_4_6_0_clk a_14195_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10720 a_14974_11471# _058_ a_14884_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X10721 a_3689_4405# a_3523_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10722 a_25849_8207# a_25302_8481# a_25502_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X10723 tdc0.o_result[162] a_10627_3035# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10724 a_15170_18111# a_15002_18365# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10725 tdc0.w_dly_sig[159] tdc0.w_dly_sig_n[158] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10726 VGND a_25571_1653# a_25578_1953# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10727 tdc0.w_dly_sig_n[167] tdc0.w_dly_sig[166] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10729 a_22093_16911# tdc0.w_dly_sig[62] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10730 VPWR tdc0.w_dly_sig[38] a_22813_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X10731 a_4222_3967# a_4054_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10732 a_16923_16885# clknet_4_12_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10734 VGND tdc0.w_dly_sig[3] tdc0.w_dly_sig_n[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10735 VPWR a_3083_4373# a_2999_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10737 a_18413_591# a_18236_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X10738 tdc0.w_dly_sig_n[192] tdc0.w_dly_sig[192] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10739 tdc0.w_dly_sig_n[164] tdc0.w_dly_sig[163] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10740 VGND tdc0.w_dly_sig[120] tdc0.w_dly_sig_n[121] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10741 uo_out[7] a_20697_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10742 VPWR tdc0.w_dly_sig[161] tdc0.w_dly_sig_n[162] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10743 VPWR a_16179_7637# _002_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X10744 VGND tdc0.w_dly_sig_n[112] tdc0.w_dly_sig[113] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10745 tdc0.w_dly_sig[30] tdc0.w_dly_sig_n[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10746 VPWR _072_ a_6357_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X10747 a_25690_15823# a_25375_15975# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X10748 clknet_4_15_0_clk a_25410_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10749 tdc0.w_dly_sig_n[133] tdc0.w_dly_sig[133] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10750 a_15565_10383# tdc0.o_result[120] a_15483_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10751 tdc0.w_dly_sig_n[180] tdc0.w_dly_sig[180] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10752 a_11398_1791# a_11230_2045# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10753 VPWR net6 a_18196_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10754 VPWR a_14255_6835# _035_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X10755 tdc0.w_dly_sig[21] tdc0.w_dly_sig_n[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10756 VPWR a_24059_7637# a_23975_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10757 VPWR a_24639_3543# tdc0.o_result[186] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10758 VGND _028_ a_17599_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10759 VPWR tdc0.w_dly_sig[95] tdc0.w_dly_sig_n[96] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10760 a_20848_4399# _017_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X10761 a_25375_8983# tdc0.o_result[10] a_25609_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10762 a_6430_13077# a_6262_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10763 a_14633_17833# a_13643_17461# a_14507_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10765 a_25019_13621# clknet_4_15_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10767 a_16881_17277# a_16543_17063# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X10768 clknet_4_13_0_clk a_19890_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10769 a_29940_12559# a_29541_12559# a_29814_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10770 a_13445_2223# tdc0.w_dly_sig[170] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10771 tdc0.w_dly_sig[125] tdc0.w_dly_sig_n[123] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10773 VGND a_19289_13441# _017_ VGND sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X10775 a_16797_3855# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10776 tdc0.o_result[43] a_30407_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10777 tdc0.w_dly_sig[69] tdc0.w_dly_sig_n[67] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10778 a_26759_4631# a_27050_4521# a_27001_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X10779 a_23999_15797# a_24283_15797# a_24218_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X10780 tdc0.w_dly_sig[28] tdc0.w_dly_sig_n[26] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10781 VPWR tdc0.w_dly_sig[121] tdc0.w_dly_sig_n[121] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10782 VPWR clknet_4_6_0_clk a_9963_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10783 VPWR a_12007_14165# a_11923_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10784 a_6262_13103# a_5989_13109# a_6177_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10785 a_7619_6031# a_7399_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X10786 a_11417_1141# a_11251_1141# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10788 VGND tdc0.w_dly_sig_n[111] tdc0.w_dly_sig[113] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10789 VPWR tdc0.w_dly_sig[138] tdc0.w_dly_sig_n[139] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10790 tdc0.w_dly_sig[72] tdc0.w_dly_sig_n[71] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10791 clknet_4_12_0_clk a_21380_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10792 VPWR a_7994_11989# a_7921_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10793 VPWR tdc0.w_dly_sig_n[189] tdc0.w_dly_sig[191] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10794 a_23907_1367# a_24198_1257# a_24149_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X10795 VPWR tdc0.w_dly_sig_n[139] tdc0.w_dly_sig[141] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10796 VPWR a_26203_7271# tdc0.o_result[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R29 VGND uio_out[7] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10797 VPWR tdc0.w_dly_sig[55] tdc0.w_dly_sig_n[55] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10798 VGND tdc0.w_dly_sig[5] a_27137_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X10799 _125_ a_12618_7983# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X10800 a_16543_17063# a_16639_16885# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X10801 a_5234_14847# a_5066_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10802 tdc0.o_result[150] a_3175_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10803 VPWR tdc0.w_dly_sig[32] tdc0.w_dly_sig_n[32] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10804 a_11471_5309# a_10773_4943# a_11214_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10805 tdc0.w_dly_sig[170] tdc0.w_dly_sig_n[168] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10806 a_19395_3543# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X10807 net1 a_30347_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10808 tdc0.w_dly_sig[67] tdc0.w_dly_sig_n[65] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10809 a_17577_14569# a_16587_14197# a_17451_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10810 a_20782_2879# a_20614_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10811 a_17967_10159# _114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X10812 VPWR a_6687_5487# a_6855_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10813 VPWR clknet_4_1_0_clk a_1131_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10814 a_13722_9295# _180_ a_13968_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X10815 tdc0.w_dly_sig[158] tdc0.w_dly_sig_n[156] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10816 VGND tdc0.w_dly_sig[51] tdc0.w_dly_sig_n[51] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10817 VGND a_4130_4373# a_4088_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10818 a_16311_3424# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10819 VPWR _050_ a_23075_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X10820 tdc0.w_dly_sig_n[124] tdc0.w_dly_sig[123] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10821 a_22457_10383# a_22291_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10823 a_19413_9545# _181_ a_19341_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X10824 VPWR tdc0.w_dly_sig_n[177] tdc0.w_dly_sig[178] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10825 VPWR a_16999_4917# a_16733_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0609 ps=0.71 w=0.42 l=0.15
X10826 VGND _130_ a_17967_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X10827 VPWR tdc0.o_result[84] a_11711_13216# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10828 VGND a_7166_14165# a_7124_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10829 VPWR tdc0.w_dly_sig_n[169] tdc0.w_dly_sig[170] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10830 tdc0.o_result[146] a_5475_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10831 tdc0.w_dly_sig[181] tdc0.w_dly_sig_n[180] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10832 a_7093_3311# a_6559_3317# a_6998_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10833 VGND a_30194_11445# a_30123_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X10834 tdc0.w_dly_sig_n[159] tdc0.w_dly_sig[159] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10836 VPWR a_1979_6299# a_1895_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10837 a_12341_14735# tdc0.w_dly_sig[72] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10838 tdc0.w_dly_sig_n[127] tdc0.w_dly_sig[126] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10839 a_19255_12335# tdc0.o_result[6] a_19777_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X10840 a_26790_7093# a_26583_7093# a_26966_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X10841 VPWR clknet_4_4_0_clk a_1867_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10842 VPWR tdc0.w_dly_sig_n[162] tdc0.w_dly_sig[164] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10844 VGND _072_ a_6077_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X10845 VPWR a_17139_8759# _054_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X10847 a_1554_6143# a_1386_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10848 VPWR tdc0.w_dly_sig_n[83] tdc0.w_dly_sig[84] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10849 tdc0.w_dly_sig_n[120] tdc0.w_dly_sig[119] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10850 a_6353_2767# a_5363_2767# a_6227_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10852 a_26571_9295# a_26351_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X10853 a_18703_14985# _065_ a_18785_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10854 tdc0.w_dly_sig[5] tdc0.w_dly_sig_n[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10855 VGND a_30347_10357# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10856 a_16645_11989# _057_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X10857 tdc0.w_dly_sig_n[41] tdc0.w_dly_sig[40] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10858 a_22790_5193# tdc0.o_result[28] a_22633_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10859 a_19741_5853# _011_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10860 VGND a_23271_6793# a_23278_6697# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10861 VGND tdc0.w_dly_sig_n[150] tdc0.w_dly_sig[152] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10862 a_16994_13103# _048_ a_16680_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X10863 a_10827_11837# a_10129_11471# a_10570_11583# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10864 a_16587_11721# _062_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X10865 VPWR tdc0.w_dly_sig[4] tdc0.w_dly_sig_n[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10866 a_6817_10383# a_6651_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10867 VPWR _075_ a_14813_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X10868 VPWR tdc0.w_dly_sig[78] tdc0.w_dly_sig_n[78] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10869 VGND a_24183_15511# _067_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X10871 a_19697_14197# a_19531_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10872 VGND _043_ a_13613_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10873 tdc0.w_dly_sig_n[104] tdc0.w_dly_sig[103] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10874 VPWR tdc0.w_dly_sig_n[18] tdc0.w_dly_sig[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10875 VGND tdc0.w_dly_sig_n[121] tdc0.w_dly_sig[123] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10876 VPWR a_21707_11145# a_21714_11049# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10877 a_11329_6031# tdc0.w_dly_sig[141] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10878 a_13061_7119# _024_ a_12989_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10879 a_18317_16367# a_17783_16373# a_18222_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10880 a_9850_2223# a_9411_2229# a_9765_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10881 tdc0.w_dly_sig[39] tdc0.w_dly_sig_n[37] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10882 VPWR a_24443_16367# a_24611_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10883 VGND _163_ a_13149_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X10885 tdc0.w_dly_sig_n[105] tdc0.w_dly_sig[105] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10886 a_16219_13647# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10887 a_11793_13469# tdc0.o_result[84] a_11711_13216# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10888 VPWR a_26571_8983# tdc0.o_result[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10889 VPWR a_21104_6005# clknet_4_8_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10890 a_13357_8029# tdc0.o_result[133] a_13275_7776# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10891 VGND a_24443_16367# a_24611_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10892 VPWR clknet_4_5_0_clk a_2787_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10893 a_16210_9839# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10894 tdc0.w_dly_sig[53] tdc0.w_dly_sig_n[51] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10895 VGND tdc0.w_dly_sig[11] tdc0.w_dly_sig_n[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10896 a_3962_4399# a_3523_4405# a_3877_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10897 VGND tdc0.w_dly_sig[66] tdc0.w_dly_sig_n[66] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10899 _088_ a_11251_4512# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X10900 a_5257_9295# tdc0.w_dly_sig[121] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10901 a_20733_13647# _003_ a_20661_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10902 VGND a_11812_13621# clknet_4_7_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10903 a_6078_4221# a_5639_3855# a_5993_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10904 a_26663_4631# a_26759_4631# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X10905 a_6550_12559# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X10906 a_23811_11293# a_23591_11305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X10907 VGND a_12115_1135# a_12283_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10909 tdc0.w_dly_sig[178] tdc0.w_dly_sig_n[177] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10910 VGND tdc0.w_dly_sig[62] tdc0.w_dly_sig_n[62] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10911 a_16762_15797# a_16562_16097# a_16911_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X10912 VPWR a_17251_15003# a_17167_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10914 tdc0.o_result[121] a_5659_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10915 a_11582_6143# a_11414_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10916 tdc0.w_dly_sig[16] tdc0.w_dly_sig_n[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10917 VPWR _060_ a_23903_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X10918 _039_ a_15333_4737# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X10919 a_5391_8573# a_4609_8207# a_5307_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10920 VPWR tdc0.w_dly_sig_n[40] tdc0.w_dly_sig[42] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10923 a_27035_10071# a_27326_9961# a_27277_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X10924 a_23903_18775# a_23999_18775# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10925 VPWR tdc0.w_dly_sig[64] tdc0.w_dly_sig_n[64] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10926 a_7470_6005# a_7270_6305# a_7619_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X10927 _148_ a_22291_14304# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X10928 a_18029_3855# _038_ a_17957_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10929 tdc0.w_dly_sig_n[59] tdc0.w_dly_sig[58] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10930 VGND a_30591_15253# a_30549_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10931 a_23838_10927# a_23591_11305# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X10932 VPWR tdc0.w_dly_sig[170] tdc0.w_dly_sig_n[171] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10933 VGND a_26583_7093# a_26590_7393# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10934 VPWR a_6476_7637# clknet_4_1_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10935 VGND tdc0.w_dly_sig[174] tdc0.w_dly_sig_n[175] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10936 a_29830_4765# a_29515_4631# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X10937 VGND a_23139_13077# a_23097_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10938 a_19797_10633# _008_ a_19881_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10939 a_7323_16367# a_6541_16373# a_7239_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10940 VGND _196_ a_20325_5089# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X10941 a_11030_8319# a_10862_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10942 a_8964_15823# a_8565_15823# a_8838_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10943 VPWR tdc0.w_dly_sig[72] tdc0.w_dly_sig_n[72] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10944 a_25431_8207# a_25302_8481# a_25011_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X10945 tdc0.w_dly_sig_n[174] tdc0.w_dly_sig[173] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10946 a_3260_15657# a_2861_15285# a_3134_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10947 VPWR tdc0.w_dly_sig[46] tdc0.w_dly_sig_n[46] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10949 VGND tdc0.w_dly_sig[109] tdc0.w_dly_sig_n[110] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10950 VPWR tdc0.w_dly_sig[35] a_22261_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X10951 a_6771_5487# a_5989_5493# a_6687_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10952 VPWR a_26767_16885# a_26774_17185# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10953 a_3778_10927# a_3339_10933# a_3693_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10954 VGND a_4647_4123# a_4605_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10955 VPWR tdc0.w_dly_sig[183] tdc0.w_dly_sig_n[184] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10956 VGND tdc0.w_dly_sig[23] tdc0.w_dly_sig_n[24] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10957 a_8491_10927# _027_ a_8573_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X10958 VPWR tdc0.w_dly_sig_n[164] tdc0.w_dly_sig[166] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10959 VPWR a_6430_4373# a_6357_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10960 VGND a_19777_12015# uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10961 VGND tdc0.w_dly_sig_n[174] tdc0.w_dly_sig[176] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10962 a_2122_12925# a_1683_12559# a_2037_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10963 VGND clknet_4_1_0_clk a_4903_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10964 VGND tdc0.w_dly_sig[107] tdc0.w_dly_sig_n[108] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10966 VPWR _132_ a_18703_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10967 a_21165_2767# a_20175_2767# a_21039_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10968 tdc0.o_result[184] a_22955_3035# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10969 VGND a_4866_8725# a_4824_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10970 tdc0.w_dly_sig[92] tdc0.w_dly_sig_n[90] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10971 a_12199_1135# a_11417_1141# a_12115_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10972 VPWR _030_ a_18751_5095# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X10973 a_25621_15101# a_25283_14887# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X10974 a_16481_591# tdc0.w_dly_sig[171] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10975 tdc0.o_result[137] a_12007_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10976 a_17773_14985# tdc0.o_result[69] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X10977 tdc0.w_dly_sig[43] tdc0.w_dly_sig_n[42] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10978 VPWR a_9431_13915# a_9347_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10979 VPWR a_4739_7637# a_4655_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10980 a_16569_17461# a_16403_17461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10981 VGND clknet_4_5_0_clk a_5823_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10982 VGND a_22955_3035# a_22913_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10983 _116_ a_12539_3424# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X10984 a_24915_8983# tdc0.o_result[14] a_25149_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10985 VGND tdc0.w_dly_sig_n[10] tdc0.w_dly_sig[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10986 a_22273_15823# a_22107_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10988 tdc0.w_dly_sig[83] tdc0.w_dly_sig_n[82] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10989 tdc0.w_dly_sig_n[40] tdc0.w_dly_sig[39] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10990 tdc0.w_dly_sig[111] tdc0.w_dly_sig_n[110] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10991 a_3413_5493# a_3247_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10992 a_1297_5493# a_1131_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10994 VGND _022_ a_14131_12353# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X10995 _035_ a_14255_6835# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X10997 a_24580_9071# tdc0.o_result[30] a_24005_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X10998 a_24443_16367# a_23579_16373# a_24186_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10999 VGND tdc0.w_dly_sig[75] tdc0.w_dly_sig_n[76] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11000 _120_ a_14103_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X11001 a_19867_6005# clknet_4_9_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11002 tdc0.w_dly_sig[63] tdc0.w_dly_sig_n[62] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11003 VPWR tdc0.o_result[70] a_18151_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11005 a_20756_5193# _195_ a_20654_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X11006 a_24419_18921# a_24290_18665# a_23999_18775# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X11007 tdc0.o_result[172] a_17619_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11008 a_20848_4399# _182_ a_20746_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X11009 a_7074_15253# a_6906_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X11011 VPWR tdc0.w_dly_sig[52] tdc0.w_dly_sig_n[52] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11012 tdc0.w_dly_sig[46] tdc0.w_dly_sig_n[44] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11013 a_22642_12925# a_22395_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X11014 a_24666_18543# a_24419_18921# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X11015 a_26422_9269# a_26222_9569# a_26571_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X11016 tdc0.o_result[73] a_11915_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11017 a_21307_2045# a_20525_1679# a_21223_2045# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11018 tdc0.w_dly_sig[133] tdc0.w_dly_sig_n[132] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11019 a_12621_6941# tdc0.o_result[147] a_12539_6688# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11020 a_23413_10927# a_23075_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X11021 a_24639_18909# a_24419_18921# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X11022 tdc0.w_dly_sig[146] tdc0.w_dly_sig_n[145] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11023 VGND a_19867_6005# a_19874_6305# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11024 VGND a_11915_9563# a_11873_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11025 VPWR tdc0.o_result[11] a_17415_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X11026 VPWR a_12226_2197# a_12153_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11027 VGND tdc0.w_dly_sig[141] tdc0.w_dly_sig_n[141] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11028 a_14379_6031# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11030 VGND tdc0.w_dly_sig_n[58] tdc0.w_dly_sig[59] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11031 a_24327_1513# a_24198_1257# a_23907_1367# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X11032 VPWR clknet_0_clk a_26514_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11033 tdc0.w_dly_sig[64] tdc0.w_dly_sig_n[63] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11034 a_20175_12559# _064_ a_20697_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11035 a_4425_12021# a_4259_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11036 a_16753_14197# a_16587_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11037 a_16769_13423# _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X11039 VGND tdc0.w_dly_sig_n[33] tdc0.w_dly_sig[35] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11040 a_9976_2601# a_9577_2229# a_9850_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11041 tdc0.w_dly_sig[179] tdc0.w_dly_sig_n[178] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11043 a_14805_6549# _077_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11044 VGND a_12254_13103# clknet_4_6_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11045 tdc0.w_dly_sig_n[59] tdc0.w_dly_sig[59] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11046 a_14415_3133# a_13551_2767# a_14158_2879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11047 a_5905_10927# _023_ a_5989_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11048 VPWR tdc0.w_dly_sig_n[53] tdc0.w_dly_sig[54] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11049 tdc0.w_dly_sig[73] tdc0.w_dly_sig_n[71] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11050 VGND tdc0.w_dly_sig_n[145] tdc0.w_dly_sig[147] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11051 uo_out[5] a_24469_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11052 VGND _202_ a_19058_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X11053 a_12999_4399# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X11054 a_8753_8207# tdc0.w_dly_sig[131] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11055 tdc0.o_result[70] a_17619_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11056 tdc0.w_dly_sig[174] tdc0.w_dly_sig_n[172] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11057 a_26483_16885# a_26774_17185# a_26725_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X11058 a_12610_5487# a_12171_5493# a_12525_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11059 a_11582_7637# a_11414_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
R30 VGND uio_oe[0] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11061 VGND tdc0.w_dly_sig_n[22] tdc0.w_dly_sig[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11062 a_3777_3689# a_2787_3317# a_3651_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11063 a_18821_8029# _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X11064 a_5970_2879# a_5802_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11065 a_6204_3855# a_5805_3855# a_6078_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11066 a_29913_15279# tdc0.w_dly_sig[46] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11067 a_7741_12015# tdc0.w_dly_sig[128] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11069 VPWR a_27123_5719# tdc0.o_result[17] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11070 a_13968_8457# _156_ a_13866_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X11071 tdc0.w_dly_sig[100] tdc0.w_dly_sig_n[98] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11072 VPWR tdc0.w_dly_sig_n[101] tdc0.w_dly_sig[103] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11073 tdc0.w_dly_sig[29] tdc0.w_dly_sig_n[28] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11074 a_15347_8001# _011_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X11075 VGND tdc0.w_dly_sig_n[185] tdc0.w_dly_sig[187] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11076 VGND _040_ a_20017_4737# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X11077 tdc0.w_dly_sig_n[1] tdc0.w_dly_sig[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11078 a_30549_3689# a_29559_3317# a_30423_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11080 VGND a_30423_7663# a_30591_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11081 a_16301_13647# tdc0.o_result[96] a_16219_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11082 a_19281_5853# _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X11083 VGND a_21879_12711# tdc0.o_result[37] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11084 a_7817_6031# a_7263_6005# a_7470_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X11085 tdc0.w_dly_sig[135] tdc0.w_dly_sig_n[133] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11086 VGND tdc0.w_dly_sig_n[95] tdc0.w_dly_sig[96] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11088 VGND a_27250_4676# a_27179_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X11089 a_3597_11471# a_3431_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11090 VGND a_17746_18111# a_17704_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11092 tdc0.w_dly_sig_n[127] tdc0.w_dly_sig[127] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11093 VGND _043_ a_13153_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11094 a_29541_12559# a_29375_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11096 tdc0.w_dly_sig_n[84] tdc0.w_dly_sig[83] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11097 a_3226_14191# a_2953_14197# a_3141_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11098 VGND clknet_4_8_0_clk a_16587_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11099 a_17329_7369# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X11100 tdc0.o_result[162] a_10627_3035# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11101 VGND tdc0.w_dly_sig_n[54] tdc0.w_dly_sig[55] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11103 a_24593_15599# _014_ a_24183_15511# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X11104 tdc0.w_dly_sig_n[106] tdc0.w_dly_sig[106] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11105 tdc0.w_dly_sig_n[79] tdc0.w_dly_sig[79] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11106 a_10309_10217# a_9319_9845# a_10183_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11107 tdc0.w_dly_sig[141] tdc0.w_dly_sig_n[139] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11108 tdc0.o_result[125] a_7867_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11109 tdc0.w_dly_sig[6] tdc0.w_dly_sig_n[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11110 VGND tdc0.w_dly_sig[155] tdc0.w_dly_sig_n[155] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11111 _069_ a_19931_4737# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X11112 VGND tdc0.w_dly_sig_n[52] tdc0.w_dly_sig[53] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11113 a_12851_11837# a_12153_11471# a_12594_11583# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11114 tdc0.w_dly_sig_n[131] tdc0.w_dly_sig[131] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11116 a_4797_6031# tdc0.w_dly_sig[147] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11117 tdc0.w_dly_sig[75] tdc0.w_dly_sig_n[73] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11118 VGND tdc0.w_dly_sig_n[129] tdc0.w_dly_sig[131] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11119 a_16833_10383# _034_ a_16761_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11120 a_2122_11837# a_1683_11471# a_2037_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11121 a_7883_10927# a_7019_10933# a_7626_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11122 tdc0.w_dly_sig_n[166] tdc0.w_dly_sig[166] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11124 VGND tdc0.w_dly_sig[142] tdc0.w_dly_sig_n[142] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11125 VGND a_17435_17429# a_17393_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11126 tdc0.w_dly_sig[90] tdc0.w_dly_sig_n[89] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11127 VPWR a_15170_2197# a_15097_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11128 VGND tdc0.w_dly_sig[140] tdc0.w_dly_sig_n[140] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11129 a_29090_13380# a_28890_13225# a_29239_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X11130 a_14865_3677# _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X11131 a_10777_8207# tdc0.w_dly_sig[78] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11132 a_13643_13647# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11133 tdc0.w_dly_sig_n[178] tdc0.w_dly_sig[178] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11134 a_22466_12533# a_22259_12533# a_22642_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X11135 VPWR a_14721_11445# _091_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X11136 a_12153_2223# a_11619_2229# a_12058_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11137 a_24490_18820# a_24283_18761# a_24666_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X11138 a_7553_10927# a_7019_10933# a_7458_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11139 VGND a_9431_9563# a_9389_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11140 a_17535_14191# a_16753_14197# a_17451_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11141 VPWR tdc0.w_dly_sig_n[143] tdc0.w_dly_sig[144] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11142 VGND tdc0.w_dly_sig[24] tdc0.w_dly_sig_n[24] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11143 clknet_4_14_0_clk a_26882_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11144 VGND _173_ a_15299_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11145 a_13633_11721# tdc0.o_result[74] a_13551_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11146 a_29703_11159# a_29987_11145# a_29922_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X11147 a_26663_4007# a_26759_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X11148 VPWR tdc0.w_dly_sig[188] a_28425_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X11149 a_21675_15101# a_20893_14735# a_21591_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11151 a_4195_5487# a_3413_5493# a_4111_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11152 a_2079_5487# a_1297_5493# a_1995_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11154 a_21707_17673# clknet_4_12_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11155 a_16555_15797# clknet_4_12_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11156 a_21561_3677# _060_ a_21489_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11157 a_24419_18921# a_24283_18761# a_23999_18775# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X11158 uo_out[4] a_19225_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11160 VGND tdc0.w_dly_sig_n[137] tdc0.w_dly_sig[139] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11161 VGND a_18659_7895# _096_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X11162 VGND _070_ a_20543_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11163 a_4697_16911# a_3707_16911# a_4571_17277# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11164 tdc0.w_dly_sig[33] tdc0.w_dly_sig_n[32] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11165 tdc0.w_dly_sig_n[126] tdc0.w_dly_sig[125] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11166 tdc0.w_dly_sig_n[128] tdc0.w_dly_sig[127] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11167 clknet_4_1_0_clk a_6476_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11168 a_20521_14569# a_19531_14197# a_20395_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11169 VPWR _034_ a_13643_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X11170 VPWR tdc0.w_dly_sig[109] tdc0.w_dly_sig_n[109] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11171 tdc0.w_dly_sig_n[27] tdc0.w_dly_sig[27] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11172 tdc0.w_dly_sig_n[33] tdc0.w_dly_sig[33] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11173 VGND tdc0.w_dly_sig[185] tdc0.w_dly_sig_n[186] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11174 tdc0.w_dly_sig[49] tdc0.w_dly_sig_n[47] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11175 tdc0.w_dly_sig[77] tdc0.w_dly_sig_n[75] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11176 a_25019_13621# clknet_4_15_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11177 a_27639_5865# a_27510_5609# a_27219_5719# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X11178 a_17023_5487# a_16495_5487# _011_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11180 VPWR tdc0.w_dly_sig_n[79] tdc0.w_dly_sig[80] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11181 a_6979_6005# a_7270_6305# a_7221_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X11182 tdc0.w_dly_sig_n[28] tdc0.w_dly_sig[27] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11183 VGND a_17619_14165# a_17577_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11184 tdc0.w_dly_sig_n[9] tdc0.w_dly_sig[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11186 a_22277_15279# tdc0.w_dly_sig[64] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11187 VGND clknet_4_0_0_clk a_3523_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11188 tdc0.w_dly_sig[23] tdc0.w_dly_sig_n[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11190 _043_ a_17231_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X11191 tdc0.w_dly_sig_n[61] tdc0.w_dly_sig[61] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11192 VGND _107_ a_23913_8353# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X11194 tdc0.w_dly_sig[97] tdc0.w_dly_sig_n[96] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11195 VGND tdc0.w_dly_sig[53] tdc0.w_dly_sig_n[53] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11196 a_12736_5865# a_12337_5493# a_12610_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11197 a_26541_11837# a_26203_11623# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X11198 a_8286_7663# a_8013_7669# a_8201_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11199 tdc0.w_dly_sig[190] tdc0.w_dly_sig_n[189] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11200 a_1669_10927# tdc0.w_dly_sig[111] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11201 VPWR tdc0.w_dly_sig[4] tdc0.w_dly_sig_n[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11202 a_15637_10383# _022_ a_15565_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11203 a_25494_11837# a_25247_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X11204 VGND a_4371_10901# a_4329_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11205 a_22374_2500# a_22174_2345# a_22523_2589# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X11206 VGND a_6246_3967# a_6204_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11207 VGND tdc0.w_dly_sig[29] tdc0.w_dly_sig_n[30] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11208 VGND tdc0.w_dly_sig_n[188] tdc0.w_dly_sig[190] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11209 VGND a_24283_2741# a_24290_3041# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11211 VGND tdc0.w_dly_sig[191] tdc0.w_dly_sig_n[191] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11212 tdc0.w_dly_sig_n[175] tdc0.w_dly_sig[175] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11213 tdc0.w_dly_sig[96] tdc0.w_dly_sig_n[94] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11214 tdc0.w_dly_sig[105] tdc0.w_dly_sig_n[103] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11215 VPWR a_8895_3311# a_9063_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11216 tdc0.w_dly_sig[95] tdc0.w_dly_sig_n[94] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11217 tdc0.o_result[158] a_7591_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11218 tdc0.w_dly_sig[120] tdc0.w_dly_sig_n[118] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11219 VPWR a_25410_13103# clknet_4_15_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11220 VGND a_7258_10495# a_7216_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11221 tdc0.w_dly_sig[148] tdc0.w_dly_sig_n[146] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11222 VPWR _072_ a_5989_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X11223 a_10018_2197# a_9850_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11224 VGND clknet_4_1_0_clk a_1131_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11226 VPWR tdc0.w_dly_sig[66] tdc0.w_dly_sig_n[67] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11227 VGND tdc0.w_dly_sig_n[81] tdc0.w_dly_sig[83] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11228 a_26203_11623# a_26299_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X11229 a_22799_17687# a_22895_17687# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11230 VPWR tdc0.o_result[26] a_24344_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X11231 a_27158_9028# a_26958_8873# a_27307_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X11232 a_15262_15935# a_15094_16189# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11233 clknet_4_4_0_clk a_6550_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11234 a_21886_5461# a_21718_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11235 a_9949_2767# tdc0.w_dly_sig[163] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11236 VPWR tdc0.w_dly_sig[86] tdc0.w_dly_sig_n[87] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11237 a_7699_15101# a_6835_14735# a_7442_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11238 tdc0.w_dly_sig_n[180] tdc0.w_dly_sig[179] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11239 tdc0.w_dly_sig[29] tdc0.w_dly_sig_n[27] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11240 VGND tdc0.w_dly_sig[5] tdc0.w_dly_sig_n[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11241 tdc0.w_dly_sig[26] tdc0.w_dly_sig_n[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11242 a_11582_14165# a_11414_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X11243 VGND tdc0.w_dly_sig_n[174] tdc0.w_dly_sig[175] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11244 tdc0.w_dly_sig_n[2] tdc0.w_dly_sig[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11245 a_23303_3424# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11246 a_9926_9813# a_9758_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11247 a_12552_14735# a_12153_14735# a_12426_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11249 VGND tdc0.w_dly_sig[151] tdc0.w_dly_sig_n[151] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11250 a_27137_7119# a_26590_7393# a_26790_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X11251 VPWR tdc0.w_dly_sig[64] tdc0.w_dly_sig_n[65] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11252 a_7369_15101# a_6835_14735# a_7274_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11253 a_14729_2229# a_14563_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11254 a_29895_4617# clknet_4_10_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11255 tdc0.o_result[146] a_5475_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11256 tdc0.w_dly_sig_n[60] tdc0.w_dly_sig[59] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11257 _132_ a_5823_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X11258 a_6633_15285# a_6467_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11259 VPWR a_19487_11159# tdc0.o_result[32] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11260 tdc0.o_result[16] a_30683_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11261 a_2582_6575# a_2143_6581# a_2497_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11262 tdc0.w_dly_sig_n[33] tdc0.w_dly_sig[32] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11263 VGND a_12391_15279# a_12559_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11265 VPWR a_7626_10901# a_7553_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11266 a_28595_7284# tdc0.w_dly_sig[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11267 VGND a_21051_8359# tdc0.o_result[29] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11268 a_17808_12335# _010_ a_17688_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X11270 clknet_4_2_0_clk a_11260_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11272 tdc0.w_dly_sig[99] tdc0.w_dly_sig_n[97] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11274 a_4613_8751# tdc0.w_dly_sig[115] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11275 tdc0.w_dly_sig[55] tdc0.w_dly_sig_n[53] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11276 tdc0.w_dly_sig[85] tdc0.w_dly_sig_n[83] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11277 a_29437_12393# a_28890_12137# a_29090_12292# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X11278 clknet_4_3_0_clk a_10506_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11279 a_18137_16367# tdc0.w_dly_sig[61] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11280 tdc0.w_dly_sig_n[35] tdc0.w_dly_sig[35] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11281 a_27158_9028# a_26951_8969# a_27334_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X11282 a_19141_2601# a_18151_2229# a_19015_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11283 VGND clknet_4_7_0_clk a_14563_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11284 tdc0.w_dly_sig_n[43] tdc0.w_dly_sig[43] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11285 tdc0.w_dly_sig_n[21] tdc0.w_dly_sig[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11287 VGND tdc0.w_dly_sig[110] tdc0.w_dly_sig_n[111] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11288 a_21603_4007# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X11289 VGND a_28503_13335# tdc0.o_result[42] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11290 tdc0.w_dly_sig[98] tdc0.w_dly_sig_n[96] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11291 a_13722_6031# _044_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X11292 VPWR tdc0.w_dly_sig[9] tdc0.w_dly_sig_n[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11293 tdc0.w_dly_sig[52] tdc0.w_dly_sig_n[51] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11294 VPWR _034_ a_14151_10535# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X11295 _203_ a_11527_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X11296 a_23315_17833# a_23186_17577# a_22895_17687# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X11297 a_12594_11583# a_12426_11837# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X11298 VGND tdc0.w_dly_sig_n[169] tdc0.w_dly_sig[171] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11300 VPWR a_29090_12292# a_29019_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X11301 VGND a_24013_11445# _015_ VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X11302 tdc0.w_dly_sig_n[144] tdc0.w_dly_sig[144] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11303 a_13725_13647# tdc0.o_result[71] a_13643_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11304 VPWR clknet_4_1_0_clk a_4167_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11305 a_24218_4943# a_23903_5095# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X11306 a_23562_17455# a_23315_17833# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X11307 a_10827_11837# a_9963_11471# a_10570_11583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11308 tdc0.w_dly_sig[188] tdc0.w_dly_sig_n[186] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11309 VGND _017_ a_18037_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X11310 VPWR a_10259_4373# a_10175_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11311 a_13809_18549# a_13643_18549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11312 VGND a_11582_14165# a_11540_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11313 tdc0.w_dly_sig_n[47] tdc0.w_dly_sig[46] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11314 tdc0.w_dly_sig_n[94] tdc0.w_dly_sig[94] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11315 a_7423_14191# a_6725_14197# a_7166_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11316 a_2547_14013# a_1849_13647# a_2290_13759# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11317 VPWR tdc0.w_dly_sig_n[86] tdc0.w_dly_sig[87] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11318 a_14082_17455# a_13643_17461# a_13997_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11319 tdc0.w_dly_sig_n[145] tdc0.w_dly_sig[145] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11320 a_30005_6031# net25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11321 a_15318_8457# _099_ a_15238_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X11322 tdc0.w_dly_sig[131] tdc0.w_dly_sig_n[129] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11323 VGND clknet_4_2_0_clk a_12171_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11324 a_5943_16189# a_5161_15823# a_5859_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11325 a_17109_15823# a_16562_16097# a_16762_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X11326 a_10497_11837# a_9963_11471# a_10402_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11327 VPWR a_14583_3035# a_14499_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11328 a_10034_4221# a_9761_3855# a_9949_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11329 VGND a_3267_7637# a_3225_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11330 a_10221_14735# a_10055_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11331 a_25318_11445# a_25111_11445# a_25494_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X11332 tdc0.w_dly_sig[159] tdc0.w_dly_sig_n[157] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11333 a_5617_14735# a_4627_14735# a_5491_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11334 tdc0.w_dly_sig_n[4] tdc0.w_dly_sig[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11335 _175_ a_18151_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X11336 a_13459_3424# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11337 VPWR a_16923_16885# a_16930_17185# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11338 tdc0.w_dly_sig[79] tdc0.w_dly_sig_n[78] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11339 VGND a_22374_2500# a_22303_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X11340 tdc0.w_dly_sig_n[26] tdc0.w_dly_sig[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11341 a_14839_13897# _020_ a_14922_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X11343 a_20009_9839# a_19671_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X11344 a_12341_15823# tdc0.w_dly_sig[88] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11345 VGND tdc0.w_dly_sig[190] tdc0.w_dly_sig_n[191] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11346 a_11865_13469# _034_ a_11793_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11347 a_16826_14847# a_16658_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X11348 VGND a_15170_2197# a_15128_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11349 a_6357_5487# a_5823_5493# a_6262_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11350 VPWR a_22603_17277# a_22771_17179# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11351 clknet_4_13_0_clk a_19890_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11352 _056_ a_16547_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11353 a_13722_12559# _199_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X11354 a_22721_2601# a_22167_2441# a_22374_2500# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X11355 tdc0.w_dly_sig_n[181] tdc0.w_dly_sig[180] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11356 a_12023_18543# a_11159_18549# a_11766_18517# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11357 a_12391_15279# a_11527_15285# a_12134_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11358 VGND clknet_4_2_0_clk a_13551_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11359 a_17187_13799# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X11360 a_25283_14887# a_25379_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11361 a_25247_11471# a_25111_11445# a_24827_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X11362 a_4387_4399# a_3523_4405# a_4130_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11363 tdc0.w_dly_sig_n[13] tdc0.w_dly_sig[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11364 VGND a_24283_18761# a_24290_18665# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11365 VGND a_5115_11159# _131_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X11366 a_13082_4399# tdc0.o_result[141] a_12999_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11367 tdc0.o_result[151] a_6855_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11368 a_13724_6895# tdc0.o_result[109] a_13149_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X11369 VPWR tdc0.w_dly_sig[56] tdc0.w_dly_sig_n[56] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11370 tdc0.w_dly_sig_n[37] tdc0.w_dly_sig[37] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11371 VPWR tdc0.w_dly_sig[34] tdc0.w_dly_sig_n[35] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11372 VPWR a_24283_2741# a_24290_3041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11373 VGND a_21207_3035# a_21165_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11374 VGND net3 a_16999_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X11375 VGND tdc0.w_dly_sig[12] tdc0.w_dly_sig_n[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11376 a_12061_15279# a_11527_15285# a_11966_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11377 a_11693_18543# a_11159_18549# a_11598_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11378 clknet_4_12_0_clk a_21380_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11379 VPWR a_30239_12925# a_30407_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11380 tdc0.w_dly_sig[19] tdc0.w_dly_sig_n[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11381 a_27505_9129# a_26951_8969# a_27158_9028# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X11382 tdc0.w_dly_sig_n[97] tdc0.w_dly_sig[97] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11383 a_14802_10901# a_14634_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11384 VGND tdc0.w_dly_sig_n[30] tdc0.w_dly_sig[31] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11385 a_19513_15285# a_19347_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11386 VPWR a_18151_1135# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X11387 a_27873_10217# a_27319_10057# a_27526_10116# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X11389 a_22809_13793# _146_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11390 a_15285_12559# tdc0.w_dly_sig[73] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11391 a_15115_9545# _129_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X11392 uo_out[1] a_24653_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11393 VGND tdc0.w_dly_sig_n[49] tdc0.w_dly_sig[51] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11394 VGND a_6982_16341# a_6940_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11395 VGND a_16916_4373# _050_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
R31 tt_um_hpretl_tt06_tdc_v1_20.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11396 VPWR a_16543_17063# tdc0.o_result[59] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11397 a_20175_12559# tdc0.o_result[7] a_20697_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X11398 tdc0.w_dly_sig[176] tdc0.w_dly_sig_n[175] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11399 a_27334_8751# a_27087_9129# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X11400 VGND clknet_4_0_0_clk a_6559_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11401 tdc0.w_dly_sig_n[64] tdc0.w_dly_sig[64] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11402 VPWR clknet_0_clk a_12254_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11403 tdc0.w_dly_sig_n[50] tdc0.w_dly_sig[50] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11404 a_18073_5847# net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.122 ps=1.08 w=0.42 l=0.15
X11405 tdc0.w_dly_sig_n[14] tdc0.w_dly_sig[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11406 VGND tdc0.w_dly_sig_n[56] tdc0.w_dly_sig[57] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11408 a_20900_4943# tdc0.o_result[191] a_20325_5089# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X11409 a_13398_6575# _164_ a_13149_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X11410 a_11329_14191# tdc0.w_dly_sig[85] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11412 VGND a_23903_5095# tdc0.o_result[23] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11413 VPWR tdc0.w_dly_sig[18] tdc0.w_dly_sig_n[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11414 a_16547_7093# _021_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X11415 VGND _114_ a_17967_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11416 tdc0.w_dly_sig_n[184] tdc0.w_dly_sig[184] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11417 a_2708_6953# a_2309_6581# a_2582_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11419 a_20881_11721# tdc0.o_result[0] a_21071_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X11420 VPWR tdc0.w_dly_sig_n[93] tdc0.w_dly_sig[95] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11421 a_26422_9269# a_26215_9269# a_26598_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X11422 a_4995_10633# _008_ a_5077_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11423 a_23075_4007# tdc0.o_result[184] a_23309_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11424 a_26882_12559# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11425 a_26387_17063# a_26483_16885# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11426 VGND a_19338_2741# a_19267_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X11427 a_8197_3317# a_8031_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11428 VPWR tdc0.w_dly_sig[176] tdc0.w_dly_sig_n[176] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11429 tdc0.w_dly_sig[151] tdc0.w_dly_sig_n[150] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11430 VPWR tdc0.w_dly_sig[84] tdc0.w_dly_sig_n[84] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11431 tdc0.w_dly_sig_n[8] tdc0.w_dly_sig[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11432 VGND _102_ a_17218_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X11433 a_2401_7669# a_2235_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11434 a_29998_8751# a_29559_8757# a_29913_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11435 VGND a_4038_11583# a_3996_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11436 tdc0.w_dly_sig_n[165] tdc0.w_dly_sig[164] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11437 a_23386_17732# a_23179_17673# a_23562_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X11438 VPWR a_17083_15101# a_17251_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11439 tdc0.w_dly_sig[43] tdc0.w_dly_sig_n[41] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11440 _055_ a_20945_13675# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X11441 VPWR _060_ a_18935_3543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X11442 VPWR tdc0.w_dly_sig_n[109] tdc0.w_dly_sig[110] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11443 a_3693_10927# tdc0.w_dly_sig[117] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11444 VPWR a_29803_5705# a_29810_5609# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11446 VGND tdc0.w_dly_sig[31] tdc0.w_dly_sig_n[32] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11447 a_20138_14165# a_19970_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11448 VPWR a_16127_4943# _060_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X11450 VGND a_2915_4399# a_3083_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11452 VGND tdc0.w_dly_sig[156] tdc0.w_dly_sig_n[157] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11453 a_19150_8207# tdc0.o_result[101] a_19069_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
C0 uio_in[7] VGND 0.182f
C1 uio_in[6] VGND 0.182f
C2 uio_in[5] VGND 0.182f
C3 uio_in[4] VGND 0.182f
C4 uio_in[3] VGND 0.182f
C5 uio_in[2] VGND 0.182f
C6 uio_in[1] VGND 0.182f
C7 uio_in[0] VGND 0.182f
C8 ui_in[2] VGND 0.182f
C9 ui_in[1] VGND 0.182f
C10 rst_n VGND 0.182f
C11 ena VGND 0.182f
C12 uio_oe[5] VGND 1.07f
C13 ui_in[5] VGND 1.18f
C14 ui_in[3] VGND 0.747f
C15 ui_in[7] VGND 1.01f
C16 ui_in[6] VGND 1.01f
C17 ui_in[4] VGND 1.2f
C18 uio_oe[4] VGND 1.24f
C19 uio_oe[0] VGND 1.13f
C20 uio_out[0] VGND 1.16f
C21 uo_out[1] VGND 3.48f
C22 uo_out[3] VGND 5.75f
C23 clk VGND 11.2f
C24 ui_in[0] VGND 1.25f
C25 uo_out[2] VGND 4.9f
C26 uo_out[0] VGND 4.85f
C27 uo_out[4] VGND 4.68f
C28 uo_out[5] VGND 3.62f
C29 uo_out[6] VGND 4.26f
C30 uo_out[7] VGND 3.87f
C31 uio_oe[1] VGND 1.04f
C32 uio_oe[2] VGND 1.21f
C33 uio_out[7] VGND 1.13f
C34 uio_oe[7] VGND 1.33f
C35 uio_out[3] VGND 1.09f
C36 uio_out[6] VGND 1.09f
C37 uio_oe[3] VGND 1.09f
C38 uio_out[2] VGND 1.09f
C39 uio_out[1] VGND 1.09f
C40 uio_out[4] VGND 1.39f
C41 uio_oe[6] VGND 1.56f
C42 uio_out[5] VGND 1.1f
C43 VPWR VGND 2.2p
C44 tt_um_hpretl_tt06_tdc_v1_12.HI VGND 0.415f $ **FLOATING
C45 a_22461_591# VGND 0.23f $ **FLOATING
C46 a_22971_957# VGND 0.609f $ **FLOATING
C47 a_23139_859# VGND 0.817f $ **FLOATING
C48 a_22546_957# VGND 0.626f $ **FLOATING
C49 a_22714_703# VGND 0.581f $ **FLOATING
C50 a_22273_591# VGND 1.43f $ **FLOATING
C51 a_22107_591# VGND 1.81f $ **FLOATING
C52 a_19057_591# VGND 0.23f $ **FLOATING
C53 a_19567_957# VGND 0.609f $ **FLOATING
C54 a_19735_859# VGND 0.817f $ **FLOATING
C55 a_19142_957# VGND 0.626f $ **FLOATING
C56 a_19310_703# VGND 0.581f $ **FLOATING
C57 a_18869_591# VGND 1.43f $ **FLOATING
C58 a_18703_591# VGND 1.81f $ **FLOATING
C59 a_18413_591# VGND 0.227f $ **FLOATING
C60 a_16481_591# VGND 0.23f $ **FLOATING
C61 a_18236_591# VGND 0.498f $ **FLOATING
C62 a_18130_591# VGND 0.578f $ **FLOATING
C63 a_17953_591# VGND 0.5f $ **FLOATING
C64 a_17634_591# VGND 0.535f $ **FLOATING
C65 a_16991_957# VGND 0.609f $ **FLOATING
C66 a_17159_859# VGND 0.817f $ **FLOATING
C67 a_16566_957# VGND 0.626f $ **FLOATING
C68 a_16734_703# VGND 0.581f $ **FLOATING
C69 a_16293_591# VGND 1.43f $ **FLOATING
C70 a_16127_591# VGND 1.81f $ **FLOATING
C71 a_15575_591# VGND 0.698f $ **FLOATING
C72 a_24745_1513# VGND 0.23f $ **FLOATING
C73 tdc0.w_dly_sig_n[178] VGND 1.99f $ **FLOATING
C74 a_11605_1135# VGND 0.23f $ **FLOATING
C75 a_24327_1513# VGND 0.581f $ **FLOATING
C76 a_24398_1412# VGND 0.626f $ **FLOATING
C77 a_24198_1257# VGND 1.43f $ **FLOATING
C78 a_24191_1353# VGND 1.81f $ **FLOATING
C79 a_23907_1367# VGND 0.609f $ **FLOATING
C80 a_23811_1367# VGND 0.817f $ **FLOATING
C81 tdc0.w_dly_sig_n[181] VGND 2.2f $ **FLOATING
C82 tdc0.w_dly_sig[180] VGND 2.84f $ **FLOATING
C83 tdc0.w_dly_sig_n[179] VGND 2.03f $ **FLOATING
C84 tdc0.w_dly_sig_n[176] VGND 1.92f $ **FLOATING
C85 a_18151_1135# VGND 1.2f $ **FLOATING
C86 a_17507_1143# VGND 0.648f $ **FLOATING
C87 a_16219_1143# VGND 0.648f $ **FLOATING
C88 tdc0.w_dly_sig[171] VGND 3.84f $ **FLOATING
C89 tdc0.w_dly_sig_n[169] VGND 2.31f $ **FLOATING
C90 a_12115_1135# VGND 0.609f $ **FLOATING
C91 a_12283_1109# VGND 0.817f $ **FLOATING
C92 a_11690_1135# VGND 0.626f $ **FLOATING
C93 a_11858_1109# VGND 0.581f $ **FLOATING
C94 a_11417_1141# VGND 1.43f $ **FLOATING
C95 a_11251_1141# VGND 1.81f $ **FLOATING
C96 tdc0.w_dly_sig_n[166] VGND 1.75f $ **FLOATING
C97 tdc0.w_dly_sig_n[163] VGND 2.04f $ **FLOATING
C98 tt_um_hpretl_tt06_tdc_v1_11.HI VGND 0.415f $ **FLOATING
C99 a_26125_1679# VGND 0.23f $ **FLOATING
C100 tdc0.w_dly_sig[181] VGND 4.06f $ **FLOATING
C101 a_20713_1679# VGND 0.23f $ **FLOATING
C102 a_25707_1679# VGND 0.581f $ **FLOATING
C103 a_25778_1653# VGND 0.626f $ **FLOATING
C104 a_25571_1653# VGND 1.81f $ **FLOATING
C105 a_25578_1953# VGND 1.43f $ **FLOATING
C106 a_25287_1653# VGND 0.609f $ **FLOATING
C107 a_25191_1831# VGND 0.817f $ **FLOATING
C108 tdc0.w_dly_sig_n[182] VGND 2.35f $ **FLOATING
C109 tdc0.w_dly_sig[183] VGND 3.72f $ **FLOATING
C110 tdc0.w_dly_sig_n[180] VGND 2.34f $ **FLOATING
C111 a_21223_2045# VGND 0.609f $ **FLOATING
C112 a_21391_1947# VGND 0.817f $ **FLOATING
C113 a_20798_2045# VGND 0.626f $ **FLOATING
C114 a_20966_1791# VGND 0.581f $ **FLOATING
C115 a_20525_1679# VGND 1.43f $ **FLOATING
C116 tdc0.w_dly_sig[179] VGND 3.32f $ **FLOATING
C117 a_20359_1679# VGND 1.81f $ **FLOATING
C118 tdc0.w_dly_sig_n[175] VGND 2.01f $ **FLOATING
C119 tdc0.w_dly_sig_n[170] VGND 1.93f $ **FLOATING
C120 tdc0.w_dly_sig_n[168] VGND 2.18f $ **FLOATING
C121 tdc0.w_dly_sig_n[167] VGND 2.12f $ **FLOATING
C122 a_11145_1679# VGND 0.23f $ **FLOATING
C123 tdc0.w_dly_sig[175] VGND 4.19f $ **FLOATING
C124 tdc0.w_dly_sig_n[174] VGND 2.31f $ **FLOATING
C125 tdc0.w_dly_sig_n[173] VGND 2.18f $ **FLOATING
C126 tdc0.w_dly_sig_n[172] VGND 1.89f $ **FLOATING
C127 tdc0.w_dly_sig_n[171] VGND 1.99f $ **FLOATING
C128 tdc0.w_dly_sig[167] VGND 3.29f $ **FLOATING
C129 a_11655_2045# VGND 0.609f $ **FLOATING
C130 a_11823_1947# VGND 0.817f $ **FLOATING
C131 a_11230_2045# VGND 0.626f $ **FLOATING
C132 a_11398_1791# VGND 0.581f $ **FLOATING
C133 a_10957_1679# VGND 1.43f $ **FLOATING
C134 tdc0.w_dly_sig[165] VGND 3.7f $ **FLOATING
C135 a_10791_1679# VGND 1.81f $ **FLOATING
C136 tdc0.w_dly_sig_n[165] VGND 1.94f $ **FLOATING
C137 tdc0.w_dly_sig_n[164] VGND 1.97f $ **FLOATING
C138 tdc0.w_dly_sig_n[162] VGND 2.42f $ **FLOATING
C139 tdc0.w_dly_sig_n[160] VGND 1.72f $ **FLOATING
C140 tdc0.w_dly_sig_n[159] VGND 1.72f $ **FLOATING
C141 tt_um_hpretl_tt06_tdc_v1_7.HI VGND 0.415f $ **FLOATING
C142 a_22721_2601# VGND 0.23f $ **FLOATING
C143 a_18505_2223# VGND 0.23f $ **FLOATING
C144 a_16941_2223# VGND 0.23f $ **FLOATING
C145 a_14917_2223# VGND 0.23f $ **FLOATING
C146 a_13445_2223# VGND 0.23f $ **FLOATING
C147 a_11973_2223# VGND 0.23f $ **FLOATING
C148 a_9765_2223# VGND 0.23f $ **FLOATING
C149 a_8293_2223# VGND 0.23f $ **FLOATING
C150 tdc0.w_dly_sig_n[161] VGND 2.24f $ **FLOATING
C151 tdc0.w_dly_sig_n[158] VGND 1.84f $ **FLOATING
C152 tdc0.w_dly_sig_n[184] VGND 2.23f $ **FLOATING
C153 tdc0.w_dly_sig_n[183] VGND 1.79f $ **FLOATING
C154 tdc0.w_dly_sig[182] VGND 3.08f $ **FLOATING
C155 a_22303_2601# VGND 0.581f $ **FLOATING
C156 a_22374_2500# VGND 0.626f $ **FLOATING
C157 a_22174_2345# VGND 1.43f $ **FLOATING
C158 a_22167_2441# VGND 1.81f $ **FLOATING
C159 a_21883_2455# VGND 0.609f $ **FLOATING
C160 a_21787_2455# VGND 0.817f $ **FLOATING
C161 tdc0.w_dly_sig_n[177] VGND 2.25f $ **FLOATING
C162 a_19015_2223# VGND 0.609f $ **FLOATING
C163 a_19183_2197# VGND 0.817f $ **FLOATING
C164 a_18590_2223# VGND 0.626f $ **FLOATING
C165 a_18758_2197# VGND 0.581f $ **FLOATING
C166 a_18317_2229# VGND 1.43f $ **FLOATING
C167 tdc0.w_dly_sig[176] VGND 3.54f $ **FLOATING
C168 a_18151_2229# VGND 1.81f $ **FLOATING
C169 a_17451_2223# VGND 0.609f $ **FLOATING
C170 a_17619_2197# VGND 0.817f $ **FLOATING
C171 a_17026_2223# VGND 0.626f $ **FLOATING
C172 a_17194_2197# VGND 0.581f $ **FLOATING
C173 a_16753_2229# VGND 1.43f $ **FLOATING
C174 tdc0.w_dly_sig[173] VGND 3.06f $ **FLOATING
C175 a_16587_2229# VGND 1.81f $ **FLOATING
C176 a_15427_2223# VGND 0.609f $ **FLOATING
C177 a_15595_2197# VGND 0.817f $ **FLOATING
C178 a_15002_2223# VGND 0.626f $ **FLOATING
C179 a_15170_2197# VGND 0.581f $ **FLOATING
C180 a_14729_2229# VGND 1.43f $ **FLOATING
C181 tdc0.w_dly_sig[169] VGND 4.39f $ **FLOATING
C182 a_14563_2229# VGND 1.81f $ **FLOATING
C183 a_13955_2223# VGND 0.609f $ **FLOATING
C184 a_14123_2197# VGND 0.817f $ **FLOATING
C185 a_13530_2223# VGND 0.626f $ **FLOATING
C186 a_13698_2197# VGND 0.581f $ **FLOATING
C187 a_13257_2229# VGND 1.43f $ **FLOATING
C188 tdc0.w_dly_sig[170] VGND 3.33f $ **FLOATING
C189 a_13091_2229# VGND 1.81f $ **FLOATING
C190 a_12483_2223# VGND 0.609f $ **FLOATING
C191 a_12651_2197# VGND 0.817f $ **FLOATING
C192 a_12058_2223# VGND 0.626f $ **FLOATING
C193 a_12226_2197# VGND 0.581f $ **FLOATING
C194 a_11785_2229# VGND 1.43f $ **FLOATING
C195 tdc0.w_dly_sig[166] VGND 3.96f $ **FLOATING
C196 a_11619_2229# VGND 1.81f $ **FLOATING
C197 a_10275_2223# VGND 0.609f $ **FLOATING
C198 a_10443_2197# VGND 0.817f $ **FLOATING
C199 a_9850_2223# VGND 0.626f $ **FLOATING
C200 a_10018_2197# VGND 0.581f $ **FLOATING
C201 a_9577_2229# VGND 1.43f $ **FLOATING
C202 tdc0.w_dly_sig[164] VGND 3.23f $ **FLOATING
C203 a_9411_2229# VGND 1.81f $ **FLOATING
C204 a_8803_2223# VGND 0.609f $ **FLOATING
C205 a_8971_2197# VGND 0.817f $ **FLOATING
C206 a_8378_2223# VGND 0.626f $ **FLOATING
C207 a_8546_2197# VGND 0.581f $ **FLOATING
C208 a_8105_2229# VGND 1.43f $ **FLOATING
C209 tdc0.w_dly_sig[162] VGND 3.2f $ **FLOATING
C210 a_7939_2229# VGND 1.81f $ **FLOATING
C211 tdc0.w_dly_sig_n[157] VGND 1.75f $ **FLOATING
C212 tdc0.w_dly_sig_n[156] VGND 1.75f $ **FLOATING
C213 tt_um_hpretl_tt06_tdc_v1_15.HI VGND 0.415f $ **FLOATING
C214 a_28425_2767# VGND 0.23f $ **FLOATING
C215 tdc0.w_dly_sig_n[186] VGND 1.97f $ **FLOATING
C216 tdc0.w_dly_sig[188] VGND 3.01f $ **FLOATING
C217 a_28007_2767# VGND 0.581f $ **FLOATING
C218 a_28078_2741# VGND 0.626f $ **FLOATING
C219 a_27871_2741# VGND 1.81f $ **FLOATING
C220 a_27878_3041# VGND 1.43f $ **FLOATING
C221 a_27587_2741# VGND 0.609f $ **FLOATING
C222 a_27491_2919# VGND 0.817f $ **FLOATING
C223 tdc0.w_dly_sig_n[185] VGND 2.04f $ **FLOATING
C224 a_24837_2767# VGND 0.23f $ **FLOATING
C225 a_22277_2767# VGND 0.23f $ **FLOATING
C226 tdc0.w_dly_sig[184] VGND 3.4f $ **FLOATING
C227 a_24419_2767# VGND 0.581f $ **FLOATING
C228 a_24490_2741# VGND 0.626f $ **FLOATING
C229 a_24283_2741# VGND 1.81f $ **FLOATING
C230 a_24290_3041# VGND 1.43f $ **FLOATING
C231 a_23999_2741# VGND 0.609f $ **FLOATING
C232 a_23903_2919# VGND 0.817f $ **FLOATING
C233 a_22787_3133# VGND 0.609f $ **FLOATING
C234 a_22955_3035# VGND 0.817f $ **FLOATING
C235 a_22362_3133# VGND 0.626f $ **FLOATING
C236 a_22530_2879# VGND 0.581f $ **FLOATING
C237 a_22089_2767# VGND 1.43f $ **FLOATING
C238 tdc0.w_dly_sig[185] VGND 4.04f $ **FLOATING
C239 a_21923_2767# VGND 1.81f $ **FLOATING
C240 a_20529_2767# VGND 0.23f $ **FLOATING
C241 a_21039_3133# VGND 0.609f $ **FLOATING
C242 a_21207_3035# VGND 0.817f $ **FLOATING
C243 a_20614_3133# VGND 0.626f $ **FLOATING
C244 a_20782_2879# VGND 0.581f $ **FLOATING
C245 a_20341_2767# VGND 1.43f $ **FLOATING
C246 tdc0.w_dly_sig[178] VGND 3.17f $ **FLOATING
C247 a_20175_2767# VGND 1.81f $ **FLOATING
C248 a_19685_2767# VGND 0.23f $ **FLOATING
C249 a_16113_2767# VGND 0.23f $ **FLOATING
C250 tdc0.w_dly_sig[177] VGND 3.91f $ **FLOATING
C251 a_19267_2767# VGND 0.581f $ **FLOATING
C252 a_19338_2741# VGND 0.626f $ **FLOATING
C253 a_19131_2741# VGND 1.81f $ **FLOATING
C254 a_19138_3041# VGND 1.43f $ **FLOATING
C255 a_18847_2741# VGND 0.609f $ **FLOATING
C256 a_18751_2919# VGND 0.817f $ **FLOATING
C257 a_16623_3133# VGND 0.609f $ **FLOATING
C258 a_16791_3035# VGND 0.817f $ **FLOATING
C259 a_16198_3133# VGND 0.626f $ **FLOATING
C260 a_16366_2879# VGND 0.581f $ **FLOATING
C261 a_15925_2767# VGND 1.43f $ **FLOATING
C262 tdc0.w_dly_sig[174] VGND 3.86f $ **FLOATING
C263 a_15759_2767# VGND 1.81f $ **FLOATING
C264 a_13905_2767# VGND 0.23f $ **FLOATING
C265 a_14415_3133# VGND 0.609f $ **FLOATING
C266 a_14583_3035# VGND 0.817f $ **FLOATING
C267 a_13990_3133# VGND 0.626f $ **FLOATING
C268 a_14158_2879# VGND 0.581f $ **FLOATING
C269 a_13717_2767# VGND 1.43f $ **FLOATING
C270 tdc0.w_dly_sig[172] VGND 4.9f $ **FLOATING
C271 a_13551_2767# VGND 1.81f $ **FLOATING
C272 tdc0.o_result[166] VGND 1.34f $ **FLOATING
C273 a_11605_2767# VGND 0.23f $ **FLOATING
C274 a_12815_2767# VGND 0.619f $ **FLOATING
C275 a_12115_3133# VGND 0.609f $ **FLOATING
C276 a_12283_3035# VGND 0.817f $ **FLOATING
C277 a_11690_3133# VGND 0.626f $ **FLOATING
C278 a_11858_2879# VGND 0.581f $ **FLOATING
C279 a_11417_2767# VGND 1.43f $ **FLOATING
C280 tdc0.w_dly_sig[168] VGND 4.26f $ **FLOATING
C281 a_11251_2767# VGND 1.81f $ **FLOATING
C282 a_9949_2767# VGND 0.23f $ **FLOATING
C283 a_10459_3133# VGND 0.609f $ **FLOATING
C284 a_10627_3035# VGND 0.817f $ **FLOATING
C285 a_10034_3133# VGND 0.626f $ **FLOATING
C286 a_10202_2879# VGND 0.581f $ **FLOATING
C287 a_9761_2767# VGND 1.43f $ **FLOATING
C288 tdc0.w_dly_sig[163] VGND 4.23f $ **FLOATING
C289 a_9595_2767# VGND 1.81f $ **FLOATING
C290 a_7189_2767# VGND 0.23f $ **FLOATING
C291 a_7699_3133# VGND 0.609f $ **FLOATING
C292 a_7867_3035# VGND 0.817f $ **FLOATING
C293 a_7274_3133# VGND 0.626f $ **FLOATING
C294 a_7442_2879# VGND 0.581f $ **FLOATING
C295 a_7001_2767# VGND 1.43f $ **FLOATING
C296 tdc0.w_dly_sig[160] VGND 3.53f $ **FLOATING
C297 a_6835_2767# VGND 1.81f $ **FLOATING
C298 a_5717_2767# VGND 0.23f $ **FLOATING
C299 a_6227_3133# VGND 0.609f $ **FLOATING
C300 a_6395_3035# VGND 0.817f $ **FLOATING
C301 a_5802_3133# VGND 0.626f $ **FLOATING
C302 a_5970_2879# VGND 0.581f $ **FLOATING
C303 a_5529_2767# VGND 1.43f $ **FLOATING
C304 tdc0.w_dly_sig[157] VGND 3.42f $ **FLOATING
C305 a_5363_2767# VGND 1.81f $ **FLOATING
C306 a_4245_2767# VGND 0.23f $ **FLOATING
C307 a_4755_3133# VGND 0.609f $ **FLOATING
C308 a_4923_3035# VGND 0.817f $ **FLOATING
C309 a_4330_3133# VGND 0.626f $ **FLOATING
C310 a_4498_2879# VGND 0.581f $ **FLOATING
C311 a_4057_2767# VGND 1.43f $ **FLOATING
C312 a_3891_2767# VGND 1.81f $ **FLOATING
C313 tdc0.w_dly_sig_n[155] VGND 2.26f $ **FLOATING
C314 tdc0.w_dly_sig[156] VGND 3.06f $ **FLOATING
C315 tdc0.w_dly_sig_n[154] VGND 1.91f $ **FLOATING
C316 a_29913_3311# VGND 0.23f $ **FLOATING
C317 a_25573_3689# VGND 0.23f $ **FLOATING
C318 a_8385_3311# VGND 0.23f $ **FLOATING
C319 a_6913_3311# VGND 0.23f $ **FLOATING
C320 a_3141_3311# VGND 0.23f $ **FLOATING
C321 a_30423_3311# VGND 0.609f $ **FLOATING
C322 a_30591_3285# VGND 0.817f $ **FLOATING
C323 a_29998_3311# VGND 0.626f $ **FLOATING
C324 a_30166_3285# VGND 0.581f $ **FLOATING
C325 a_29725_3317# VGND 1.43f $ **FLOATING
C326 a_29559_3317# VGND 1.81f $ **FLOATING
C327 tdc0.w_dly_sig_n[189] VGND 1.9f $ **FLOATING
C328 tdc0.w_dly_sig_n[187] VGND 2.46f $ **FLOATING
C329 tdc0.w_dly_sig_n[188] VGND 2.3f $ **FLOATING
C330 tdc0.w_dly_sig[187] VGND 3.86f $ **FLOATING
C331 a_25155_3689# VGND 0.581f $ **FLOATING
C332 a_25226_3588# VGND 0.626f $ **FLOATING
C333 a_25026_3433# VGND 1.43f $ **FLOATING
C334 a_25019_3529# VGND 1.81f $ **FLOATING
C335 a_24735_3543# VGND 0.609f $ **FLOATING
C336 a_24639_3543# VGND 0.817f $ **FLOATING
C337 a_23303_3424# VGND 0.619f $ **FLOATING
C338 tdc0.o_result[187] VGND 2.77f $ **FLOATING
C339 tdc0.o_result[178] VGND 1.5f $ **FLOATING
C340 a_21787_3543# VGND 0.619f $ **FLOATING
C341 tdc0.o_result[177] VGND 0.956f $ **FLOATING
C342 a_21327_3543# VGND 0.619f $ **FLOATING
C343 a_19899_3424# VGND 0.619f $ **FLOATING
C344 tdc0.o_result[174] VGND 1.85f $ **FLOATING
C345 tdc0.o_result[175] VGND 1.22f $ **FLOATING
C346 a_19395_3543# VGND 0.619f $ **FLOATING
C347 tdc0.o_result[176] VGND 1.16f $ **FLOATING
C348 a_18935_3543# VGND 0.619f $ **FLOATING
C349 a_17047_3424# VGND 0.619f $ **FLOATING
C350 tdc0.o_result[170] VGND 1.97f $ **FLOATING
C351 a_16311_3424# VGND 0.619f $ **FLOATING
C352 tdc0.o_result[168] VGND 1.28f $ **FLOATING
C353 tdc0.o_result[171] VGND 1.16f $ **FLOATING
C354 a_15163_3543# VGND 0.619f $ **FLOATING
C355 tdc0.o_result[169] VGND 1.37f $ **FLOATING
C356 a_14703_3543# VGND 0.619f $ **FLOATING
C357 a_14195_3424# VGND 0.619f $ **FLOATING
C358 tdc0.o_result[161] VGND 3.39f $ **FLOATING
C359 a_13459_3424# VGND 0.619f $ **FLOATING
C360 tdc0.o_result[160] VGND 2.53f $ **FLOATING
C361 a_12999_3424# VGND 0.619f $ **FLOATING
C362 tdc0.o_result[167] VGND 1.1f $ **FLOATING
C363 a_12539_3424# VGND 0.619f $ **FLOATING
C364 tdc0.o_result[163] VGND 1.88f $ **FLOATING
C365 a_8895_3311# VGND 0.609f $ **FLOATING
C366 a_9063_3285# VGND 0.817f $ **FLOATING
C367 a_8470_3311# VGND 0.626f $ **FLOATING
C368 a_8638_3285# VGND 0.581f $ **FLOATING
C369 a_8197_3317# VGND 1.43f $ **FLOATING
C370 tdc0.w_dly_sig[161] VGND 3.9f $ **FLOATING
C371 a_8031_3317# VGND 1.81f $ **FLOATING
C372 a_7423_3311# VGND 0.609f $ **FLOATING
C373 a_7591_3285# VGND 0.817f $ **FLOATING
C374 a_6998_3311# VGND 0.626f $ **FLOATING
C375 a_7166_3285# VGND 0.581f $ **FLOATING
C376 a_6725_3317# VGND 1.43f $ **FLOATING
C377 tdc0.w_dly_sig[159] VGND 3.8f $ **FLOATING
C378 a_6559_3317# VGND 1.81f $ **FLOATING
C379 a_3651_3311# VGND 0.609f $ **FLOATING
C380 a_3819_3285# VGND 0.817f $ **FLOATING
C381 a_3226_3311# VGND 0.626f $ **FLOATING
C382 a_3394_3285# VGND 0.581f $ **FLOATING
C383 a_2953_3317# VGND 1.43f $ **FLOATING
C384 tdc0.w_dly_sig[155] VGND 3.55f $ **FLOATING
C385 a_2787_3317# VGND 1.81f $ **FLOATING
C386 tdc0.w_dly_sig_n[153] VGND 1.86f $ **FLOATING
C387 tdc0.w_dly_sig[193] VGND 1.16f $ **FLOATING
C388 tdc0.w_dly_sig_n[191] VGND 2.16f $ **FLOATING
C389 tdc0.w_dly_sig_n[190] VGND 1.99f $ **FLOATING
C390 a_27597_3855# VGND 0.23f $ **FLOATING
C391 tdc0.w_dly_sig[190] VGND 3.53f $ **FLOATING
C392 a_27179_3855# VGND 0.581f $ **FLOATING
C393 a_27250_3829# VGND 0.626f $ **FLOATING
C394 a_27043_3829# VGND 1.81f $ **FLOATING
C395 a_27050_4129# VGND 1.43f $ **FLOATING
C396 a_26759_3829# VGND 0.609f $ **FLOATING
C397 a_26663_4007# VGND 0.817f $ **FLOATING
C398 a_25757_3855# VGND 0.23f $ **FLOATING
C399 tdc0.o_result[186] VGND 0.876f $ **FLOATING
C400 tdc0.o_result[179] VGND 2.3f $ **FLOATING
C401 tdc0.o_result[184] VGND 1.09f $ **FLOATING
C402 tdc0.o_result[189] VGND 2.47f $ **FLOATING
C403 tdc0.o_result[182] VGND 2.9f $ **FLOATING
C404 tdc0.o_result[190] VGND 5.94f $ **FLOATING
C405 tdc0.w_dly_sig[186] VGND 3.41f $ **FLOATING
C406 a_25339_3855# VGND 0.581f $ **FLOATING
C407 a_25410_3829# VGND 0.626f $ **FLOATING
C408 a_25203_3829# VGND 1.81f $ **FLOATING
C409 a_25210_4129# VGND 1.43f $ **FLOATING
C410 a_24919_3829# VGND 0.609f $ **FLOATING
C411 a_24823_4007# VGND 0.817f $ **FLOATING
C412 a_24363_4007# VGND 0.619f $ **FLOATING
C413 a_23903_4007# VGND 0.619f $ **FLOATING
C414 a_23075_4007# VGND 0.619f $ **FLOATING
C415 a_22615_4007# VGND 0.619f $ **FLOATING
C416 a_21603_4007# VGND 0.619f $ **FLOATING
C417 a_20359_3855# VGND 0.648f $ **FLOATING
C418 tdc0.o_result[172] VGND 1.3f $ **FLOATING
C419 tdc0.o_result[173] VGND 1.13f $ **FLOATING
C420 a_17048_4105# VGND 0.259f $ **FLOATING
C421 tdc0.o_result[154] VGND 5.77f $ **FLOATING
C422 tdc0.o_result[158] VGND 3.79f $ **FLOATING
C423 tdc0.o_result[159] VGND 2.45f $ **FLOATING
C424 a_9949_3855# VGND 0.23f $ **FLOATING
C425 a_19947_4007# VGND 0.619f $ **FLOATING
C426 a_17875_3855# VGND 0.619f $ **FLOATING
C427 a_17218_3855# VGND 0.672f $ **FLOATING
C428 _104_ VGND 0.91f $ **FLOATING
C429 _103_ VGND 2.78f $ **FLOATING
C430 _102_ VGND 1.29f $ **FLOATING
C431 tdc0.o_result[138] VGND 3.35f $ **FLOATING
C432 a_16635_4007# VGND 0.619f $ **FLOATING
C433 a_15391_3855# VGND 0.619f $ **FLOATING
C434 a_14931_3855# VGND 0.619f $ **FLOATING
C435 a_14287_3855# VGND 0.619f $ **FLOATING
C436 a_11527_3855# VGND 0.619f $ **FLOATING
C437 a_10459_4221# VGND 0.609f $ **FLOATING
C438 a_10627_4123# VGND 0.817f $ **FLOATING
C439 a_10034_4221# VGND 0.626f $ **FLOATING
C440 a_10202_3967# VGND 0.581f $ **FLOATING
C441 a_9761_3855# VGND 1.43f $ **FLOATING
C442 a_9595_3855# VGND 1.81f $ **FLOATING
C443 a_5993_3855# VGND 0.23f $ **FLOATING
C444 a_6503_4221# VGND 0.609f $ **FLOATING
C445 a_6671_4123# VGND 0.817f $ **FLOATING
C446 a_6078_4221# VGND 0.626f $ **FLOATING
C447 a_6246_3967# VGND 0.581f $ **FLOATING
C448 a_5805_3855# VGND 1.43f $ **FLOATING
C449 tdc0.w_dly_sig[158] VGND 4.13f $ **FLOATING
C450 a_5639_3855# VGND 1.81f $ **FLOATING
C451 a_3969_3855# VGND 0.23f $ **FLOATING
C452 a_4479_4221# VGND 0.609f $ **FLOATING
C453 a_4647_4123# VGND 0.817f $ **FLOATING
C454 a_4054_4221# VGND 0.626f $ **FLOATING
C455 a_4222_3967# VGND 0.581f $ **FLOATING
C456 a_3781_3855# VGND 1.43f $ **FLOATING
C457 tdc0.w_dly_sig[154] VGND 3.74f $ **FLOATING
C458 a_3615_3855# VGND 1.81f $ **FLOATING
C459 tdc0.w_dly_sig_n[152] VGND 2.1f $ **FLOATING
C460 a_30449_4777# VGND 0.23f $ **FLOATING
C461 tdc0.w_dly_sig_n[192] VGND 2.57f $ **FLOATING
C462 a_27597_4777# VGND 0.23f $ **FLOATING
C463 a_20848_4399# VGND 0.259f $ **FLOATING
C464 a_22001_4399# VGND 0.23f $ **FLOATING
C465 a_18888_4399# VGND 0.259f $ **FLOATING
C466 a_17876_4399# VGND 0.259f $ **FLOATING
C467 _056_ VGND 9.43f $ **FLOATING
C468 a_12999_4399# VGND 0.333f $ **FLOATING
C469 a_9581_4399# VGND 0.23f $ **FLOATING
C470 tdc0.o_result[143] VGND 3.71f $ **FLOATING
C471 a_7649_4399# VGND 0.23f $ **FLOATING
C472 a_6177_4399# VGND 0.23f $ **FLOATING
C473 a_3877_4399# VGND 0.23f $ **FLOATING
C474 a_2405_4399# VGND 0.23f $ **FLOATING
C475 tdc0.w_dly_sig[192] VGND 2.31f $ **FLOATING
C476 a_30031_4777# VGND 0.581f $ **FLOATING
C477 a_30102_4676# VGND 0.626f $ **FLOATING
C478 a_29902_4521# VGND 1.43f $ **FLOATING
C479 a_29895_4617# VGND 1.81f $ **FLOATING
C480 a_29611_4631# VGND 0.609f $ **FLOATING
C481 a_29515_4631# VGND 0.817f $ **FLOATING
C482 tdc0.w_dly_sig[191] VGND 2.99f $ **FLOATING
C483 tdc0.w_dly_sig[189] VGND 3.13f $ **FLOATING
C484 a_27179_4777# VGND 0.581f $ **FLOATING
C485 a_27250_4676# VGND 0.626f $ **FLOATING
C486 a_27050_4521# VGND 1.43f $ **FLOATING
C487 a_27043_4617# VGND 1.81f $ **FLOATING
C488 a_26759_4631# VGND 0.609f $ **FLOATING
C489 a_26663_4631# VGND 0.817f $ **FLOATING
C490 a_22511_4399# VGND 0.609f $ **FLOATING
C491 a_22679_4373# VGND 0.817f $ **FLOATING
C492 a_22086_4399# VGND 0.626f $ **FLOATING
C493 a_22254_4373# VGND 0.581f $ **FLOATING
C494 a_21813_4405# VGND 1.43f $ **FLOATING
C495 a_21647_4405# VGND 1.81f $ **FLOATING
C496 _182_ VGND 4.7f $ **FLOATING
C497 _183_ VGND 1.16f $ **FLOATING
C498 _184_ VGND 1.19f $ **FLOATING
C499 a_20417_4373# VGND 0.672f $ **FLOATING
C500 a_19931_4737# VGND 0.56f $ **FLOATING
C501 a_19058_4719# VGND 0.672f $ **FLOATING
C502 _204_ VGND 1.02f $ **FLOATING
C503 _203_ VGND 4.61f $ **FLOATING
C504 tdc0.o_result[151] VGND 5.98f $ **FLOATING
C505 a_18046_4719# VGND 0.672f $ **FLOATING
C506 _144_ VGND 0.857f $ **FLOATING
C507 _143_ VGND 3.07f $ **FLOATING
C508 tdc0.o_result[148] VGND 6.54f $ **FLOATING
C509 a_17231_4399# VGND 0.698f $ **FLOATING
C510 a_16916_4373# VGND 0.648f $ **FLOATING
C511 a_16547_4373# VGND 0.698f $ **FLOATING
C512 a_15333_4737# VGND 0.713f $ **FLOATING
C513 tdc0.o_result[181] VGND 4.45f $ **FLOATING
C514 a_14887_4631# VGND 0.619f $ **FLOATING
C515 a_13735_4512# VGND 0.619f $ **FLOATING
C516 tdc0.o_result[152] VGND 5.54f $ **FLOATING
C517 a_13082_4399# VGND 0.723f $ **FLOATING
C518 tdc0.o_result[165] VGND 1.59f $ **FLOATING
C519 tdc0.o_result[141] VGND 1.66f $ **FLOATING
C520 a_12171_4512# VGND 0.619f $ **FLOATING
C521 tdc0.o_result[156] VGND 4.16f $ **FLOATING
C522 a_11711_4512# VGND 0.619f $ **FLOATING
C523 tdc0.o_result[157] VGND 3.05f $ **FLOATING
C524 a_11251_4512# VGND 0.619f $ **FLOATING
C525 tdc0.o_result[153] VGND 3.72f $ **FLOATING
C526 a_10091_4399# VGND 0.609f $ **FLOATING
C527 a_10259_4373# VGND 0.817f $ **FLOATING
C528 a_9666_4399# VGND 0.626f $ **FLOATING
C529 a_9834_4373# VGND 0.581f $ **FLOATING
C530 a_9393_4405# VGND 1.43f $ **FLOATING
C531 a_9227_4405# VGND 1.81f $ **FLOATING
C532 a_8159_4399# VGND 0.609f $ **FLOATING
C533 a_8327_4373# VGND 0.817f $ **FLOATING
C534 a_7734_4399# VGND 0.626f $ **FLOATING
C535 a_7902_4373# VGND 0.581f $ **FLOATING
C536 a_7461_4405# VGND 1.43f $ **FLOATING
C537 a_7295_4405# VGND 1.81f $ **FLOATING
C538 a_6687_4399# VGND 0.609f $ **FLOATING
C539 a_6855_4373# VGND 0.817f $ **FLOATING
C540 a_6262_4399# VGND 0.626f $ **FLOATING
C541 a_6430_4373# VGND 0.581f $ **FLOATING
C542 a_5989_4405# VGND 1.43f $ **FLOATING
C543 tdc0.w_dly_sig[152] VGND 4.99f $ **FLOATING
C544 a_5823_4405# VGND 1.81f $ **FLOATING
C545 a_4387_4399# VGND 0.609f $ **FLOATING
C546 a_4555_4373# VGND 0.817f $ **FLOATING
C547 a_3962_4399# VGND 0.626f $ **FLOATING
C548 a_4130_4373# VGND 0.581f $ **FLOATING
C549 a_3689_4405# VGND 1.43f $ **FLOATING
C550 a_3523_4405# VGND 1.81f $ **FLOATING
C551 a_2915_4399# VGND 0.609f $ **FLOATING
C552 a_3083_4373# VGND 0.817f $ **FLOATING
C553 a_2490_4399# VGND 0.626f $ **FLOATING
C554 a_2658_4373# VGND 0.581f $ **FLOATING
C555 a_2217_4405# VGND 1.43f $ **FLOATING
C556 tdc0.w_dly_sig[153] VGND 4.07f $ **FLOATING
C557 a_2051_4405# VGND 1.81f $ **FLOATING
C558 tdc0.w_dly_sig_n[151] VGND 2.22f $ **FLOATING
C559 a_29361_4943# VGND 0.23f $ **FLOATING
C560 a_29871_5309# VGND 0.609f $ **FLOATING
C561 a_30039_5211# VGND 0.817f $ **FLOATING
C562 a_29446_5309# VGND 0.626f $ **FLOATING
C563 a_29614_5055# VGND 0.581f $ **FLOATING
C564 a_29173_4943# VGND 1.43f $ **FLOATING
C565 a_29007_4943# VGND 1.81f $ **FLOATING
C566 a_26309_4943# VGND 0.23f $ **FLOATING
C567 a_25891_4943# VGND 0.581f $ **FLOATING
C568 a_25962_4917# VGND 0.626f $ **FLOATING
C569 a_25755_4917# VGND 1.81f $ **FLOATING
C570 a_25762_5217# VGND 1.43f $ **FLOATING
C571 a_25471_4917# VGND 0.609f $ **FLOATING
C572 a_25375_5095# VGND 0.817f $ **FLOATING
C573 a_24837_4943# VGND 0.23f $ **FLOATING
C574 a_22790_5193# VGND 0.333f $ **FLOATING
C575 a_20756_5193# VGND 0.259f $ **FLOATING
C576 a_19928_5193# VGND 0.259f $ **FLOATING
C577 tdc0.o_result[12] VGND 6.07f $ **FLOATING
C578 _142_ VGND 1.1f $ **FLOATING
C579 _040_ VGND 6.68f $ **FLOATING
C580 _038_ VGND 8.54f $ **FLOATING
C581 a_24419_4943# VGND 0.581f $ **FLOATING
C582 a_24490_4917# VGND 0.626f $ **FLOATING
C583 a_24283_4917# VGND 1.81f $ **FLOATING
C584 a_24290_5217# VGND 1.43f $ **FLOATING
C585 a_23999_4917# VGND 0.609f $ **FLOATING
C586 a_23903_5095# VGND 0.817f $ **FLOATING
C587 tdc0.o_result[180] VGND 2.48f $ **FLOATING
C588 a_22633_4917# VGND 0.723f $ **FLOATING
C589 tdc0.o_result[191] VGND 4.52f $ **FLOATING
C590 _195_ VGND 3.59f $ **FLOATING
C591 a_20325_5089# VGND 0.672f $ **FLOATING
C592 tdc0.o_result[188] VGND 3.82f $ **FLOATING
C593 a_19497_5089# VGND 0.672f $ **FLOATING
C594 a_18751_5095# VGND 0.619f $ **FLOATING
C595 a_17383_5095# VGND 0.56f $ **FLOATING
C596 a_16999_4917# VGND 0.604f $ **FLOATING
C597 a_16733_4917# VGND 0.672f $ **FLOATING
C598 a_16127_4943# VGND 0.648f $ **FLOATING
C599 _005_ VGND 2.26f $ **FLOATING
C600 tdc0.o_result[162] VGND 2.83f $ **FLOATING
C601 _135_ VGND 3.54f $ **FLOATING
C602 _043_ VGND 9.27f $ **FLOATING
C603 tdc0.o_result[164] VGND 2.25f $ **FLOATING
C604 a_10961_4943# VGND 0.23f $ **FLOATING
C605 a_15609_4971# VGND 0.713f $ **FLOATING
C606 a_15203_5309# VGND 0.508f $ **FLOATING
C607 a_15023_5309# VGND 0.604f $ **FLOATING
C608 a_14103_4943# VGND 0.619f $ **FLOATING
C609 a_12999_4943# VGND 0.619f $ **FLOATING
C610 a_11471_5309# VGND 0.609f $ **FLOATING
C611 a_11639_5211# VGND 0.817f $ **FLOATING
C612 a_11046_5309# VGND 0.626f $ **FLOATING
C613 a_11214_5055# VGND 0.581f $ **FLOATING
C614 a_10773_4943# VGND 1.43f $ **FLOATING
C615 a_10607_4943# VGND 1.81f $ **FLOATING
C616 tdc0.w_dly_sig_n[141] VGND 1.99f $ **FLOATING
C617 tdc0.w_dly_sig_n[142] VGND 1.75f $ **FLOATING
C618 tdc0.w_dly_sig_n[144] VGND 1.72f $ **FLOATING
C619 tdc0.w_dly_sig[144] VGND 2.97f $ **FLOATING
C620 tdc0.w_dly_sig_n[150] VGND 1.9f $ **FLOATING
C621 a_30357_5865# VGND 0.23f $ **FLOATING
C622 a_28057_5865# VGND 0.23f $ **FLOATING
C623 a_23027_5487# VGND 0.333f $ **FLOATING
C624 tdc0.o_result[28] VGND 1.03f $ **FLOATING
C625 a_21633_5487# VGND 0.23f $ **FLOATING
C626 _196_ VGND 0.886f $ **FLOATING
C627 _136_ VGND 0.886f $ **FLOATING
C628 a_17023_5487# VGND 0.495f $ **FLOATING
C629 a_16665_5487# VGND 0.422f $ **FLOATING
C630 _202_ VGND 1.48f $ **FLOATING
C631 a_29939_5865# VGND 0.581f $ **FLOATING
C632 a_30010_5764# VGND 0.626f $ **FLOATING
C633 a_29810_5609# VGND 1.43f $ **FLOATING
C634 a_29803_5705# VGND 1.81f $ **FLOATING
C635 a_29519_5719# VGND 0.609f $ **FLOATING
C636 a_29423_5719# VGND 0.817f $ **FLOATING
C637 a_27639_5865# VGND 0.581f $ **FLOATING
C638 a_27710_5764# VGND 0.626f $ **FLOATING
C639 a_27510_5609# VGND 1.43f $ **FLOATING
C640 a_27503_5705# VGND 1.81f $ **FLOATING
C641 a_27219_5719# VGND 0.609f $ **FLOATING
C642 a_27123_5719# VGND 0.817f $ **FLOATING
C643 a_23110_5487# VGND 0.723f $ **FLOATING
C644 _050_ VGND 12.6f $ **FLOATING
C645 tdc0.o_result[183] VGND 1.9f $ **FLOATING
C646 tdc0.o_result[31] VGND 1f $ **FLOATING
C647 a_22143_5487# VGND 0.609f $ **FLOATING
C648 a_22311_5461# VGND 0.817f $ **FLOATING
C649 a_21718_5487# VGND 0.626f $ **FLOATING
C650 a_21886_5461# VGND 0.581f $ **FLOATING
C651 a_21445_5493# VGND 1.43f $ **FLOATING
C652 a_21279_5493# VGND 1.81f $ **FLOATING
C653 tdc0.o_result[23] VGND 2.27f $ **FLOATING
C654 a_20499_5719# VGND 0.619f $ **FLOATING
C655 tdc0.o_result[20] VGND 3.1f $ **FLOATING
C656 a_20039_5719# VGND 0.619f $ **FLOATING
C657 tdc0.o_result[15] VGND 4.97f $ **FLOATING
C658 a_19579_5719# VGND 0.619f $ **FLOATING
C659 tdc0.o_result[17] VGND 4.27f $ **FLOATING
C660 a_19119_5719# VGND 0.619f $ **FLOATING
C661 a_18196_5719# VGND 0.488f $ **FLOATING
C662 a_12525_5487# VGND 0.23f $ **FLOATING
C663 tdc0.w_dly_sig_n[143] VGND 2.04f $ **FLOATING
C664 a_6177_5487# VGND 0.23f $ **FLOATING
C665 a_3601_5487# VGND 0.23f $ **FLOATING
C666 a_1485_5487# VGND 0.23f $ **FLOATING
C667 a_17923_5719# VGND 0.601f $ **FLOATING
C668 a_16495_5487# VGND 1.45f $ **FLOATING
C669 a_14011_5487# VGND 0.698f $ **FLOATING
C670 a_13035_5487# VGND 0.609f $ **FLOATING
C671 a_13203_5461# VGND 0.817f $ **FLOATING
C672 a_12610_5487# VGND 0.626f $ **FLOATING
C673 a_12778_5461# VGND 0.581f $ **FLOATING
C674 a_12337_5493# VGND 1.43f $ **FLOATING
C675 a_12171_5493# VGND 1.81f $ **FLOATING
C676 clknet_4_2_0_clk VGND 14.3f $ **FLOATING
C677 a_11260_5461# VGND 1.98f $ **FLOATING
C678 tdc0.w_dly_sig_n[140] VGND 2.04f $ **FLOATING
C679 tdc0.w_dly_sig[142] VGND 3.78f $ **FLOATING
C680 tdc0.w_dly_sig[143] VGND 4.29f $ **FLOATING
C681 a_6687_5487# VGND 0.609f $ **FLOATING
C682 a_6855_5461# VGND 0.817f $ **FLOATING
C683 a_6262_5487# VGND 0.626f $ **FLOATING
C684 a_6430_5461# VGND 0.581f $ **FLOATING
C685 a_5989_5493# VGND 1.43f $ **FLOATING
C686 a_5823_5493# VGND 1.81f $ **FLOATING
C687 tdc0.w_dly_sig[145] VGND 6.08f $ **FLOATING
C688 tdc0.w_dly_sig_n[145] VGND 1.97f $ **FLOATING
C689 a_4111_5487# VGND 0.609f $ **FLOATING
C690 a_4279_5461# VGND 0.817f $ **FLOATING
C691 a_3686_5487# VGND 0.626f $ **FLOATING
C692 a_3854_5461# VGND 0.581f $ **FLOATING
C693 a_3413_5493# VGND 1.43f $ **FLOATING
C694 tdc0.w_dly_sig[148] VGND 2.92f $ **FLOATING
C695 a_3247_5493# VGND 1.81f $ **FLOATING
C696 a_1995_5487# VGND 0.609f $ **FLOATING
C697 a_2163_5461# VGND 0.817f $ **FLOATING
C698 a_1570_5487# VGND 0.626f $ **FLOATING
C699 a_1738_5461# VGND 0.581f $ **FLOATING
C700 a_1297_5493# VGND 1.43f $ **FLOATING
C701 tdc0.w_dly_sig[150] VGND 3.54f $ **FLOATING
C702 a_1131_5493# VGND 1.81f $ **FLOATING
C703 a_30005_6031# VGND 0.23f $ **FLOATING
C704 a_30515_6397# VGND 0.609f $ **FLOATING
C705 a_30683_6299# VGND 0.817f $ **FLOATING
C706 a_30090_6397# VGND 0.626f $ **FLOATING
C707 a_30258_6143# VGND 0.581f $ **FLOATING
C708 a_29817_6031# VGND 1.43f $ **FLOATING
C709 a_29651_6031# VGND 1.81f $ **FLOATING
C710 net28 VGND 1.5f $ **FLOATING
C711 clknet_4_8_0_clk VGND 13.2f $ **FLOATING
C712 a_29423_6196# VGND 0.524f $ **FLOATING
C713 tdc0.w_dly_sig_n[21] VGND 1.72f $ **FLOATING
C714 tdc0.w_dly_sig_n[22] VGND 2.46f $ **FLOATING
C715 tdc0.w_dly_sig_n[23] VGND 2.37f $ **FLOATING
C716 tdc0.w_dly_sig_n[24] VGND 2.43f $ **FLOATING
C717 tdc0.w_dly_sig_n[25] VGND 2.09f $ **FLOATING
C718 tdc0.w_dly_sig[24] VGND 3.07f $ **FLOATING
C719 a_21104_6005# VGND 1.98f $ **FLOATING
C720 a_20421_6031# VGND 0.23f $ **FLOATING
C721 a_17773_6281# VGND 0.214f $ **FLOATING
C722 tdc0.o_result[145] VGND 4.07f $ **FLOATING
C723 a_13552_6281# VGND 0.259f $ **FLOATING
C724 tdc0.o_result[149] VGND 5.34f $ **FLOATING
C725 a_11329_6031# VGND 0.23f $ **FLOATING
C726 tdc0.w_dly_sig[26] VGND 3.82f $ **FLOATING
C727 a_20003_6031# VGND 0.581f $ **FLOATING
C728 a_20074_6005# VGND 0.626f $ **FLOATING
C729 a_19867_6005# VGND 1.81f $ **FLOATING
C730 a_19874_6305# VGND 1.43f $ **FLOATING
C731 a_19583_6005# VGND 0.609f $ **FLOATING
C732 a_19487_6183# VGND 0.817f $ **FLOATING
C733 a_18737_6059# VGND 0.713f $ **FLOATING
C734 a_17691_6281# VGND 1.01f $ **FLOATING
C735 net3 VGND 8.2f $ **FLOATING
C736 a_15530_6077# VGND 0.611f $ **FLOATING
C737 net2 VGND 8.65f $ **FLOATING
C738 a_14379_6031# VGND 0.619f $ **FLOATING
C739 a_13722_6031# VGND 0.672f $ **FLOATING
C740 _044_ VGND 1.75f $ **FLOATING
C741 _041_ VGND 1.4f $ **FLOATING
C742 a_12723_6031# VGND 0.619f $ **FLOATING
C743 a_11839_6397# VGND 0.609f $ **FLOATING
C744 a_12007_6299# VGND 0.817f $ **FLOATING
C745 a_11414_6397# VGND 0.626f $ **FLOATING
C746 a_11582_6143# VGND 0.581f $ **FLOATING
C747 a_11141_6031# VGND 1.43f $ **FLOATING
C748 tdc0.w_dly_sig[141] VGND 3.74f $ **FLOATING
C749 a_10975_6031# VGND 1.81f $ **FLOATING
C750 tdc0.w_dly_sig[139] VGND 4.23f $ **FLOATING
C751 tdc0.w_dly_sig_n[139] VGND 1.97f $ **FLOATING
C752 tdc0.w_dly_sig_n[138] VGND 2.14f $ **FLOATING
C753 a_7817_6031# VGND 0.23f $ **FLOATING
C754 tdc0.o_result[136] VGND 3.74f $ **FLOATING
C755 a_4797_6031# VGND 0.23f $ **FLOATING
C756 a_7399_6031# VGND 0.581f $ **FLOATING
C757 a_7470_6005# VGND 0.626f $ **FLOATING
C758 a_7263_6005# VGND 1.81f $ **FLOATING
C759 a_7270_6305# VGND 1.43f $ **FLOATING
C760 a_6979_6005# VGND 0.609f $ **FLOATING
C761 a_6883_6183# VGND 0.817f $ **FLOATING
C762 a_5307_6397# VGND 0.609f $ **FLOATING
C763 a_5475_6299# VGND 0.817f $ **FLOATING
C764 a_4882_6397# VGND 0.626f $ **FLOATING
C765 a_5050_6143# VGND 0.581f $ **FLOATING
C766 a_4609_6031# VGND 1.43f $ **FLOATING
C767 a_4443_6031# VGND 1.81f $ **FLOATING
C768 tdc0.w_dly_sig_n[146] VGND 2.5f $ **FLOATING
C769 tdc0.w_dly_sig_n[147] VGND 2.53f $ **FLOATING
C770 tdc0.w_dly_sig_n[149] VGND 3.1f $ **FLOATING
C771 a_1301_6031# VGND 0.23f $ **FLOATING
C772 tdc0.w_dly_sig[146] VGND 3.82f $ **FLOATING
C773 tdc0.w_dly_sig[147] VGND 3.83f $ **FLOATING
C774 tdc0.w_dly_sig[149] VGND 3.93f $ **FLOATING
C775 tdc0.w_dly_sig_n[148] VGND 2.13f $ **FLOATING
C776 a_1811_6397# VGND 0.609f $ **FLOATING
C777 a_1979_6299# VGND 0.817f $ **FLOATING
C778 a_1386_6397# VGND 0.626f $ **FLOATING
C779 a_1554_6143# VGND 0.581f $ **FLOATING
C780 a_1113_6031# VGND 1.43f $ **FLOATING
C781 a_947_6031# VGND 1.81f $ **FLOATING
C782 net24 VGND 1.22f $ **FLOATING
C783 net25 VGND 1.24f $ **FLOATING
C784 tdc0.w_dly_sig[18] VGND 3.73f $ **FLOATING
C785 tdc0.w_dly_sig[21] VGND 4.81f $ **FLOATING
C786 a_23825_6953# VGND 0.23f $ **FLOATING
C787 a_17695_6575# VGND 1.29f $ **FLOATING
C788 _045_ VGND 3.21f $ **FLOATING
C789 a_18479_6895# VGND 0.473f $ **FLOATING
C790 a_15236_6575# VGND 0.259f $ **FLOATING
C791 a_17703_6895# VGND 0.473f $ **FLOATING
C792 _042_ VGND 2.38f $ **FLOATING
C793 a_13580_6575# VGND 0.259f $ **FLOATING
C794 a_30711_6794# VGND 0.524f $ **FLOATING
C795 a_29099_6575# VGND 0.524f $ **FLOATING
C796 tdc0.w_dly_sig_n[17] VGND 2.62f $ **FLOATING
C797 tdc0.w_dly_sig_n[18] VGND 3.15f $ **FLOATING
C798 tdc0.w_dly_sig_n[19] VGND 2.74f $ **FLOATING
C799 a_26514_6575# VGND 1.98f $ **FLOATING
C800 tdc0.w_dly_sig_n[20] VGND 2.9f $ **FLOATING
C801 tdc0.w_dly_sig[25] VGND 3.12f $ **FLOATING
C802 a_23407_6953# VGND 0.581f $ **FLOATING
C803 a_23478_6852# VGND 0.626f $ **FLOATING
C804 a_23278_6697# VGND 1.43f $ **FLOATING
C805 a_23271_6793# VGND 1.81f $ **FLOATING
C806 a_22987_6807# VGND 0.609f $ **FLOATING
C807 a_22891_6807# VGND 0.817f $ **FLOATING
C808 tdc0.w_dly_sig_n[26] VGND 2.12f $ **FLOATING
C809 tdc0.w_dly_sig_n[27] VGND 2.08f $ **FLOATING
C810 tdc0.o_result[16] VGND 5.87f $ **FLOATING
C811 a_19395_6807# VGND 0.619f $ **FLOATING
C812 a_17323_6575# VGND 0.698f $ **FLOATING
C813 a_16401_6691# VGND 0.601f $ **FLOATING
C814 a_16301_6575# VGND 0.488f $ **FLOATING
C815 a_11329_6575# VGND 0.23f $ **FLOATING
C816 tdc0.w_dly_sig_n[137] VGND 2.18f $ **FLOATING
C817 tdc0.w_dly_sig[137] VGND 3.18f $ **FLOATING
C818 clknet_4_0_0_clk VGND 19.2f $ **FLOATING
C819 a_2497_6575# VGND 0.23f $ **FLOATING
C820 tdc0.o_result[25] VGND 2.66f $ **FLOATING
C821 _078_ VGND 2.7f $ **FLOATING
C822 _079_ VGND 2.21f $ **FLOATING
C823 a_14805_6549# VGND 0.672f $ **FLOATING
C824 a_14255_6835# VGND 1.2f $ **FLOATING
C825 tdc0.o_result[109] VGND 5.97f $ **FLOATING
C826 _162_ VGND 2f $ **FLOATING
C827 _163_ VGND 7.27f $ **FLOATING
C828 _164_ VGND 0.935f $ **FLOATING
C829 a_13149_6549# VGND 0.672f $ **FLOATING
C830 a_12539_6688# VGND 0.619f $ **FLOATING
C831 _060_ VGND 12.8f $ **FLOATING
C832 tdc0.o_result[147] VGND 4.63f $ **FLOATING
C833 a_11839_6575# VGND 0.609f $ **FLOATING
C834 a_12007_6549# VGND 0.817f $ **FLOATING
C835 a_11414_6575# VGND 0.626f $ **FLOATING
C836 a_11582_6549# VGND 0.581f $ **FLOATING
C837 a_11141_6581# VGND 1.43f $ **FLOATING
C838 tdc0.w_dly_sig[140] VGND 3.48f $ **FLOATING
C839 a_10975_6581# VGND 1.81f $ **FLOATING
C840 tdc0.w_dly_sig_n[135] VGND 2.17f $ **FLOATING
C841 a_6476_6549# VGND 1.98f $ **FLOATING
C842 a_3007_6575# VGND 0.609f $ **FLOATING
C843 a_3175_6549# VGND 0.817f $ **FLOATING
C844 a_2582_6575# VGND 0.626f $ **FLOATING
C845 a_2750_6549# VGND 0.581f $ **FLOATING
C846 a_2309_6581# VGND 1.43f $ **FLOATING
C847 tdc0.w_dly_sig[151] VGND 3.77f $ **FLOATING
C848 a_2143_6581# VGND 1.81f $ **FLOATING
C849 net23 VGND 1.61f $ **FLOATING
C850 tdc0.w_dly_sig[16] VGND 5.08f $ **FLOATING
C851 a_30343_7284# VGND 0.524f $ **FLOATING
C852 a_29331_7284# VGND 0.524f $ **FLOATING
C853 tdc0.w_dly_sig_n[14] VGND 2.55f $ **FLOATING
C854 tdc0.w_dly_sig[19] VGND 3.74f $ **FLOATING
C855 a_28595_7284# VGND 0.524f $ **FLOATING
C856 a_27137_7119# VGND 0.23f $ **FLOATING
C857 tdc0.w_dly_sig[20] VGND 2.7f $ **FLOATING
C858 a_26719_7119# VGND 0.581f $ **FLOATING
C859 a_26790_7093# VGND 0.626f $ **FLOATING
C860 a_26583_7093# VGND 1.81f $ **FLOATING
C861 a_26590_7393# VGND 1.43f $ **FLOATING
C862 a_26299_7093# VGND 0.609f $ **FLOATING
C863 a_26203_7271# VGND 0.817f $ **FLOATING
C864 a_25665_7119# VGND 0.23f $ **FLOATING
C865 tdc0.w_dly_sig[22] VGND 3.66f $ **FLOATING
C866 a_25247_7119# VGND 0.581f $ **FLOATING
C867 a_25318_7093# VGND 0.626f $ **FLOATING
C868 a_25111_7093# VGND 1.81f $ **FLOATING
C869 a_25118_7393# VGND 1.43f $ **FLOATING
C870 a_24827_7093# VGND 0.609f $ **FLOATING
C871 a_24731_7271# VGND 0.817f $ **FLOATING
C872 a_22852_7093# VGND 1.98f $ **FLOATING
C873 tdc0.w_dly_sig[29] VGND 3.46f $ **FLOATING
C874 tdc0.w_dly_sig_n[28] VGND 1.93f $ **FLOATING
C875 a_20145_7119# VGND 0.23f $ **FLOATING
C876 net6 VGND 9.34f $ **FLOATING
C877 _077_ VGND 1.06f $ **FLOATING
C878 tdc0.w_dly_sig[28] VGND 3.61f $ **FLOATING
C879 a_19727_7119# VGND 0.581f $ **FLOATING
C880 a_19798_7093# VGND 0.626f $ **FLOATING
C881 a_19591_7093# VGND 1.81f $ **FLOATING
C882 a_19598_7393# VGND 1.43f $ **FLOATING
C883 a_19307_7093# VGND 0.609f $ **FLOATING
C884 a_19211_7271# VGND 0.817f $ **FLOATING
C885 a_17691_7119# VGND 1.2f $ **FLOATING
C886 _009_ VGND 1.45f $ **FLOATING
C887 a_16547_7093# VGND 0.698f $ **FLOATING
C888 a_15731_7271# VGND 0.611f $ **FLOATING
C889 a_15351_7093# VGND 0.698f $ **FLOATING
C890 _006_ VGND 1.27f $ **FLOATING
C891 a_14983_7093# VGND 0.698f $ **FLOATING
C892 a_14379_7119# VGND 0.619f $ **FLOATING
C893 tdc0.o_result[134] VGND 1.74f $ **FLOATING
C894 a_9305_7119# VGND 0.23f $ **FLOATING
C895 a_14064_7093# VGND 0.648f $ **FLOATING
C896 a_12907_7119# VGND 0.619f $ **FLOATING
C897 a_11435_7119# VGND 0.619f $ **FLOATING
C898 a_10506_7119# VGND 1.98f $ **FLOATING
C899 a_9815_7485# VGND 0.609f $ **FLOATING
C900 a_9983_7387# VGND 0.817f $ **FLOATING
C901 a_9390_7485# VGND 0.626f $ **FLOATING
C902 a_9558_7231# VGND 0.581f $ **FLOATING
C903 a_9117_7119# VGND 1.43f $ **FLOATING
C904 a_8951_7119# VGND 1.81f $ **FLOATING
C905 tdc0.w_dly_sig_n[136] VGND 1.98f $ **FLOATING
C906 a_7097_7119# VGND 0.23f $ **FLOATING
C907 a_7607_7485# VGND 0.609f $ **FLOATING
C908 a_7775_7387# VGND 0.817f $ **FLOATING
C909 a_7182_7485# VGND 0.626f $ **FLOATING
C910 a_7350_7231# VGND 0.581f $ **FLOATING
C911 a_6909_7119# VGND 1.43f $ **FLOATING
C912 a_6743_7119# VGND 1.81f $ **FLOATING
C913 tdc0.w_dly_sig[135] VGND 3.92f $ **FLOATING
C914 tdc0.w_dly_sig[136] VGND 3.43f $ **FLOATING
C915 a_4521_7119# VGND 0.23f $ **FLOATING
C916 tdc0.w_dly_sig_n[134] VGND 2.19f $ **FLOATING
C917 a_5031_7485# VGND 0.609f $ **FLOATING
C918 a_5199_7387# VGND 0.817f $ **FLOATING
C919 a_4606_7485# VGND 0.626f $ **FLOATING
C920 a_4774_7231# VGND 0.581f $ **FLOATING
C921 a_4333_7119# VGND 1.43f $ **FLOATING
C922 a_4167_7119# VGND 1.81f $ **FLOATING
C923 tdc0.o_result[113] VGND 5.77f $ **FLOATING
C924 a_1485_7119# VGND 0.23f $ **FLOATING
C925 a_1995_7485# VGND 0.609f $ **FLOATING
C926 a_2163_7387# VGND 0.817f $ **FLOATING
C927 a_1570_7485# VGND 0.626f $ **FLOATING
C928 a_1738_7231# VGND 0.581f $ **FLOATING
C929 a_1297_7119# VGND 1.43f $ **FLOATING
C930 a_1131_7119# VGND 1.81f $ **FLOATING
C931 a_29913_7663# VGND 0.23f $ **FLOATING
C932 tdc0.w_dly_sig[17] VGND 3.33f $ **FLOATING
C933 a_27689_8041# VGND 0.23f $ **FLOATING
C934 clknet_4_10_0_clk VGND 18.1f $ **FLOATING
C935 a_23381_7663# VGND 0.23f $ **FLOATING
C936 a_12448_7663# VGND 0.259f $ **FLOATING
C937 a_11329_7663# VGND 0.23f $ **FLOATING
C938 tdc0.o_result[131] VGND 1.86f $ **FLOATING
C939 a_8201_7663# VGND 0.23f $ **FLOATING
C940 tdc0.w_dly_sig[134] VGND 3.98f $ **FLOATING
C941 a_4061_7663# VGND 0.23f $ **FLOATING
C942 a_2589_7663# VGND 0.23f $ **FLOATING
C943 a_30423_7663# VGND 0.609f $ **FLOATING
C944 a_30591_7637# VGND 0.817f $ **FLOATING
C945 a_29998_7663# VGND 0.626f $ **FLOATING
C946 a_30166_7637# VGND 0.581f $ **FLOATING
C947 a_29725_7669# VGND 1.43f $ **FLOATING
C948 a_29559_7669# VGND 1.81f $ **FLOATING
C949 net27 VGND 1.28f $ **FLOATING
C950 a_27271_8041# VGND 0.581f $ **FLOATING
C951 a_27342_7940# VGND 0.626f $ **FLOATING
C952 a_27142_7785# VGND 1.43f $ **FLOATING
C953 a_27135_7881# VGND 1.81f $ **FLOATING
C954 a_26851_7895# VGND 0.609f $ **FLOATING
C955 a_26755_7895# VGND 0.817f $ **FLOATING
C956 a_25428_7637# VGND 1.98f $ **FLOATING
C957 a_23891_7663# VGND 0.609f $ **FLOATING
C958 a_24059_7637# VGND 0.817f $ **FLOATING
C959 a_23466_7663# VGND 0.626f $ **FLOATING
C960 a_23634_7637# VGND 0.581f $ **FLOATING
C961 a_23193_7669# VGND 1.43f $ **FLOATING
C962 tdc0.w_dly_sig[27] VGND 4.64f $ **FLOATING
C963 a_23027_7669# VGND 1.81f $ **FLOATING
C964 tdc0.w_dly_sig_n[29] VGND 1.87f $ **FLOATING
C965 tdc0.w_dly_sig_n[30] VGND 2.63f $ **FLOATING
C966 tdc0.o_result[21] VGND 2.67f $ **FLOATING
C967 a_20315_7895# VGND 0.619f $ **FLOATING
C968 tdc0.o_result[19] VGND 3.52f $ **FLOATING
C969 a_19855_7895# VGND 0.619f $ **FLOATING
C970 tdc0.o_result[13] VGND 5.7f $ **FLOATING
C971 a_19395_7895# VGND 0.619f $ **FLOATING
C972 tdc0.o_result[18] VGND 4.23f $ **FLOATING
C973 a_18659_7895# VGND 0.619f $ **FLOATING
C974 a_18059_7663# VGND 1.2f $ **FLOATING
C975 _000_ VGND 2.28f $ **FLOATING
C976 a_17503_7663# VGND 0.508f $ **FLOATING
C977 a_17323_7663# VGND 0.604f $ **FLOATING
C978 a_16739_7895# VGND 0.56f $ **FLOATING
C979 net5 VGND 8.37f $ **FLOATING
C980 a_16355_7969# VGND 0.604f $ **FLOATING
C981 net4 VGND 7.71f $ **FLOATING
C982 a_16179_7637# VGND 0.508f $ **FLOATING
C983 a_15101_7637# VGND 0.713f $ **FLOATING
C984 a_13997_7637# VGND 0.713f $ **FLOATING
C985 a_13275_7776# VGND 0.619f $ **FLOATING
C986 _024_ VGND 4.76f $ **FLOATING
C987 tdc0.o_result[133] VGND 4.7f $ **FLOATING
C988 a_12618_7983# VGND 0.672f $ **FLOATING
C989 _124_ VGND 1.29f $ **FLOATING
C990 _123_ VGND 3.47f $ **FLOATING
C991 _122_ VGND 1.3f $ **FLOATING
C992 tdc0.o_result[115] VGND 4.57f $ **FLOATING
C993 a_11839_7663# VGND 0.609f $ **FLOATING
C994 a_12007_7637# VGND 0.817f $ **FLOATING
C995 a_11414_7663# VGND 0.626f $ **FLOATING
C996 a_11582_7637# VGND 0.581f $ **FLOATING
C997 a_11141_7669# VGND 1.43f $ **FLOATING
C998 tdc0.w_dly_sig[138] VGND 4.01f $ **FLOATING
C999 a_10975_7669# VGND 1.81f $ **FLOATING
C1000 a_8711_7663# VGND 0.609f $ **FLOATING
C1001 a_8879_7637# VGND 0.817f $ **FLOATING
C1002 a_8286_7663# VGND 0.626f $ **FLOATING
C1003 a_8454_7637# VGND 0.581f $ **FLOATING
C1004 a_8013_7669# VGND 1.43f $ **FLOATING
C1005 a_7847_7669# VGND 1.81f $ **FLOATING
C1006 a_6476_7637# VGND 1.98f $ **FLOATING
C1007 tdc0.w_dly_sig_n[133] VGND 2.66f $ **FLOATING
C1008 a_4571_7663# VGND 0.609f $ **FLOATING
C1009 a_4739_7637# VGND 0.817f $ **FLOATING
C1010 a_4146_7663# VGND 0.626f $ **FLOATING
C1011 a_4314_7637# VGND 0.581f $ **FLOATING
C1012 a_3873_7669# VGND 1.43f $ **FLOATING
C1013 a_3707_7669# VGND 1.81f $ **FLOATING
C1014 a_3099_7663# VGND 0.609f $ **FLOATING
C1015 a_3267_7637# VGND 0.817f $ **FLOATING
C1016 a_2674_7663# VGND 0.626f $ **FLOATING
C1017 a_2842_7637# VGND 0.581f $ **FLOATING
C1018 a_2401_7669# VGND 1.43f $ **FLOATING
C1019 a_2235_7669# VGND 1.81f $ **FLOATING
C1020 tdc0.w_dly_sig_n[15] VGND 3.47f $ **FLOATING
C1021 tdc0.w_dly_sig_n[16] VGND 3.76f $ **FLOATING
C1022 tdc0.w_dly_sig_n[13] VGND 2.27f $ **FLOATING
C1023 tdc0.w_dly_sig[14] VGND 3.34f $ **FLOATING
C1024 tdc0.w_dly_sig[15] VGND 3.87f $ **FLOATING
C1025 tdc0.w_dly_sig[13] VGND 3.13f $ **FLOATING
C1026 a_27505_8207# VGND 0.23f $ **FLOATING
C1027 net26 VGND 2.36f $ **FLOATING
C1028 a_27087_8207# VGND 0.581f $ **FLOATING
C1029 a_27158_8181# VGND 0.626f $ **FLOATING
C1030 a_26951_8181# VGND 1.81f $ **FLOATING
C1031 a_26958_8481# VGND 1.43f $ **FLOATING
C1032 a_26667_8181# VGND 0.609f $ **FLOATING
C1033 a_26571_8359# VGND 0.817f $ **FLOATING
C1034 a_25849_8207# VGND 0.23f $ **FLOATING
C1035 a_24344_8457# VGND 0.259f $ **FLOATING
C1036 tdc0.o_result[22] VGND 1.32f $ **FLOATING
C1037 tdc0.w_dly_sig[23] VGND 3.28f $ **FLOATING
C1038 a_25431_8207# VGND 0.581f $ **FLOATING
C1039 a_25502_8181# VGND 0.626f $ **FLOATING
C1040 a_25295_8181# VGND 1.81f $ **FLOATING
C1041 a_25302_8481# VGND 1.43f $ **FLOATING
C1042 a_25011_8181# VGND 0.609f $ **FLOATING
C1043 a_24915_8359# VGND 0.817f $ **FLOATING
C1044 tdc0.o_result[26] VGND 0.863f $ **FLOATING
C1045 _108_ VGND 2.43f $ **FLOATING
C1046 a_23913_8353# VGND 0.672f $ **FLOATING
C1047 a_23303_8207# VGND 0.619f $ **FLOATING
C1048 a_21985_8207# VGND 0.23f $ **FLOATING
C1049 tdc0.o_result[29] VGND 1.01f $ **FLOATING
C1050 _030_ VGND 7.73f $ **FLOATING
C1051 a_18980_8457# VGND 0.259f $ **FLOATING
C1052 _105_ VGND 2.49f $ **FLOATING
C1053 _109_ VGND 3.48f $ **FLOATING
C1054 _021_ VGND 1.59f $ **FLOATING
C1055 _013_ VGND 4.16f $ **FLOATING
C1056 a_15420_8457# VGND 0.259f $ **FLOATING
C1057 _101_ VGND 1.76f $ **FLOATING
C1058 _007_ VGND 9.31f $ **FLOATING
C1059 a_13552_8457# VGND 0.259f $ **FLOATING
C1060 a_12264_8457# VGND 0.259f $ **FLOATING
C1061 a_10777_8207# VGND 0.23f $ **FLOATING
C1062 a_21567_8207# VGND 0.581f $ **FLOATING
C1063 a_21638_8181# VGND 0.626f $ **FLOATING
C1064 a_21431_8181# VGND 1.81f $ **FLOATING
C1065 a_21438_8481# VGND 1.43f $ **FLOATING
C1066 a_21147_8181# VGND 0.609f $ **FLOATING
C1067 a_21051_8359# VGND 0.817f $ **FLOATING
C1068 a_19855_8359# VGND 0.619f $ **FLOATING
C1069 a_19150_8207# VGND 0.672f $ **FLOATING
C1070 _160_ VGND 1.23f $ **FLOATING
C1071 _159_ VGND 0.815f $ **FLOATING
C1072 _158_ VGND 0.903f $ **FLOATING
C1073 a_17231_8457# VGND 0.702f $ **FLOATING
C1074 a_16713_8235# VGND 0.713f $ **FLOATING
C1075 a_15837_8181# VGND 0.713f $ **FLOATING
C1076 _098_ VGND 2.31f $ **FLOATING
C1077 _099_ VGND 0.854f $ **FLOATING
C1078 a_14989_8353# VGND 0.672f $ **FLOATING
C1079 a_14379_8207# VGND 0.619f $ **FLOATING
C1080 a_13722_8207# VGND 0.672f $ **FLOATING
C1081 _155_ VGND 0.942f $ **FLOATING
C1082 tdc0.o_result[117] VGND 4.74f $ **FLOATING
C1083 a_12434_8207# VGND 0.672f $ **FLOATING
C1084 _168_ VGND 4.31f $ **FLOATING
C1085 _167_ VGND 2.64f $ **FLOATING
C1086 tdc0.o_result[77] VGND 0.972f $ **FLOATING
C1087 a_11287_8573# VGND 0.609f $ **FLOATING
C1088 a_11455_8475# VGND 0.817f $ **FLOATING
C1089 a_10862_8573# VGND 0.626f $ **FLOATING
C1090 a_11030_8319# VGND 0.581f $ **FLOATING
C1091 a_10589_8207# VGND 1.43f $ **FLOATING
C1092 a_10423_8207# VGND 1.81f $ **FLOATING
C1093 tdc0.o_result[130] VGND 2.72f $ **FLOATING
C1094 a_8753_8207# VGND 0.23f $ **FLOATING
C1095 a_9263_8573# VGND 0.609f $ **FLOATING
C1096 a_9431_8475# VGND 0.817f $ **FLOATING
C1097 a_8838_8573# VGND 0.626f $ **FLOATING
C1098 a_9006_8319# VGND 0.581f $ **FLOATING
C1099 a_8565_8207# VGND 1.43f $ **FLOATING
C1100 a_8399_8207# VGND 1.81f $ **FLOATING
C1101 tdc0.w_dly_sig[132] VGND 2.96f $ **FLOATING
C1102 a_4797_8207# VGND 0.23f $ **FLOATING
C1103 tdc0.w_dly_sig_n[132] VGND 2.15f $ **FLOATING
C1104 a_5307_8573# VGND 0.609f $ **FLOATING
C1105 a_5475_8475# VGND 0.817f $ **FLOATING
C1106 a_4882_8573# VGND 0.626f $ **FLOATING
C1107 a_5050_8319# VGND 0.581f $ **FLOATING
C1108 a_4609_8207# VGND 1.43f $ **FLOATING
C1109 tdc0.w_dly_sig[133] VGND 3.51f $ **FLOATING
C1110 a_4443_8207# VGND 1.81f $ **FLOATING
C1111 a_29913_8751# VGND 0.23f $ **FLOATING
C1112 tdc0.w_dly_sig_n[12] VGND 2.54f $ **FLOATING
C1113 a_27505_9129# VGND 0.23f $ **FLOATING
C1114 a_24436_8751# VGND 0.259f $ **FLOATING
C1115 _106_ VGND 1.24f $ **FLOATING
C1116 a_19899_8751# VGND 0.333f $ **FLOATING
C1117 a_22829_8751# VGND 0.23f $ **FLOATING
C1118 a_17996_8751# VGND 0.259f $ **FLOATING
C1119 a_16350_8751# VGND 0.333f $ **FLOATING
C1120 a_14868_8751# VGND 0.259f $ **FLOATING
C1121 _097_ VGND 1.27f $ **FLOATING
C1122 a_30423_8751# VGND 0.609f $ **FLOATING
C1123 a_30591_8725# VGND 0.817f $ **FLOATING
C1124 a_29998_8751# VGND 0.626f $ **FLOATING
C1125 a_30166_8725# VGND 0.581f $ **FLOATING
C1126 a_29725_8757# VGND 1.43f $ **FLOATING
C1127 a_29559_8757# VGND 1.81f $ **FLOATING
C1128 tdc0.w_dly_sig_n[11] VGND 1.92f $ **FLOATING
C1129 a_27087_9129# VGND 0.581f $ **FLOATING
C1130 a_27158_9028# VGND 0.626f $ **FLOATING
C1131 a_26958_8873# VGND 1.43f $ **FLOATING
C1132 a_26951_8969# VGND 1.81f $ **FLOATING
C1133 a_26667_8983# VGND 0.609f $ **FLOATING
C1134 a_26571_8983# VGND 0.817f $ **FLOATING
C1135 tdc0.o_result[10] VGND 1.01f $ **FLOATING
C1136 a_25375_8983# VGND 0.619f $ **FLOATING
C1137 tdc0.o_result[14] VGND 1.47f $ **FLOATING
C1138 a_24915_8983# VGND 0.619f $ **FLOATING
C1139 tdc0.o_result[30] VGND 0.948f $ **FLOATING
C1140 _186_ VGND 0.818f $ **FLOATING
C1141 _188_ VGND 1.08f $ **FLOATING
C1142 a_24005_8725# VGND 0.672f $ **FLOATING
C1143 a_23339_8751# VGND 0.609f $ **FLOATING
C1144 a_23507_8725# VGND 0.817f $ **FLOATING
C1145 a_22914_8751# VGND 0.626f $ **FLOATING
C1146 a_23082_8725# VGND 0.581f $ **FLOATING
C1147 a_22641_8757# VGND 1.43f $ **FLOATING
C1148 a_22475_8757# VGND 1.81f $ **FLOATING
C1149 clknet_4_9_0_clk VGND 9.02f $ **FLOATING
C1150 tdc0.w_dly_sig[30] VGND 2.97f $ **FLOATING
C1151 a_19982_8751# VGND 0.723f $ **FLOATING
C1152 tdc0.o_result[9] VGND 5.42f $ **FLOATING
C1153 tdc0.o_result[137] VGND 4.43f $ **FLOATING
C1154 a_18383_8983# VGND 0.619f $ **FLOATING
C1155 _095_ VGND 0.779f $ **FLOATING
C1156 _096_ VGND 1.33f $ **FLOATING
C1157 a_17565_8725# VGND 0.672f $ **FLOATING
C1158 a_17139_8759# VGND 0.648f $ **FLOATING
C1159 tdc0.o_result[155] VGND 8.14f $ **FLOATING
C1160 _051_ VGND 14f $ **FLOATING
C1161 a_16193_8725# VGND 0.723f $ **FLOATING
C1162 _115_ VGND 3.28f $ **FLOATING
C1163 _116_ VGND 3.69f $ **FLOATING
C1164 a_14437_8725# VGND 0.672f $ **FLOATING
C1165 a_12999_8867# VGND 0.858f $ **FLOATING
C1166 _157_ VGND 1.24f $ **FLOATING
C1167 _161_ VGND 4.29f $ **FLOATING
C1168 _165_ VGND 1.63f $ **FLOATING
C1169 _169_ VGND 0.849f $ **FLOATING
C1170 a_9213_8751# VGND 0.23f $ **FLOATING
C1171 tdc0.w_dly_sig[131] VGND 3.16f $ **FLOATING
C1172 tdc0.w_dly_sig_n[131] VGND 2f $ **FLOATING
C1173 a_4613_8751# VGND 0.23f $ **FLOATING
C1174 a_11679_8983# VGND 0.56f $ **FLOATING
C1175 a_11159_8864# VGND 0.619f $ **FLOATING
C1176 _026_ VGND 10.1f $ **FLOATING
C1177 _025_ VGND 10.5f $ **FLOATING
C1178 tdc0.o_result[129] VGND 1.04f $ **FLOATING
C1179 a_9723_8751# VGND 0.609f $ **FLOATING
C1180 a_9891_8725# VGND 0.817f $ **FLOATING
C1181 a_9298_8751# VGND 0.626f $ **FLOATING
C1182 a_9466_8725# VGND 0.581f $ **FLOATING
C1183 a_9025_8757# VGND 1.43f $ **FLOATING
C1184 a_8859_8757# VGND 1.81f $ **FLOATING
C1185 a_5123_8751# VGND 0.609f $ **FLOATING
C1186 a_5291_8725# VGND 0.817f $ **FLOATING
C1187 a_4698_8751# VGND 0.626f $ **FLOATING
C1188 a_4866_8725# VGND 0.581f $ **FLOATING
C1189 a_4425_8757# VGND 1.43f $ **FLOATING
C1190 a_4259_8757# VGND 1.81f $ **FLOATING
C1191 tdc0.w_dly_sig_n[116] VGND 1.87f $ **FLOATING
C1192 tdc0.w_dly_sig[116] VGND 2.86f $ **FLOATING
C1193 tdc0.w_dly_sig_n[115] VGND 1.96f $ **FLOATING
C1194 tdc0.w_dly_sig[115] VGND 3.43f $ **FLOATING
C1195 tdc0.w_dly_sig_n[114] VGND 2.12f $ **FLOATING
C1196 tdc0.w_dly_sig[11] VGND 3.1f $ **FLOATING
C1197 a_24131_9295# VGND 0.594f $ **FLOATING
C1198 tdc0.w_dly_sig_n[10] VGND 2.08f $ **FLOATING
C1199 a_26769_9295# VGND 0.23f $ **FLOATING
C1200 a_24843_9545# VGND 0.399f $ **FLOATING
C1201 a_24381_9545# VGND 0.384f $ **FLOATING
C1202 a_24131_9545# VGND 0.388f $ **FLOATING
C1203 a_20709_9545# VGND 0.214f $ **FLOATING
C1204 a_20625_9545# VGND 0.167f $ **FLOATING
C1205 a_20204_9545# VGND 0.259f $ **FLOATING
C1206 _177_ VGND 0.666f $ **FLOATING
C1207 _185_ VGND 3.09f $ **FLOATING
C1208 _189_ VGND 3.03f $ **FLOATING
C1209 a_17168_9545# VGND 0.259f $ **FLOATING
C1210 a_16109_9545# VGND 0.214f $ **FLOATING
C1211 a_16025_9545# VGND 0.167f $ **FLOATING
C1212 _117_ VGND 1.25f $ **FLOATING
C1213 _125_ VGND 2.23f $ **FLOATING
C1214 _080_ VGND 1.93f $ **FLOATING
C1215 _181_ VGND 4.6f $ **FLOATING
C1216 a_13552_9545# VGND 0.259f $ **FLOATING
C1217 _089_ VGND 1.21f $ **FLOATING
C1218 a_12356_9545# VGND 0.259f $ **FLOATING
C1219 a_11237_9295# VGND 0.23f $ **FLOATING
C1220 a_26351_9295# VGND 0.581f $ **FLOATING
C1221 a_26422_9269# VGND 0.626f $ **FLOATING
C1222 a_26215_9269# VGND 1.81f $ **FLOATING
C1223 a_26222_9569# VGND 1.43f $ **FLOATING
C1224 a_25931_9269# VGND 0.609f $ **FLOATING
C1225 a_25835_9447# VGND 0.817f $ **FLOATING
C1226 a_24653_9545# VGND 1.44f $ **FLOATING
C1227 tdc0.o_result[1] VGND 1.02f $ **FLOATING
C1228 _090_ VGND 5.8f $ **FLOATING
C1229 _071_ VGND 2.06f $ **FLOATING
C1230 tdc0.w_dly_sig[31] VGND 3.05f $ **FLOATING
C1231 tdc0.w_dly_sig_n[31] VGND 1.92f $ **FLOATING
C1232 a_20543_9295# VGND 0.972f $ **FLOATING
C1233 _069_ VGND 3.83f $ **FLOATING
C1234 tdc0.o_result[185] VGND 4.84f $ **FLOATING
C1235 _070_ VGND 0.759f $ **FLOATING
C1236 _176_ VGND 2.93f $ **FLOATING
C1237 a_19773_9441# VGND 0.672f $ **FLOATING
C1238 a_19163_9545# VGND 0.702f $ **FLOATING
C1239 a_17567_9447# VGND 0.56f $ **FLOATING
C1240 tdc0.o_result[24] VGND 4.32f $ **FLOATING
C1241 a_16737_9441# VGND 0.672f $ **FLOATING
C1242 a_15943_9295# VGND 0.972f $ **FLOATING
C1243 _031_ VGND 10.8f $ **FLOATING
C1244 tdc0.o_result[27] VGND 2.74f $ **FLOATING
C1245 _113_ VGND 1.2f $ **FLOATING
C1246 a_15115_9545# VGND 0.702f $ **FLOATING
C1247 a_14563_9545# VGND 0.702f $ **FLOATING
C1248 a_13722_9295# VGND 0.672f $ **FLOATING
C1249 _179_ VGND 3.53f $ **FLOATING
C1250 _178_ VGND 1.9f $ **FLOATING
C1251 a_12526_9295# VGND 0.672f $ **FLOATING
C1252 _088_ VGND 3.24f $ **FLOATING
C1253 _087_ VGND 1.37f $ **FLOATING
C1254 tdc0.o_result[73] VGND 0.714f $ **FLOATING
C1255 a_11747_9661# VGND 0.609f $ **FLOATING
C1256 a_11915_9563# VGND 0.817f $ **FLOATING
C1257 a_11322_9661# VGND 0.626f $ **FLOATING
C1258 a_11490_9407# VGND 0.581f $ **FLOATING
C1259 a_11049_9295# VGND 1.43f $ **FLOATING
C1260 a_10883_9295# VGND 1.81f $ **FLOATING
C1261 clknet_4_3_0_clk VGND 8.41f $ **FLOATING
C1262 tdc0.o_result[126] VGND 2.45f $ **FLOATING
C1263 a_8753_9295# VGND 0.23f $ **FLOATING
C1264 a_9263_9661# VGND 0.609f $ **FLOATING
C1265 a_9431_9563# VGND 0.817f $ **FLOATING
C1266 a_8838_9661# VGND 0.626f $ **FLOATING
C1267 a_9006_9407# VGND 0.581f $ **FLOATING
C1268 a_8565_9295# VGND 1.43f $ **FLOATING
C1269 a_8399_9295# VGND 1.81f $ **FLOATING
C1270 tdc0.w_dly_sig[130] VGND 3f $ **FLOATING
C1271 tdc0.w_dly_sig_n[130] VGND 2.55f $ **FLOATING
C1272 a_5257_9295# VGND 0.23f $ **FLOATING
C1273 tdc0.w_dly_sig_n[129] VGND 2.14f $ **FLOATING
C1274 a_5767_9661# VGND 0.609f $ **FLOATING
C1275 a_5935_9563# VGND 0.817f $ **FLOATING
C1276 a_5342_9661# VGND 0.626f $ **FLOATING
C1277 a_5510_9407# VGND 0.581f $ **FLOATING
C1278 a_5069_9295# VGND 1.43f $ **FLOATING
C1279 a_4903_9295# VGND 1.81f $ **FLOATING
C1280 clknet_4_1_0_clk VGND 15.2f $ **FLOATING
C1281 tdc0.w_dly_sig_n[113] VGND 2.09f $ **FLOATING
C1282 tdc0.w_dly_sig[114] VGND 3.54f $ **FLOATING
C1283 tdc0.w_dly_sig_n[117] VGND 2.05f $ **FLOATING
C1284 a_29729_9839# VGND 0.23f $ **FLOATING
C1285 tdc0.w_dly_sig[10] VGND 3.47f $ **FLOATING
C1286 a_27873_10217# VGND 0.23f $ **FLOATING
C1287 a_23700_9839# VGND 0.259f $ **FLOATING
C1288 _129_ VGND 5.41f $ **FLOATING
C1289 a_20605_10217# VGND 0.23f $ **FLOATING
C1290 a_18679_9839# VGND 0.399f $ **FLOATING
C1291 a_18217_9839# VGND 0.384f $ **FLOATING
C1292 a_17967_9839# VGND 0.388f $ **FLOATING
C1293 a_15328_9839# VGND 0.259f $ **FLOATING
C1294 a_14012_9839# VGND 0.259f $ **FLOATING
C1295 a_17967_10159# VGND 0.594f $ **FLOATING
C1296 _084_ VGND 0.889f $ **FLOATING
C1297 _075_ VGND 0.848f $ **FLOATING
C1298 _180_ VGND 0.966f $ **FLOATING
C1299 tdc0.o_result[75] VGND 2.27f $ **FLOATING
C1300 a_12249_9839# VGND 0.23f $ **FLOATING
C1301 a_9673_9839# VGND 0.23f $ **FLOATING
C1302 tdc0.w_dly_sig_n[128] VGND 1.83f $ **FLOATING
C1303 a_2221_9839# VGND 0.23f $ **FLOATING
C1304 tdc0.w_dly_sig_n[112] VGND 1.99f $ **FLOATING
C1305 a_30239_9839# VGND 0.609f $ **FLOATING
C1306 a_30407_9813# VGND 0.817f $ **FLOATING
C1307 a_29814_9839# VGND 0.626f $ **FLOATING
C1308 a_29982_9813# VGND 0.581f $ **FLOATING
C1309 a_29541_9845# VGND 1.43f $ **FLOATING
C1310 tdc0.w_dly_sig[12] VGND 3.9f $ **FLOATING
C1311 a_29375_9845# VGND 1.81f $ **FLOATING
C1312 tdc0.w_dly_sig_n[9] VGND 2.41f $ **FLOATING
C1313 clknet_4_11_0_clk VGND 11.3f $ **FLOATING
C1314 a_27455_10217# VGND 0.581f $ **FLOATING
C1315 a_27526_10116# VGND 0.626f $ **FLOATING
C1316 a_27326_9961# VGND 1.43f $ **FLOATING
C1317 a_27319_10057# VGND 1.81f $ **FLOATING
C1318 a_27035_10071# VGND 0.609f $ **FLOATING
C1319 a_26939_10071# VGND 0.817f $ **FLOATING
C1320 _126_ VGND 3.89f $ **FLOATING
C1321 _128_ VGND 3.37f $ **FLOATING
C1322 a_23269_9813# VGND 0.672f $ **FLOATING
C1323 tdc0.w_dly_sig[32] VGND 4.85f $ **FLOATING
C1324 tdc0.w_dly_sig_n[32] VGND 2.33f $ **FLOATING
C1325 a_20187_10217# VGND 0.581f $ **FLOATING
C1326 a_20258_10116# VGND 0.626f $ **FLOATING
C1327 a_20058_9961# VGND 1.43f $ **FLOATING
C1328 a_20051_10057# VGND 1.81f $ **FLOATING
C1329 a_19767_10071# VGND 0.609f $ **FLOATING
C1330 a_19671_10071# VGND 0.817f $ **FLOATING
C1331 a_18489_9839# VGND 1.44f $ **FLOATING
C1332 tdc0.o_result[3] VGND 4.52f $ **FLOATING
C1333 _130_ VGND 2.42f $ **FLOATING
C1334 _114_ VGND 1.61f $ **FLOATING
C1335 a_16210_9839# VGND 4.03f $ **FLOATING
C1336 tdc0.o_result[33] VGND 2.55f $ **FLOATING
C1337 _082_ VGND 6.11f $ **FLOATING
C1338 _083_ VGND 2.56f $ **FLOATING
C1339 a_14897_9813# VGND 0.672f $ **FLOATING
C1340 a_14182_10159# VGND 0.672f $ **FLOATING
C1341 _033_ VGND 10.9f $ **FLOATING
C1342 _073_ VGND 3.98f $ **FLOATING
C1343 a_13367_9952# VGND 0.619f $ **FLOATING
C1344 tdc0.o_result[78] VGND 1.84f $ **FLOATING
C1345 a_12759_9839# VGND 0.609f $ **FLOATING
C1346 a_12927_9813# VGND 0.817f $ **FLOATING
C1347 a_12334_9839# VGND 0.626f $ **FLOATING
C1348 a_12502_9813# VGND 0.581f $ **FLOATING
C1349 a_12061_9845# VGND 1.43f $ **FLOATING
C1350 a_11895_9845# VGND 1.81f $ **FLOATING
C1351 a_10183_9839# VGND 0.609f $ **FLOATING
C1352 a_10351_9813# VGND 0.817f $ **FLOATING
C1353 a_9758_9839# VGND 0.626f $ **FLOATING
C1354 a_9926_9813# VGND 0.581f $ **FLOATING
C1355 a_9485_9845# VGND 1.43f $ **FLOATING
C1356 a_9319_9845# VGND 1.81f $ **FLOATING
C1357 tdc0.w_dly_sig[118] VGND 3.48f $ **FLOATING
C1358 tdc0.w_dly_sig_n[118] VGND 1.83f $ **FLOATING
C1359 a_2731_9839# VGND 0.609f $ **FLOATING
C1360 a_2899_9813# VGND 0.817f $ **FLOATING
C1361 a_2306_9839# VGND 0.626f $ **FLOATING
C1362 a_2474_9813# VGND 0.581f $ **FLOATING
C1363 a_2033_9845# VGND 1.43f $ **FLOATING
C1364 tdc0.w_dly_sig[113] VGND 3.05f $ **FLOATING
C1365 a_1867_9845# VGND 1.81f $ **FLOATING
C1366 a_30347_10357# VGND 1.33f $ **FLOATING
C1367 tdc0.w_dly_sig_n[8] VGND 1.92f $ **FLOATING
C1368 tdc0.w_dly_sig_n[2] VGND 1.83f $ **FLOATING
C1369 _638_.X VGND 0.226f $ **FLOATING
C1370 tdc0.w_dly_sig_n[1] VGND 2.45f $ **FLOATING
C1371 tdc0.o_result[35] VGND 0.902f $ **FLOATING
C1372 a_22645_10383# VGND 0.23f $ **FLOATING
C1373 a_25288_10357# VGND 0.648f $ **FLOATING
C1374 net1 VGND 4.98f $ **FLOATING
C1375 a_23155_10749# VGND 0.609f $ **FLOATING
C1376 a_23323_10651# VGND 0.817f $ **FLOATING
C1377 a_22730_10749# VGND 0.626f $ **FLOATING
C1378 a_22898_10495# VGND 0.581f $ **FLOATING
C1379 a_22457_10383# VGND 1.43f $ **FLOATING
C1380 a_22291_10383# VGND 1.81f $ **FLOATING
C1381 a_19881_10633# VGND 0.214f $ **FLOATING
C1382 a_19797_10633# VGND 0.167f $ **FLOATING
C1383 tdc0.w_dly_sig_n[33] VGND 2.04f $ **FLOATING
C1384 a_19715_10383# VGND 0.972f $ **FLOATING
C1385 tdc0.o_result[144] VGND 5.45f $ **FLOATING
C1386 a_18703_10383# VGND 0.648f $ **FLOATING
C1387 _175_ VGND 1.78f $ **FLOATING
C1388 _036_ VGND 1.07f $ **FLOATING
C1389 a_16109_10633# VGND 0.214f $ **FLOATING
C1390 a_16025_10633# VGND 0.167f $ **FLOATING
C1391 _032_ VGND 1.67f $ **FLOATING
C1392 _019_ VGND 7.93f $ **FLOATING
C1393 tdc0.o_result[120] VGND 5.63f $ **FLOATING
C1394 _081_ VGND 0.982f $ **FLOATING
C1395 _100_ VGND 1.57f $ **FLOATING
C1396 _074_ VGND 1.06f $ **FLOATING
C1397 _166_ VGND 1.6f $ **FLOATING
C1398 a_8481_10633# VGND 0.206f $ **FLOATING
C1399 a_7005_10383# VGND 0.23f $ **FLOATING
C1400 a_18151_10383# VGND 0.619f $ **FLOATING
C1401 _018_ VGND 3.95f $ **FLOATING
C1402 a_17467_10357# VGND 0.698f $ **FLOATING
C1403 a_16679_10383# VGND 0.619f $ **FLOATING
C1404 a_15943_10383# VGND 0.972f $ **FLOATING
C1405 _133_ VGND 5.75f $ **FLOATING
C1406 a_15483_10383# VGND 0.619f $ **FLOATING
C1407 a_15023_10383# VGND 0.619f $ **FLOATING
C1408 a_14563_10383# VGND 0.619f $ **FLOATING
C1409 a_14151_10535# VGND 0.619f $ **FLOATING
C1410 a_12539_10383# VGND 0.619f $ **FLOATING
C1411 a_8399_10633# VGND 0.804f $ **FLOATING
C1412 tdc0.o_result[112] VGND 3.22f $ **FLOATING
C1413 tdc0.o_result[128] VGND 0.747f $ **FLOATING
C1414 a_7515_10749# VGND 0.609f $ **FLOATING
C1415 a_7683_10651# VGND 0.817f $ **FLOATING
C1416 a_7090_10749# VGND 0.626f $ **FLOATING
C1417 a_7258_10495# VGND 0.581f $ **FLOATING
C1418 a_6817_10383# VGND 1.43f $ **FLOATING
C1419 a_6651_10383# VGND 1.81f $ **FLOATING
C1420 a_5077_10633# VGND 0.206f $ **FLOATING
C1421 a_4995_10633# VGND 0.804f $ **FLOATING
C1422 tdc0.o_result[150] VGND 2.81f $ **FLOATING
C1423 tdc0.w_dly_sig_n[119] VGND 1.94f $ **FLOATING
C1424 tdc0.w_dly_sig_n[111] VGND 1.98f $ **FLOATING
C1425 a_30541_11305# VGND 0.23f $ **FLOATING
C1426 tdc0.w_dly_sig[2] VGND 3.8f $ **FLOATING
C1427 a_24009_11305# VGND 0.23f $ **FLOATING
C1428 a_22261_11305# VGND 0.23f $ **FLOATING
C1429 a_20421_11305# VGND 0.23f $ **FLOATING
C1430 a_18127_10927# VGND 0.399f $ **FLOATING
C1431 a_17665_10927# VGND 0.384f $ **FLOATING
C1432 a_17415_10927# VGND 0.388f $ **FLOATING
C1433 a_16845_10927# VGND 0.214f $ **FLOATING
C1434 a_16761_10927# VGND 0.167f $ **FLOATING
C1435 tdc0.o_result[32] VGND 1.1f $ **FLOATING
C1436 a_17415_11247# VGND 0.594f $ **FLOATING
C1437 tdc0.o_result[76] VGND 1.23f $ **FLOATING
C1438 a_8573_10927# VGND 0.206f $ **FLOATING
C1439 a_14549_10927# VGND 0.23f $ **FLOATING
C1440 tdc0.w_dly_sig_n[77] VGND 2.04f $ **FLOATING
C1441 a_5989_10927# VGND 0.214f $ **FLOATING
C1442 a_5905_10927# VGND 0.167f $ **FLOATING
C1443 a_5261_10927# VGND 0.206f $ **FLOATING
C1444 a_7373_10927# VGND 0.23f $ **FLOATING
C1445 a_3693_10927# VGND 0.23f $ **FLOATING
C1446 tdc0.o_result[110] VGND 1.99f $ **FLOATING
C1447 a_1669_10927# VGND 0.23f $ **FLOATING
C1448 tdc0.w_dly_sig[9] VGND 3.86f $ **FLOATING
C1449 a_30123_11305# VGND 0.581f $ **FLOATING
C1450 a_30194_11204# VGND 0.626f $ **FLOATING
C1451 a_29994_11049# VGND 1.43f $ **FLOATING
C1452 a_29987_11145# VGND 1.81f $ **FLOATING
C1453 a_29703_11159# VGND 0.609f $ **FLOATING
C1454 a_29607_11159# VGND 0.817f $ **FLOATING
C1455 tdc0.w_dly_sig_n[5] VGND 2f $ **FLOATING
C1456 tdc0.w_dly_sig_n[4] VGND 1.75f $ **FLOATING
C1457 tdc0.w_dly_sig[4] VGND 2.89f $ **FLOATING
C1458 tdc0.w_dly_sig_n[3] VGND 2.22f $ **FLOATING
C1459 tdc0.w_dly_sig_n[0] VGND 2.69f $ **FLOATING
C1460 tdc0.w_dly_sig[3] VGND 4.22f $ **FLOATING
C1461 a_23591_11305# VGND 0.581f $ **FLOATING
C1462 a_23662_11204# VGND 0.626f $ **FLOATING
C1463 a_23462_11049# VGND 1.43f $ **FLOATING
C1464 a_23455_11145# VGND 1.81f $ **FLOATING
C1465 a_23171_11159# VGND 0.609f $ **FLOATING
C1466 a_23075_11159# VGND 0.817f $ **FLOATING
C1467 tdc0.w_dly_sig_n[34] VGND 2.81f $ **FLOATING
C1468 a_21843_11305# VGND 0.581f $ **FLOATING
C1469 a_21914_11204# VGND 0.626f $ **FLOATING
C1470 a_21714_11049# VGND 1.43f $ **FLOATING
C1471 a_21707_11145# VGND 1.81f $ **FLOATING
C1472 a_21423_11159# VGND 0.609f $ **FLOATING
C1473 a_21327_11159# VGND 0.817f $ **FLOATING
C1474 tdc0.w_dly_sig[33] VGND 3.51f $ **FLOATING
C1475 a_20003_11305# VGND 0.581f $ **FLOATING
C1476 a_20074_11204# VGND 0.626f $ **FLOATING
C1477 a_19874_11049# VGND 1.43f $ **FLOATING
C1478 a_19867_11145# VGND 1.81f $ **FLOATING
C1479 a_19583_11159# VGND 0.609f $ **FLOATING
C1480 a_19487_11159# VGND 0.817f $ **FLOATING
C1481 a_17937_10927# VGND 1.44f $ **FLOATING
C1482 tdc0.o_result[2] VGND 2.7f $ **FLOATING
C1483 _110_ VGND 1.96f $ **FLOATING
C1484 _094_ VGND 0.854f $ **FLOATING
C1485 a_16679_10927# VGND 0.972f $ **FLOATING
C1486 _008_ VGND 13.2f $ **FLOATING
C1487 tdc0.o_result[146] VGND 7.75f $ **FLOATING
C1488 a_16205_10901# VGND 0.713f $ **FLOATING
C1489 a_15059_10927# VGND 0.609f $ **FLOATING
C1490 a_15227_10901# VGND 0.817f $ **FLOATING
C1491 a_14634_10927# VGND 0.626f $ **FLOATING
C1492 a_14802_10901# VGND 0.581f $ **FLOATING
C1493 a_14361_10933# VGND 1.43f $ **FLOATING
C1494 a_14195_10933# VGND 1.81f $ **FLOATING
C1495 tdc0.w_dly_sig_n[75] VGND 1.72f $ **FLOATING
C1496 tdc0.w_dly_sig_n[76] VGND 1.82f $ **FLOATING
C1497 tdc0.w_dly_sig[77] VGND 4.02f $ **FLOATING
C1498 tdc0.w_dly_sig_n[78] VGND 1.91f $ **FLOATING
C1499 a_8491_10927# VGND 0.804f $ **FLOATING
C1500 tdc0.o_result[79] VGND 0.818f $ **FLOATING
C1501 tdc0.o_result[135] VGND 2.33f $ **FLOATING
C1502 a_7883_10927# VGND 0.609f $ **FLOATING
C1503 a_8051_10901# VGND 0.817f $ **FLOATING
C1504 a_7458_10927# VGND 0.626f $ **FLOATING
C1505 a_7626_10901# VGND 0.581f $ **FLOATING
C1506 a_7185_10933# VGND 1.43f $ **FLOATING
C1507 a_7019_10933# VGND 1.81f $ **FLOATING
C1508 a_5823_10927# VGND 0.972f $ **FLOATING
C1509 tdc0.o_result[116] VGND 1.12f $ **FLOATING
C1510 _131_ VGND 0.894f $ **FLOATING
C1511 tdc0.o_result[132] VGND 1.73f $ **FLOATING
C1512 _027_ VGND 5.05f $ **FLOATING
C1513 a_5115_11159# VGND 0.804f $ **FLOATING
C1514 a_4203_10927# VGND 0.609f $ **FLOATING
C1515 a_4371_10901# VGND 0.817f $ **FLOATING
C1516 a_3778_10927# VGND 0.626f $ **FLOATING
C1517 a_3946_10901# VGND 0.581f $ **FLOATING
C1518 a_3505_10933# VGND 1.43f $ **FLOATING
C1519 tdc0.w_dly_sig[117] VGND 3.51f $ **FLOATING
C1520 a_3339_10933# VGND 1.81f $ **FLOATING
C1521 a_2179_10927# VGND 0.609f $ **FLOATING
C1522 a_2347_10901# VGND 0.817f $ **FLOATING
C1523 a_1754_10927# VGND 0.626f $ **FLOATING
C1524 a_1922_10901# VGND 0.581f $ **FLOATING
C1525 a_1481_10933# VGND 1.43f $ **FLOATING
C1526 a_1315_10933# VGND 1.81f $ **FLOATING
C1527 a_30541_11471# VGND 0.23f $ **FLOATING
C1528 tdc0.w_dly_sig_n[7] VGND 3.2f $ **FLOATING
C1529 a_30123_11471# VGND 0.581f $ **FLOATING
C1530 a_30194_11445# VGND 0.626f $ **FLOATING
C1531 a_29987_11445# VGND 1.81f $ **FLOATING
C1532 a_29994_11745# VGND 1.43f $ **FLOATING
C1533 a_29703_11445# VGND 0.609f $ **FLOATING
C1534 a_29607_11623# VGND 0.817f $ **FLOATING
C1535 a_27137_11471# VGND 0.23f $ **FLOATING
C1536 a_20359_11471# VGND 0.594f $ **FLOATING
C1537 a_18703_11471# VGND 0.594f $ **FLOATING
C1538 tdc0.w_dly_sig[5] VGND 3.2f $ **FLOATING
C1539 a_26719_11471# VGND 0.581f $ **FLOATING
C1540 a_26790_11445# VGND 0.626f $ **FLOATING
C1541 a_26583_11445# VGND 1.81f $ **FLOATING
C1542 a_26590_11745# VGND 1.43f $ **FLOATING
C1543 a_26299_11445# VGND 0.609f $ **FLOATING
C1544 a_26203_11623# VGND 0.817f $ **FLOATING
C1545 a_25665_11471# VGND 0.23f $ **FLOATING
C1546 a_24170_11721# VGND 0.333f $ **FLOATING
C1547 _015_ VGND 3.17f $ **FLOATING
C1548 a_21071_11721# VGND 0.399f $ **FLOATING
C1549 a_20609_11721# VGND 0.384f $ **FLOATING
C1550 a_20359_11721# VGND 0.388f $ **FLOATING
C1551 a_19415_11721# VGND 0.399f $ **FLOATING
C1552 a_18953_11721# VGND 0.384f $ **FLOATING
C1553 a_18703_11721# VGND 0.388f $ **FLOATING
C1554 _137_ VGND 3.66f $ **FLOATING
C1555 _145_ VGND 3.62f $ **FLOATING
C1556 _037_ VGND 1.59f $ **FLOATING
C1557 _046_ VGND 3.92f $ **FLOATING
C1558 a_14878_11721# VGND 0.333f $ **FLOATING
C1559 _093_ VGND 2.28f $ **FLOATING
C1560 a_13633_11721# VGND 0.206f $ **FLOATING
C1561 a_12341_11471# VGND 0.23f $ **FLOATING
C1562 tdc0.w_dly_sig[1] VGND 2.91f $ **FLOATING
C1563 a_25247_11471# VGND 0.581f $ **FLOATING
C1564 a_25318_11445# VGND 0.626f $ **FLOATING
C1565 a_25111_11445# VGND 1.81f $ **FLOATING
C1566 a_25118_11745# VGND 1.43f $ **FLOATING
C1567 a_24827_11445# VGND 0.609f $ **FLOATING
C1568 a_24731_11623# VGND 0.817f $ **FLOATING
C1569 tdc0.o_result[8] VGND 3.09f $ **FLOATING
C1570 a_24013_11445# VGND 0.723f $ **FLOATING
C1571 tdc0.w_dly_sig_n[35] VGND 1.9f $ **FLOATING
C1572 tdc0.w_dly_sig[35] VGND 3.26f $ **FLOATING
C1573 tdc0.w_dly_sig[34] VGND 3.77f $ **FLOATING
C1574 a_20881_11721# VGND 1.44f $ **FLOATING
C1575 tdc0.o_result[0] VGND 2.41f $ **FLOATING
C1576 _063_ VGND 2.41f $ **FLOATING
C1577 _016_ VGND 1.16f $ **FLOATING
C1578 a_19225_11721# VGND 1.44f $ **FLOATING
C1579 tdc0.o_result[4] VGND 3.75f $ **FLOATING
C1580 _150_ VGND 1.03f $ **FLOATING
C1581 _134_ VGND 2.23f $ **FLOATING
C1582 _132_ VGND 6.72f $ **FLOATING
C1583 a_18059_11721# VGND 0.702f $ **FLOATING
C1584 a_16587_11721# VGND 0.702f $ **FLOATING
C1585 tdc0.o_result[34] VGND 3.74f $ **FLOATING
C1586 a_14721_11445# VGND 0.723f $ **FLOATING
C1587 a_13551_11721# VGND 0.804f $ **FLOATING
C1588 _085_ VGND 8.6f $ **FLOATING
C1589 tdc0.o_result[74] VGND 0.669f $ **FLOATING
C1590 a_12851_11837# VGND 0.609f $ **FLOATING
C1591 a_13019_11739# VGND 0.817f $ **FLOATING
C1592 a_12426_11837# VGND 0.626f $ **FLOATING
C1593 a_12594_11583# VGND 0.581f $ **FLOATING
C1594 a_12153_11471# VGND 1.43f $ **FLOATING
C1595 a_11987_11471# VGND 1.81f $ **FLOATING
C1596 tdc0.w_dly_sig[76] VGND 3.86f $ **FLOATING
C1597 tdc0.o_result[80] VGND 3.95f $ **FLOATING
C1598 a_10317_11471# VGND 0.23f $ **FLOATING
C1599 a_10827_11837# VGND 0.609f $ **FLOATING
C1600 a_10995_11739# VGND 0.817f $ **FLOATING
C1601 a_10402_11837# VGND 0.626f $ **FLOATING
C1602 a_10570_11583# VGND 0.581f $ **FLOATING
C1603 a_10129_11471# VGND 1.43f $ **FLOATING
C1604 a_9963_11471# VGND 1.81f $ **FLOATING
C1605 _092_ VGND 5.26f $ **FLOATING
C1606 a_7645_11721# VGND 0.214f $ **FLOATING
C1607 a_7561_11721# VGND 0.167f $ **FLOATING
C1608 a_5805_11721# VGND 0.214f $ **FLOATING
C1609 a_5721_11721# VGND 0.167f $ **FLOATING
C1610 a_3785_11471# VGND 0.23f $ **FLOATING
C1611 tdc0.w_dly_sig[78] VGND 3.95f $ **FLOATING
C1612 a_7479_11471# VGND 0.972f $ **FLOATING
C1613 tdc0.o_result[114] VGND 2.5f $ **FLOATING
C1614 _091_ VGND 3.77f $ **FLOATING
C1615 a_5639_11471# VGND 0.972f $ **FLOATING
C1616 tdc0.o_result[118] VGND 0.98f $ **FLOATING
C1617 _171_ VGND 1.01f $ **FLOATING
C1618 a_4295_11837# VGND 0.609f $ **FLOATING
C1619 a_4463_11739# VGND 0.817f $ **FLOATING
C1620 a_3870_11837# VGND 0.626f $ **FLOATING
C1621 a_4038_11583# VGND 0.581f $ **FLOATING
C1622 a_3597_11471# VGND 1.43f $ **FLOATING
C1623 a_3431_11471# VGND 1.81f $ **FLOATING
C1624 tdc0.o_result[108] VGND 1.77f $ **FLOATING
C1625 a_2037_11471# VGND 0.23f $ **FLOATING
C1626 a_2547_11837# VGND 0.609f $ **FLOATING
C1627 a_2715_11739# VGND 0.817f $ **FLOATING
C1628 a_2122_11837# VGND 0.626f $ **FLOATING
C1629 a_2290_11583# VGND 0.581f $ **FLOATING
C1630 a_1849_11471# VGND 1.43f $ **FLOATING
C1631 a_1683_11471# VGND 1.81f $ **FLOATING
C1632 tdc0.w_dly_sig[8] VGND 3.99f $ **FLOATING
C1633 a_29437_12393# VGND 0.23f $ **FLOATING
C1634 a_27873_12393# VGND 0.23f $ **FLOATING
C1635 a_24659_12015# VGND 0.399f $ **FLOATING
C1636 a_24197_12015# VGND 0.384f $ **FLOATING
C1637 a_23947_12015# VGND 0.388f $ **FLOATING
C1638 a_22917_12015# VGND 0.214f $ **FLOATING
C1639 a_22833_12015# VGND 0.167f $ **FLOATING
C1640 a_19967_12015# VGND 0.399f $ **FLOATING
C1641 a_19505_12015# VGND 0.384f $ **FLOATING
C1642 a_19255_12015# VGND 0.388f $ **FLOATING
C1643 a_17415_12015# VGND 0.333f $ **FLOATING
C1644 a_17076_12015# VGND 0.259f $ **FLOATING
C1645 a_15465_12015# VGND 0.214f $ **FLOATING
C1646 a_15381_12015# VGND 0.167f $ **FLOATING
C1647 a_23947_12335# VGND 0.594f $ **FLOATING
C1648 a_19255_12335# VGND 0.594f $ **FLOATING
C1649 _062_ VGND 0.892f $ **FLOATING
C1650 _156_ VGND 2.34f $ **FLOATING
C1651 a_6357_12015# VGND 0.214f $ **FLOATING
C1652 a_6273_12015# VGND 0.167f $ **FLOATING
C1653 a_7741_12015# VGND 0.23f $ **FLOATING
C1654 tdc0.w_dly_sig[129] VGND 3.42f $ **FLOATING
C1655 a_4613_12015# VGND 0.23f $ **FLOATING
C1656 tdc0.w_dly_sig[111] VGND 3.56f $ **FLOATING
C1657 tdc0.w_dly_sig_n[110] VGND 1.91f $ **FLOATING
C1658 a_29019_12393# VGND 0.581f $ **FLOATING
C1659 a_29090_12292# VGND 0.626f $ **FLOATING
C1660 a_28890_12137# VGND 1.43f $ **FLOATING
C1661 a_28883_12233# VGND 1.81f $ **FLOATING
C1662 a_28599_12247# VGND 0.609f $ **FLOATING
C1663 a_28503_12247# VGND 0.817f $ **FLOATING
C1664 tdc0.w_dly_sig[6] VGND 3.22f $ **FLOATING
C1665 a_27455_12393# VGND 0.581f $ **FLOATING
C1666 a_27526_12292# VGND 0.626f $ **FLOATING
C1667 a_27326_12137# VGND 1.43f $ **FLOATING
C1668 a_27319_12233# VGND 1.81f $ **FLOATING
C1669 a_27035_12247# VGND 0.609f $ **FLOATING
C1670 a_26939_12247# VGND 0.817f $ **FLOATING
C1671 a_24469_12015# VGND 1.44f $ **FLOATING
C1672 tdc0.o_result[5] VGND 1.57f $ **FLOATING
C1673 _170_ VGND 7.51f $ **FLOATING
C1674 _154_ VGND 1.05f $ **FLOATING
C1675 a_22751_12015# VGND 0.972f $ **FLOATING
C1676 _153_ VGND 7.91f $ **FLOATING
C1677 tdc0.w_dly_sig_n[36] VGND 2.47f $ **FLOATING
C1678 a_19777_12015# VGND 1.44f $ **FLOATING
C1679 tdc0.o_result[6] VGND 4.28f $ **FLOATING
C1680 _190_ VGND 1.95f $ **FLOATING
C1681 _174_ VGND 2.53f $ **FLOATING
C1682 _172_ VGND 6.94f $ **FLOATING
C1683 a_17498_12015# VGND 0.723f $ **FLOATING
C1684 _010_ VGND 14.3f $ **FLOATING
C1685 tdc0.o_result[11] VGND 7.5f $ **FLOATING
C1686 _057_ VGND 4.48f $ **FLOATING
C1687 _061_ VGND 5.02f $ **FLOATING
C1688 a_16645_11989# VGND 0.672f $ **FLOATING
C1689 a_15299_12015# VGND 0.972f $ **FLOATING
C1690 tdc0.o_result[142] VGND 5.15f $ **FLOATING
C1691 a_14045_12353# VGND 0.713f $ **FLOATING
C1692 a_12999_12128# VGND 0.619f $ **FLOATING
C1693 tdc0.w_dly_sig[79] VGND 3.46f $ **FLOATING
C1694 tdc0.w_dly_sig_n[79] VGND 1.92f $ **FLOATING
C1695 a_8251_12015# VGND 0.609f $ **FLOATING
C1696 a_8419_11989# VGND 0.817f $ **FLOATING
C1697 a_7826_12015# VGND 0.626f $ **FLOATING
C1698 a_7994_11989# VGND 0.581f $ **FLOATING
C1699 a_7553_12021# VGND 1.43f $ **FLOATING
C1700 a_7387_12021# VGND 1.81f $ **FLOATING
C1701 a_6191_12015# VGND 0.972f $ **FLOATING
C1702 _023_ VGND 9.18f $ **FLOATING
C1703 tdc0.o_result[119] VGND 0.863f $ **FLOATING
C1704 _191_ VGND 2.22f $ **FLOATING
C1705 a_5123_12015# VGND 0.609f $ **FLOATING
C1706 a_5291_11989# VGND 0.817f $ **FLOATING
C1707 a_4698_12015# VGND 0.626f $ **FLOATING
C1708 a_4866_11989# VGND 0.581f $ **FLOATING
C1709 a_4425_12021# VGND 1.43f $ **FLOATING
C1710 a_4259_12021# VGND 1.81f $ **FLOATING
C1711 tdc0.w_dly_sig[119] VGND 3.51f $ **FLOATING
C1712 a_29729_12559# VGND 0.23f $ **FLOATING
C1713 a_30239_12925# VGND 0.609f $ **FLOATING
C1714 a_30407_12827# VGND 0.817f $ **FLOATING
C1715 a_29814_12925# VGND 0.626f $ **FLOATING
C1716 a_29982_12671# VGND 0.581f $ **FLOATING
C1717 a_29541_12559# VGND 1.43f $ **FLOATING
C1718 a_29375_12559# VGND 1.81f $ **FLOATING
C1719 tdc0.w_dly_sig[7] VGND 3.29f $ **FLOATING
C1720 tdc0.w_dly_sig_n[6] VGND 2.79f $ **FLOATING
C1721 a_26882_12559# VGND 1.98f $ **FLOATING
C1722 a_26309_12559# VGND 0.23f $ **FLOATING
C1723 tdc0.o_result[38] VGND 5.64f $ **FLOATING
C1724 a_20175_12559# VGND 0.594f $ **FLOATING
C1725 a_25891_12559# VGND 0.581f $ **FLOATING
C1726 a_25962_12533# VGND 0.626f $ **FLOATING
C1727 a_25755_12533# VGND 1.81f $ **FLOATING
C1728 a_25762_12833# VGND 1.43f $ **FLOATING
C1729 a_25471_12533# VGND 0.609f $ **FLOATING
C1730 a_25375_12711# VGND 0.817f $ **FLOATING
C1731 tdc0.w_dly_sig_n[37] VGND 1.75f $ **FLOATING
C1732 tdc0.w_dly_sig[36] VGND 3.78f $ **FLOATING
C1733 a_22813_12559# VGND 0.23f $ **FLOATING
C1734 tdc0.o_result[37] VGND 1.2f $ **FLOATING
C1735 a_20887_12809# VGND 0.399f $ **FLOATING
C1736 a_20425_12809# VGND 0.384f $ **FLOATING
C1737 a_20175_12809# VGND 0.388f $ **FLOATING
C1738 a_22395_12559# VGND 0.581f $ **FLOATING
C1739 a_22466_12533# VGND 0.626f $ **FLOATING
C1740 a_22259_12533# VGND 1.81f $ **FLOATING
C1741 a_22266_12833# VGND 1.43f $ **FLOATING
C1742 a_21975_12533# VGND 0.609f $ **FLOATING
C1743 a_21879_12711# VGND 0.817f $ **FLOATING
C1744 a_20697_12809# VGND 1.44f $ **FLOATING
C1745 tdc0.o_result[7] VGND 4.93f $ **FLOATING
C1746 _064_ VGND 12.3f $ **FLOATING
C1747 _192_ VGND 6.98f $ **FLOATING
C1748 a_19807_12559# VGND 0.648f $ **FLOATING
C1749 _210_ VGND 1.15f $ **FLOATING
C1750 _197_ VGND 3.86f $ **FLOATING
C1751 _205_ VGND 3.9f $ **FLOATING
C1752 a_17887_12809# VGND 0.167f $ **FLOATING
C1753 a_17685_12809# VGND 0.214f $ **FLOATING
C1754 _112_ VGND 2.19f $ **FLOATING
C1755 _059_ VGND 0.9f $ **FLOATING
C1756 tdc0.o_result[72] VGND 0.732f $ **FLOATING
C1757 a_15285_12559# VGND 0.23f $ **FLOATING
C1758 a_19255_12809# VGND 0.702f $ **FLOATING
C1759 a_18703_12559# VGND 0.698f $ **FLOATING
C1760 _002_ VGND 5.18f $ **FLOATING
C1761 _111_ VGND 0.805f $ **FLOATING
C1762 _072_ VGND 12.3f $ **FLOATING
C1763 a_17559_12711# VGND 0.972f $ **FLOATING
C1764 a_16495_12559# VGND 0.619f $ **FLOATING
C1765 a_15795_12925# VGND 0.609f $ **FLOATING
C1766 a_15963_12827# VGND 0.817f $ **FLOATING
C1767 a_15370_12925# VGND 0.626f $ **FLOATING
C1768 a_15538_12671# VGND 0.581f $ **FLOATING
C1769 a_15097_12559# VGND 1.43f $ **FLOATING
C1770 a_14931_12559# VGND 1.81f $ **FLOATING
C1771 _201_ VGND 3.26f $ **FLOATING
C1772 a_13552_12809# VGND 0.259f $ **FLOATING
C1773 tdc0.w_dly_sig_n[74] VGND 2.22f $ **FLOATING
C1774 _086_ VGND 2.19f $ **FLOATING
C1775 tdc0.o_result[81] VGND 0.888f $ **FLOATING
C1776 a_10225_12559# VGND 0.23f $ **FLOATING
C1777 a_13722_12559# VGND 0.672f $ **FLOATING
C1778 _199_ VGND 4.89f $ **FLOATING
C1779 _198_ VGND 0.818f $ **FLOATING
C1780 tdc0.o_result[127] VGND 3.16f $ **FLOATING
C1781 a_12999_12559# VGND 0.619f $ **FLOATING
C1782 a_11803_12559# VGND 0.619f $ **FLOATING
C1783 a_10735_12925# VGND 0.609f $ **FLOATING
C1784 a_10903_12827# VGND 0.817f $ **FLOATING
C1785 a_10310_12925# VGND 0.626f $ **FLOATING
C1786 a_10478_12671# VGND 0.581f $ **FLOATING
C1787 a_10037_12559# VGND 1.43f $ **FLOATING
C1788 a_9871_12559# VGND 1.81f $ **FLOATING
C1789 tdc0.w_dly_sig[128] VGND 4.12f $ **FLOATING
C1790 tdc0.o_result[107] VGND 7.14f $ **FLOATING
C1791 a_2037_12559# VGND 0.23f $ **FLOATING
C1792 tdc0.w_dly_sig_n[80] VGND 1.98f $ **FLOATING
C1793 tdc0.w_dly_sig[80] VGND 4.15f $ **FLOATING
C1794 a_6550_12559# VGND 1.98f $ **FLOATING
C1795 tdc0.w_dly_sig_n[127] VGND 2.77f $ **FLOATING
C1796 tdc0.w_dly_sig[120] VGND 3.75f $ **FLOATING
C1797 a_2547_12925# VGND 0.609f $ **FLOATING
C1798 a_2715_12827# VGND 0.817f $ **FLOATING
C1799 a_2122_12925# VGND 0.626f $ **FLOATING
C1800 a_2290_12671# VGND 0.581f $ **FLOATING
C1801 a_1849_12559# VGND 1.43f $ **FLOATING
C1802 a_1683_12559# VGND 1.81f $ **FLOATING
C1803 tdc0.w_dly_sig_n[109] VGND 2.17f $ **FLOATING
C1804 a_29437_13481# VGND 0.23f $ **FLOATING
C1805 tdc0.o_result[42] VGND 6.57f $ **FLOATING
C1806 a_27965_13481# VGND 0.23f $ **FLOATING
C1807 a_22461_13103# VGND 0.23f $ **FLOATING
C1808 a_17765_13103# VGND 0.214f $ **FLOATING
C1809 a_17681_13103# VGND 0.167f $ **FLOATING
C1810 a_16680_13103# VGND 0.259f $ **FLOATING
C1811 a_14104_13103# VGND 0.259f $ **FLOATING
C1812 a_13184_13103# VGND 0.259f $ **FLOATING
C1813 _029_ VGND 2.68f $ **FLOATING
C1814 _053_ VGND 1.55f $ **FLOATING
C1815 _121_ VGND 2.28f $ **FLOATING
C1816 _141_ VGND 3.34f $ **FLOATING
C1817 tdc0.o_result[122] VGND 7.35f $ **FLOATING
C1818 a_6177_13103# VGND 0.23f $ **FLOATING
C1819 a_2037_13103# VGND 0.23f $ **FLOATING
C1820 tdc0.w_dly_sig[110] VGND 5.71f $ **FLOATING
C1821 clknet_4_14_0_clk VGND 12.9f $ **FLOATING
C1822 a_29019_13481# VGND 0.581f $ **FLOATING
C1823 a_29090_13380# VGND 0.626f $ **FLOATING
C1824 a_28890_13225# VGND 1.43f $ **FLOATING
C1825 a_28883_13321# VGND 1.81f $ **FLOATING
C1826 a_28599_13335# VGND 0.609f $ **FLOATING
C1827 a_28503_13335# VGND 0.817f $ **FLOATING
C1828 a_27547_13481# VGND 0.581f $ **FLOATING
C1829 a_27618_13380# VGND 0.626f $ **FLOATING
C1830 a_27418_13225# VGND 1.43f $ **FLOATING
C1831 a_27411_13321# VGND 1.81f $ **FLOATING
C1832 a_27127_13335# VGND 0.609f $ **FLOATING
C1833 a_27031_13335# VGND 0.817f $ **FLOATING
C1834 a_25410_13103# VGND 1.98f $ **FLOATING
C1835 tdc0.w_dly_sig_n[38] VGND 2.28f $ **FLOATING
C1836 a_22971_13103# VGND 0.609f $ **FLOATING
C1837 a_23139_13077# VGND 0.817f $ **FLOATING
C1838 a_22546_13103# VGND 0.626f $ **FLOATING
C1839 a_22714_13077# VGND 0.581f $ **FLOATING
C1840 a_22273_13109# VGND 1.43f $ **FLOATING
C1841 tdc0.w_dly_sig[37] VGND 4.11f $ **FLOATING
C1842 a_22107_13109# VGND 1.81f $ **FLOATING
C1843 a_21313_13441# VGND 0.713f $ **FLOATING
C1844 a_19890_13103# VGND 1.98f $ **FLOATING
C1845 a_19289_13441# VGND 0.713f $ **FLOATING
C1846 a_18843_13335# VGND 0.619f $ **FLOATING
C1847 a_17599_13103# VGND 0.972f $ **FLOATING
C1848 tdc0.o_result[40] VGND 4.8f $ **FLOATING
C1849 _028_ VGND 5.68f $ **FLOATING
C1850 a_16850_13423# VGND 0.672f $ **FLOATING
C1851 _052_ VGND 7.45f $ **FLOATING
C1852 _047_ VGND 12.5f $ **FLOATING
C1853 a_14274_13423# VGND 0.672f $ **FLOATING
C1854 tdc0.o_result[139] VGND 4.52f $ **FLOATING
C1855 a_13354_13423# VGND 0.672f $ **FLOATING
C1856 _140_ VGND 3.02f $ **FLOATING
C1857 _138_ VGND 1.21f $ **FLOATING
C1858 tdc0.o_result[140] VGND 4.33f $ **FLOATING
C1859 _039_ VGND 13.9f $ **FLOATING
C1860 a_12254_13103# VGND 1.98f $ **FLOATING
C1861 a_11711_13216# VGND 0.619f $ **FLOATING
C1862 _076_ VGND 12.9f $ **FLOATING
C1863 tdc0.w_dly_sig_n[81] VGND 2.19f $ **FLOATING
C1864 a_7378_13103# VGND 1.98f $ **FLOATING
C1865 a_6687_13103# VGND 0.609f $ **FLOATING
C1866 a_6855_13077# VGND 0.817f $ **FLOATING
C1867 a_6262_13103# VGND 0.626f $ **FLOATING
C1868 a_6430_13077# VGND 0.581f $ **FLOATING
C1869 a_5989_13109# VGND 1.43f $ **FLOATING
C1870 a_5823_13109# VGND 1.81f $ **FLOATING
C1871 tdc0.w_dly_sig_n[120] VGND 2.37f $ **FLOATING
C1872 tdc0.w_dly_sig[121] VGND 4.37f $ **FLOATING
C1873 tdc0.w_dly_sig_n[121] VGND 2.05f $ **FLOATING
C1874 a_2547_13103# VGND 0.609f $ **FLOATING
C1875 a_2715_13077# VGND 0.817f $ **FLOATING
C1876 a_2122_13103# VGND 0.626f $ **FLOATING
C1877 a_2290_13077# VGND 0.581f $ **FLOATING
C1878 a_1849_13109# VGND 1.43f $ **FLOATING
C1879 tdc0.w_dly_sig[112] VGND 4.01f $ **FLOATING
C1880 a_1683_13109# VGND 1.81f $ **FLOATING
C1881 clknet_4_4_0_clk VGND 13.3f $ **FLOATING
C1882 tdc0.w_dly_sig[39] VGND 3.59f $ **FLOATING
C1883 tdc0.w_dly_sig_n[39] VGND 2f $ **FLOATING
C1884 tdc0.w_dly_sig[38] VGND 4.46f $ **FLOATING
C1885 a_25573_13647# VGND 0.23f $ **FLOATING
C1886 _187_ VGND 2.75f $ **FLOATING
C1887 a_23240_13897# VGND 0.259f $ **FLOATING
C1888 _149_ VGND 3.65f $ **FLOATING
C1889 _107_ VGND 3.58f $ **FLOATING
C1890 tdc0.o_result[43] VGND 5.62f $ **FLOATING
C1891 _011_ VGND 13.2f $ **FLOATING
C1892 _118_ VGND 3.39f $ **FLOATING
C1893 a_19652_13897# VGND 0.259f $ **FLOATING
C1894 _209_ VGND 1.11f $ **FLOATING
C1895 _049_ VGND 0.9f $ **FLOATING
C1896 _048_ VGND 1.1f $ **FLOATING
C1897 tdc0.o_result[111] VGND 6.41f $ **FLOATING
C1898 _173_ VGND 1.29f $ **FLOATING
C1899 a_14839_13897# VGND 0.333f $ **FLOATING
C1900 _120_ VGND 1.15f $ **FLOATING
C1901 _200_ VGND 1.02f $ **FLOATING
C1902 _034_ VGND 10.1f $ **FLOATING
C1903 tdc0.w_dly_sig[74] VGND 5.53f $ **FLOATING
C1904 _139_ VGND 1.11f $ **FLOATING
C1905 tdc0.w_dly_sig[75] VGND 4.27f $ **FLOATING
C1906 tdc0.o_result[82] VGND 3.18f $ **FLOATING
C1907 a_10225_13647# VGND 0.23f $ **FLOATING
C1908 a_25155_13647# VGND 0.581f $ **FLOATING
C1909 a_25226_13621# VGND 0.626f $ **FLOATING
C1910 a_25019_13621# VGND 1.81f $ **FLOATING
C1911 a_25026_13921# VGND 1.43f $ **FLOATING
C1912 a_24735_13621# VGND 0.609f $ **FLOATING
C1913 a_24639_13799# VGND 0.817f $ **FLOATING
C1914 a_23855_13647# VGND 0.619f $ **FLOATING
C1915 tdc0.o_result[36] VGND 0.863f $ **FLOATING
C1916 a_22809_13793# VGND 0.672f $ **FLOATING
C1917 a_21923_13647# VGND 0.619f $ **FLOATING
C1918 a_21523_13799# VGND 0.56f $ **FLOATING
C1919 a_20945_13675# VGND 0.713f $ **FLOATING
C1920 a_20499_13799# VGND 0.619f $ **FLOATING
C1921 a_20039_13799# VGND 0.619f $ **FLOATING
C1922 _004_ VGND 12.4f $ **FLOATING
C1923 tdc0.o_result[39] VGND 2.82f $ **FLOATING
C1924 _206_ VGND 2.21f $ **FLOATING
C1925 _207_ VGND 1.01f $ **FLOATING
C1926 _208_ VGND 0.786f $ **FLOATING
C1927 a_19221_13793# VGND 0.672f $ **FLOATING
C1928 a_18703_13647# VGND 0.619f $ **FLOATING
C1929 a_17187_13799# VGND 0.619f $ **FLOATING
C1930 a_16219_13647# VGND 0.619f $ **FLOATING
C1931 a_15575_13647# VGND 0.619f $ **FLOATING
C1932 a_14922_13897# VGND 0.723f $ **FLOATING
C1933 _020_ VGND 7.75f $ **FLOATING
C1934 a_14103_13647# VGND 0.619f $ **FLOATING
C1935 a_13643_13647# VGND 0.619f $ **FLOATING
C1936 a_12723_13647# VGND 0.619f $ **FLOATING
C1937 a_11812_13621# VGND 1.98f $ **FLOATING
C1938 a_10735_14013# VGND 0.609f $ **FLOATING
C1939 a_10903_13915# VGND 0.817f $ **FLOATING
C1940 a_10310_14013# VGND 0.626f $ **FLOATING
C1941 a_10478_13759# VGND 0.581f $ **FLOATING
C1942 a_10037_13647# VGND 1.43f $ **FLOATING
C1943 a_9871_13647# VGND 1.81f $ **FLOATING
C1944 tdc0.o_result[124] VGND 2.08f $ **FLOATING
C1945 a_8753_13647# VGND 0.23f $ **FLOATING
C1946 a_9263_14013# VGND 0.609f $ **FLOATING
C1947 a_9431_13915# VGND 0.817f $ **FLOATING
C1948 a_8838_14013# VGND 0.626f $ **FLOATING
C1949 a_9006_13759# VGND 0.581f $ **FLOATING
C1950 a_8565_13647# VGND 1.43f $ **FLOATING
C1951 a_8399_13647# VGND 1.81f $ **FLOATING
C1952 tdc0.w_dly_sig[127] VGND 4.78f $ **FLOATING
C1953 tdc0.o_result[106] VGND 6.33f $ **FLOATING
C1954 a_2037_13647# VGND 0.23f $ **FLOATING
C1955 tdc0.w_dly_sig_n[126] VGND 2.43f $ **FLOATING
C1956 tdc0.w_dly_sig_n[125] VGND 2.33f $ **FLOATING
C1957 tdc0.w_dly_sig[125] VGND 3.75f $ **FLOATING
C1958 tdc0.w_dly_sig[123] VGND 3.18f $ **FLOATING
C1959 tdc0.w_dly_sig_n[122] VGND 2.21f $ **FLOATING
C1960 a_2547_14013# VGND 0.609f $ **FLOATING
C1961 a_2715_13915# VGND 0.817f $ **FLOATING
C1962 a_2122_14013# VGND 0.626f $ **FLOATING
C1963 a_2290_13759# VGND 0.581f $ **FLOATING
C1964 a_1849_13647# VGND 1.43f $ **FLOATING
C1965 a_1683_13647# VGND 1.81f $ **FLOATING
C1966 tdc0.w_dly_sig_n[108] VGND 1.88f $ **FLOATING
C1967 a_29913_14191# VGND 0.23f $ **FLOATING
C1968 a_24113_14191# VGND 0.214f $ **FLOATING
C1969 a_24029_14191# VGND 0.167f $ **FLOATING
C1970 _127_ VGND 2.94f $ **FLOATING
C1971 _152_ VGND 1.82f $ **FLOATING
C1972 _146_ VGND 0.85f $ **FLOATING
C1973 _147_ VGND 0.925f $ **FLOATING
C1974 _148_ VGND 1.01f $ **FLOATING
C1975 a_19885_14191# VGND 0.23f $ **FLOATING
C1976 tdc0.o_result[70] VGND 2.25f $ **FLOATING
C1977 a_16941_14191# VGND 0.23f $ **FLOATING
C1978 _119_ VGND 1.29f $ **FLOATING
C1979 tdc0.w_dly_sig_n[73] VGND 2.78f $ **FLOATING
C1980 tdc0.o_result[84] VGND 1.33f $ **FLOATING
C1981 a_11329_14191# VGND 0.23f $ **FLOATING
C1982 a_6913_14191# VGND 0.23f $ **FLOATING
C1983 tdc0.o_result[105] VGND 7.05f $ **FLOATING
C1984 a_3141_14191# VGND 0.23f $ **FLOATING
C1985 tdc0.w_dly_sig[109] VGND 3.52f $ **FLOATING
C1986 tdc0.w_dly_sig[108] VGND 3.54f $ **FLOATING
C1987 a_30423_14191# VGND 0.609f $ **FLOATING
C1988 a_30591_14165# VGND 0.817f $ **FLOATING
C1989 a_29998_14191# VGND 0.626f $ **FLOATING
C1990 a_30166_14165# VGND 0.581f $ **FLOATING
C1991 a_29725_14197# VGND 1.43f $ **FLOATING
C1992 a_29559_14197# VGND 1.81f $ **FLOATING
C1993 tdc0.w_dly_sig[43] VGND 3.23f $ **FLOATING
C1994 tdc0.w_dly_sig_n[42] VGND 2.05f $ **FLOATING
C1995 tdc0.w_dly_sig[41] VGND 2.97f $ **FLOATING
C1996 tdc0.w_dly_sig_n[41] VGND 1.95f $ **FLOATING
C1997 tdc0.w_dly_sig_n[40] VGND 2.08f $ **FLOATING
C1998 tdc0.w_dly_sig[40] VGND 3.42f $ **FLOATING
C1999 a_24731_14423# VGND 0.619f $ **FLOATING
C2000 a_23947_14191# VGND 0.972f $ **FLOATING
C2001 tdc0.o_result[44] VGND 4.12f $ **FLOATING
C2002 _012_ VGND 16.5f $ **FLOATING
C2003 a_23351_14423# VGND 0.619f $ **FLOATING
C2004 _003_ VGND 8.66f $ **FLOATING
C2005 _035_ VGND 20f $ **FLOATING
C2006 a_22891_14423# VGND 0.619f $ **FLOATING
C2007 a_22291_14304# VGND 0.619f $ **FLOATING
C2008 _058_ VGND 13f $ **FLOATING
C2009 _001_ VGND 15.2f $ **FLOATING
C2010 tdc0.o_result[68] VGND 1.4f $ **FLOATING
C2011 clknet_0_clk VGND 34.2f $ **FLOATING
C2012 a_21380_14165# VGND 1.98f $ **FLOATING
C2013 a_20395_14191# VGND 0.609f $ **FLOATING
C2014 a_20563_14165# VGND 0.817f $ **FLOATING
C2015 a_19970_14191# VGND 0.626f $ **FLOATING
C2016 a_20138_14165# VGND 0.581f $ **FLOATING
C2017 a_19697_14197# VGND 1.43f $ **FLOATING
C2018 a_19531_14197# VGND 1.81f $ **FLOATING
C2019 a_17451_14191# VGND 0.609f $ **FLOATING
C2020 a_17619_14165# VGND 0.817f $ **FLOATING
C2021 a_17026_14191# VGND 0.626f $ **FLOATING
C2022 a_17194_14165# VGND 0.581f $ **FLOATING
C2023 a_16753_14197# VGND 1.43f $ **FLOATING
C2024 a_16587_14197# VGND 1.81f $ **FLOATING
C2025 tdc0.w_dly_sig_n[72] VGND 2.23f $ **FLOATING
C2026 a_13735_14304# VGND 0.619f $ **FLOATING
C2027 _054_ VGND 17.4f $ **FLOATING
C2028 _022_ VGND 11.7f $ **FLOATING
C2029 tdc0.o_result[123] VGND 3.11f $ **FLOATING
C2030 tdc0.w_dly_sig[73] VGND 5f $ **FLOATING
C2031 a_11839_14191# VGND 0.609f $ **FLOATING
C2032 a_12007_14165# VGND 0.817f $ **FLOATING
C2033 a_11414_14191# VGND 0.626f $ **FLOATING
C2034 a_11582_14165# VGND 0.581f $ **FLOATING
C2035 a_11141_14197# VGND 1.43f $ **FLOATING
C2036 a_10975_14197# VGND 1.81f $ **FLOATING
C2037 tdc0.w_dly_sig_n[82] VGND 1.75f $ **FLOATING
C2038 tdc0.w_dly_sig[81] VGND 3.59f $ **FLOATING
C2039 tdc0.w_dly_sig[82] VGND 3.14f $ **FLOATING
C2040 a_7423_14191# VGND 0.609f $ **FLOATING
C2041 a_7591_14165# VGND 0.817f $ **FLOATING
C2042 a_6998_14191# VGND 0.626f $ **FLOATING
C2043 a_7166_14165# VGND 0.581f $ **FLOATING
C2044 a_6725_14197# VGND 1.43f $ **FLOATING
C2045 a_6559_14197# VGND 1.81f $ **FLOATING
C2046 tdc0.w_dly_sig_n[124] VGND 2.09f $ **FLOATING
C2047 tdc0.w_dly_sig[124] VGND 3.53f $ **FLOATING
C2048 tdc0.w_dly_sig_n[123] VGND 2.37f $ **FLOATING
C2049 a_3651_14191# VGND 0.609f $ **FLOATING
C2050 a_3819_14165# VGND 0.817f $ **FLOATING
C2051 a_3226_14191# VGND 0.626f $ **FLOATING
C2052 a_3394_14165# VGND 0.581f $ **FLOATING
C2053 a_2953_14197# VGND 1.43f $ **FLOATING
C2054 a_2787_14197# VGND 1.81f $ **FLOATING
C2055 tdc0.w_dly_sig_n[107] VGND 1.74f $ **FLOATING
C2056 tdc0.w_dly_sig[44] VGND 3.47f $ **FLOATING
C2057 tdc0.w_dly_sig_n[43] VGND 2.28f $ **FLOATING
C2058 tdc0.w_dly_sig_n[44] VGND 2.18f $ **FLOATING
C2059 a_26217_14735# VGND 0.23f $ **FLOATING
C2060 _194_ VGND 3.46f $ **FLOATING
C2061 a_24021_14985# VGND 0.214f $ **FLOATING
C2062 a_23937_14985# VGND 0.167f $ **FLOATING
C2063 tdc0.o_result[66] VGND 1.21f $ **FLOATING
C2064 a_21081_14735# VGND 0.23f $ **FLOATING
C2065 tdc0.w_dly_sig[42] VGND 3.15f $ **FLOATING
C2066 a_25799_14735# VGND 0.581f $ **FLOATING
C2067 a_25870_14709# VGND 0.626f $ **FLOATING
C2068 a_25663_14709# VGND 1.81f $ **FLOATING
C2069 a_25670_15009# VGND 1.43f $ **FLOATING
C2070 a_25379_14709# VGND 0.609f $ **FLOATING
C2071 a_25283_14887# VGND 0.817f $ **FLOATING
C2072 a_23855_14735# VGND 0.972f $ **FLOATING
C2073 _193_ VGND 4.86f $ **FLOATING
C2074 a_21591_15101# VGND 0.609f $ **FLOATING
C2075 a_21759_15003# VGND 0.817f $ **FLOATING
C2076 a_21166_15101# VGND 0.626f $ **FLOATING
C2077 a_21334_14847# VGND 0.581f $ **FLOATING
C2078 a_20893_14735# VGND 1.43f $ **FLOATING
C2079 a_20727_14735# VGND 1.81f $ **FLOATING
C2080 a_18785_14985# VGND 0.206f $ **FLOATING
C2081 _151_ VGND 3.41f $ **FLOATING
C2082 a_17773_14985# VGND 0.206f $ **FLOATING
C2083 a_16573_14735# VGND 0.23f $ **FLOATING
C2084 a_18703_14985# VGND 0.804f $ **FLOATING
C2085 _055_ VGND 7.91f $ **FLOATING
C2086 a_17691_14985# VGND 0.804f $ **FLOATING
C2087 _068_ VGND 7.62f $ **FLOATING
C2088 tdc0.o_result[69] VGND 0.76f $ **FLOATING
C2089 _065_ VGND 9.23f $ **FLOATING
C2090 a_17083_15101# VGND 0.609f $ **FLOATING
C2091 a_17251_15003# VGND 0.817f $ **FLOATING
C2092 a_16658_15101# VGND 0.626f $ **FLOATING
C2093 a_16826_14847# VGND 0.581f $ **FLOATING
C2094 a_16385_14735# VGND 1.43f $ **FLOATING
C2095 a_16219_14735# VGND 1.81f $ **FLOATING
C2096 tdc0.w_dly_sig[71] VGND 4.27f $ **FLOATING
C2097 tdc0.w_dly_sig_n[71] VGND 2.03f $ **FLOATING
C2098 tdc0.o_result[71] VGND 1.25f $ **FLOATING
C2099 a_12341_14735# VGND 0.23f $ **FLOATING
C2100 a_12851_15101# VGND 0.609f $ **FLOATING
C2101 a_13019_15003# VGND 0.817f $ **FLOATING
C2102 a_12426_15101# VGND 0.626f $ **FLOATING
C2103 a_12594_14847# VGND 0.581f $ **FLOATING
C2104 a_12153_14735# VGND 1.43f $ **FLOATING
C2105 tdc0.w_dly_sig[72] VGND 3.86f $ **FLOATING
C2106 a_11987_14735# VGND 1.81f $ **FLOATING
C2107 clknet_4_6_0_clk VGND 12.4f $ **FLOATING
C2108 tdc0.o_result[83] VGND 2.43f $ **FLOATING
C2109 a_10409_14735# VGND 0.23f $ **FLOATING
C2110 a_10919_15101# VGND 0.609f $ **FLOATING
C2111 a_11087_15003# VGND 0.817f $ **FLOATING
C2112 a_10494_15101# VGND 0.626f $ **FLOATING
C2113 a_10662_14847# VGND 0.581f $ **FLOATING
C2114 a_10221_14735# VGND 1.43f $ **FLOATING
C2115 a_10055_14735# VGND 1.81f $ **FLOATING
C2116 tdc0.o_result[125] VGND 4.86f $ **FLOATING
C2117 a_7189_14735# VGND 0.23f $ **FLOATING
C2118 tdc0.w_dly_sig[83] VGND 3f $ **FLOATING
C2119 a_7699_15101# VGND 0.609f $ **FLOATING
C2120 a_7867_15003# VGND 0.817f $ **FLOATING
C2121 a_7274_15101# VGND 0.626f $ **FLOATING
C2122 a_7442_14847# VGND 0.581f $ **FLOATING
C2123 a_7001_14735# VGND 1.43f $ **FLOATING
C2124 tdc0.w_dly_sig[126] VGND 4.22f $ **FLOATING
C2125 a_6835_14735# VGND 1.81f $ **FLOATING
C2126 tdc0.o_result[121] VGND 6.24f $ **FLOATING
C2127 a_4981_14735# VGND 0.23f $ **FLOATING
C2128 a_5491_15101# VGND 0.609f $ **FLOATING
C2129 a_5659_15003# VGND 0.817f $ **FLOATING
C2130 a_5066_15101# VGND 0.626f $ **FLOATING
C2131 a_5234_14847# VGND 0.581f $ **FLOATING
C2132 a_4793_14735# VGND 1.43f $ **FLOATING
C2133 tdc0.w_dly_sig[122] VGND 3.24f $ **FLOATING
C2134 a_4627_14735# VGND 1.81f $ **FLOATING
C2135 tdc0.w_dly_sig[107] VGND 3.08f $ **FLOATING
C2136 tdc0.o_result[45] VGND 4.32f $ **FLOATING
C2137 a_29913_15279# VGND 0.23f $ **FLOATING
C2138 a_27413_15657# VGND 0.23f $ **FLOATING
C2139 a_24511_15279# VGND 0.167f $ **FLOATING
C2140 a_24309_15279# VGND 0.214f $ **FLOATING
C2141 tdc0.o_result[47] VGND 1.8f $ **FLOATING
C2142 _067_ VGND 3.1f $ **FLOATING
C2143 tdc0.o_result[63] VGND 1.08f $ **FLOATING
C2144 a_22277_15279# VGND 0.23f $ **FLOATING
C2145 tdc0.o_result[65] VGND 3.02f $ **FLOATING
C2146 a_19701_15279# VGND 0.23f $ **FLOATING
C2147 tdc0.w_dly_sig[69] VGND 4.82f $ **FLOATING
C2148 tdc0.w_dly_sig_n[69] VGND 2.02f $ **FLOATING
C2149 tdc0.w_dly_sig_n[70] VGND 2.51f $ **FLOATING
C2150 tdc0.o_result[86] VGND 1.32f $ **FLOATING
C2151 a_13997_15279# VGND 0.23f $ **FLOATING
C2152 tdc0.o_result[85] VGND 1.95f $ **FLOATING
C2153 a_11881_15279# VGND 0.23f $ **FLOATING
C2154 tdc0.o_result[101] VGND 8.81f $ **FLOATING
C2155 a_6821_15279# VGND 0.23f $ **FLOATING
C2156 tdc0.o_result[102] VGND 2.29f $ **FLOATING
C2157 a_4521_15279# VGND 0.23f $ **FLOATING
C2158 tdc0.o_result[104] VGND 7.09f $ **FLOATING
C2159 a_3049_15279# VGND 0.23f $ **FLOATING
C2160 tdc0.w_dly_sig[106] VGND 2.91f $ **FLOATING
C2161 tdc0.w_dly_sig_n[106] VGND 2.22f $ **FLOATING
C2162 a_30423_15279# VGND 0.609f $ **FLOATING
C2163 a_30591_15253# VGND 0.817f $ **FLOATING
C2164 a_29998_15279# VGND 0.626f $ **FLOATING
C2165 a_30166_15253# VGND 0.581f $ **FLOATING
C2166 a_29725_15285# VGND 1.43f $ **FLOATING
C2167 a_29559_15285# VGND 1.81f $ **FLOATING
C2168 tdc0.w_dly_sig[45] VGND 3.14f $ **FLOATING
C2169 tdc0.w_dly_sig_n[46] VGND 2.09f $ **FLOATING
C2170 a_26995_15657# VGND 0.581f $ **FLOATING
C2171 a_27066_15556# VGND 0.626f $ **FLOATING
C2172 a_26866_15401# VGND 1.43f $ **FLOATING
C2173 a_26859_15497# VGND 1.81f $ **FLOATING
C2174 a_26575_15511# VGND 0.609f $ **FLOATING
C2175 a_26479_15511# VGND 0.817f $ **FLOATING
C2176 _066_ VGND 3.14f $ **FLOATING
C2177 _014_ VGND 9.62f $ **FLOATING
C2178 tdc0.o_result[41] VGND 1.18f $ **FLOATING
C2179 _017_ VGND 12.5f $ **FLOATING
C2180 a_24183_15511# VGND 0.972f $ **FLOATING
C2181 a_22787_15279# VGND 0.609f $ **FLOATING
C2182 a_22955_15253# VGND 0.817f $ **FLOATING
C2183 a_22362_15279# VGND 0.626f $ **FLOATING
C2184 a_22530_15253# VGND 0.581f $ **FLOATING
C2185 a_22089_15285# VGND 1.43f $ **FLOATING
C2186 a_21923_15285# VGND 1.81f $ **FLOATING
C2187 a_20211_15279# VGND 0.609f $ **FLOATING
C2188 a_20379_15253# VGND 0.817f $ **FLOATING
C2189 a_19786_15279# VGND 0.626f $ **FLOATING
C2190 a_19954_15253# VGND 0.581f $ **FLOATING
C2191 a_19513_15285# VGND 1.43f $ **FLOATING
C2192 a_19347_15285# VGND 1.81f $ **FLOATING
C2193 tdc0.w_dly_sig[67] VGND 3.61f $ **FLOATING
C2194 tdc0.w_dly_sig_n[68] VGND 1.72f $ **FLOATING
C2195 tdc0.w_dly_sig[70] VGND 3.7f $ **FLOATING
C2196 a_14507_15279# VGND 0.609f $ **FLOATING
C2197 a_14675_15253# VGND 0.817f $ **FLOATING
C2198 a_14082_15279# VGND 0.626f $ **FLOATING
C2199 a_14250_15253# VGND 0.581f $ **FLOATING
C2200 a_13809_15285# VGND 1.43f $ **FLOATING
C2201 a_13643_15285# VGND 1.81f $ **FLOATING
C2202 a_12391_15279# VGND 0.609f $ **FLOATING
C2203 a_12559_15253# VGND 0.817f $ **FLOATING
C2204 a_11966_15279# VGND 0.626f $ **FLOATING
C2205 a_12134_15253# VGND 0.581f $ **FLOATING
C2206 a_11693_15285# VGND 1.43f $ **FLOATING
C2207 a_11527_15285# VGND 1.81f $ **FLOATING
C2208 tdc0.w_dly_sig[84] VGND 2.77f $ **FLOATING
C2209 tdc0.w_dly_sig_n[83] VGND 2.17f $ **FLOATING
C2210 tdc0.w_dly_sig_n[84] VGND 2.22f $ **FLOATING
C2211 a_7331_15279# VGND 0.609f $ **FLOATING
C2212 a_7499_15253# VGND 0.817f $ **FLOATING
C2213 a_6906_15279# VGND 0.626f $ **FLOATING
C2214 a_7074_15253# VGND 0.581f $ **FLOATING
C2215 a_6633_15285# VGND 1.43f $ **FLOATING
C2216 a_6467_15285# VGND 1.81f $ **FLOATING
C2217 a_5031_15279# VGND 0.609f $ **FLOATING
C2218 a_5199_15253# VGND 0.817f $ **FLOATING
C2219 a_4606_15279# VGND 0.626f $ **FLOATING
C2220 a_4774_15253# VGND 0.581f $ **FLOATING
C2221 a_4333_15285# VGND 1.43f $ **FLOATING
C2222 a_4167_15285# VGND 1.81f $ **FLOATING
C2223 a_3559_15279# VGND 0.609f $ **FLOATING
C2224 a_3727_15253# VGND 0.817f $ **FLOATING
C2225 a_3134_15279# VGND 0.626f $ **FLOATING
C2226 a_3302_15253# VGND 0.581f $ **FLOATING
C2227 a_2861_15285# VGND 1.43f $ **FLOATING
C2228 a_2695_15285# VGND 1.81f $ **FLOATING
C2229 tdc0.w_dly_sig_n[105] VGND 2.19f $ **FLOATING
C2230 tdc0.w_dly_sig[46] VGND 3.51f $ **FLOATING
C2231 tdc0.w_dly_sig_n[45] VGND 2.61f $ **FLOATING
C2232 tdc0.w_dly_sig_n[47] VGND 1.81f $ **FLOATING
C2233 tdc0.w_dly_sig[48] VGND 2.9f $ **FLOATING
C2234 a_26309_15823# VGND 0.23f $ **FLOATING
C2235 tdc0.o_result[48] VGND 2.6f $ **FLOATING
C2236 a_25891_15823# VGND 0.581f $ **FLOATING
C2237 a_25962_15797# VGND 0.626f $ **FLOATING
C2238 a_25755_15797# VGND 1.81f $ **FLOATING
C2239 a_25762_16097# VGND 1.43f $ **FLOATING
C2240 a_25471_15797# VGND 0.609f $ **FLOATING
C2241 a_25375_15975# VGND 0.817f $ **FLOATING
C2242 a_24837_15823# VGND 0.23f $ **FLOATING
C2243 tdc0.o_result[49] VGND 1.1f $ **FLOATING
C2244 tdc0.o_result[62] VGND 1.89f $ **FLOATING
C2245 a_22461_15823# VGND 0.23f $ **FLOATING
C2246 a_24419_15823# VGND 0.581f $ **FLOATING
C2247 a_24490_15797# VGND 0.626f $ **FLOATING
C2248 a_24283_15797# VGND 1.81f $ **FLOATING
C2249 a_24290_16097# VGND 1.43f $ **FLOATING
C2250 a_23999_15797# VGND 0.609f $ **FLOATING
C2251 a_23903_15975# VGND 0.817f $ **FLOATING
C2252 a_22971_16189# VGND 0.609f $ **FLOATING
C2253 a_23139_16091# VGND 0.817f $ **FLOATING
C2254 a_22546_16189# VGND 0.626f $ **FLOATING
C2255 a_22714_15935# VGND 0.581f $ **FLOATING
C2256 a_22273_15823# VGND 1.43f $ **FLOATING
C2257 a_22107_15823# VGND 1.81f $ **FLOATING
C2258 tdc0.w_dly_sig_n[67] VGND 1.81f $ **FLOATING
C2259 tdc0.w_dly_sig_n[65] VGND 2.03f $ **FLOATING
C2260 tdc0.w_dly_sig[66] VGND 3.2f $ **FLOATING
C2261 tdc0.w_dly_sig_n[66] VGND 2.31f $ **FLOATING
C2262 a_17109_15823# VGND 0.23f $ **FLOATING
C2263 tdc0.o_result[64] VGND 2.14f $ **FLOATING
C2264 tdc0.o_result[67] VGND 3.93f $ **FLOATING
C2265 a_15009_15823# VGND 0.23f $ **FLOATING
C2266 a_16691_15823# VGND 0.581f $ **FLOATING
C2267 a_16762_15797# VGND 0.626f $ **FLOATING
C2268 a_16555_15797# VGND 1.81f $ **FLOATING
C2269 a_16562_16097# VGND 1.43f $ **FLOATING
C2270 a_16271_15797# VGND 0.609f $ **FLOATING
C2271 a_16175_15975# VGND 0.817f $ **FLOATING
C2272 a_15519_16189# VGND 0.609f $ **FLOATING
C2273 a_15687_16091# VGND 0.817f $ **FLOATING
C2274 a_15094_16189# VGND 0.626f $ **FLOATING
C2275 a_15262_15935# VGND 0.581f $ **FLOATING
C2276 a_14821_15823# VGND 1.43f $ **FLOATING
C2277 tdc0.w_dly_sig[68] VGND 4.02f $ **FLOATING
C2278 a_14655_15823# VGND 1.81f $ **FLOATING
C2279 tdc0.o_result[87] VGND 2.27f $ **FLOATING
C2280 a_12341_15823# VGND 0.23f $ **FLOATING
C2281 a_12851_16189# VGND 0.609f $ **FLOATING
C2282 a_13019_16091# VGND 0.817f $ **FLOATING
C2283 a_12426_16189# VGND 0.626f $ **FLOATING
C2284 a_12594_15935# VGND 0.581f $ **FLOATING
C2285 a_12153_15823# VGND 1.43f $ **FLOATING
C2286 a_11987_15823# VGND 1.81f $ **FLOATING
C2287 tdc0.o_result[99] VGND 5.56f $ **FLOATING
C2288 a_8753_15823# VGND 0.23f $ **FLOATING
C2289 tdc0.w_dly_sig[85] VGND 3.72f $ **FLOATING
C2290 tdc0.w_dly_sig_n[86] VGND 1.71f $ **FLOATING
C2291 a_9263_16189# VGND 0.609f $ **FLOATING
C2292 a_9431_16091# VGND 0.817f $ **FLOATING
C2293 a_8838_16189# VGND 0.626f $ **FLOATING
C2294 a_9006_15935# VGND 0.581f $ **FLOATING
C2295 a_8565_15823# VGND 1.43f $ **FLOATING
C2296 a_8399_15823# VGND 1.81f $ **FLOATING
C2297 tdc0.o_result[103] VGND 2.11f $ **FLOATING
C2298 a_5349_15823# VGND 0.23f $ **FLOATING
C2299 a_5859_16189# VGND 0.609f $ **FLOATING
C2300 a_6027_16091# VGND 0.817f $ **FLOATING
C2301 a_5434_16189# VGND 0.626f $ **FLOATING
C2302 a_5602_15935# VGND 0.581f $ **FLOATING
C2303 a_5161_15823# VGND 1.43f $ **FLOATING
C2304 a_4995_15823# VGND 1.81f $ **FLOATING
C2305 tdc0.w_dly_sig[105] VGND 3.18f $ **FLOATING
C2306 tdc0.w_dly_sig_n[103] VGND 1.72f $ **FLOATING
C2307 a_29621_16745# VGND 0.23f $ **FLOATING
C2308 tdc0.o_result[46] VGND 8.58f $ **FLOATING
C2309 tdc0.o_result[51] VGND 1.51f $ **FLOATING
C2310 a_23933_16367# VGND 0.23f $ **FLOATING
C2311 tdc0.w_dly_sig[64] VGND 3.61f $ **FLOATING
C2312 tdc0.w_dly_sig[65] VGND 4.61f $ **FLOATING
C2313 tdc0.o_result[60] VGND 1.89f $ **FLOATING
C2314 a_18137_16367# VGND 0.23f $ **FLOATING
C2315 tdc0.o_result[89] VGND 3.15f $ **FLOATING
C2316 a_13537_16367# VGND 0.23f $ **FLOATING
C2317 tdc0.w_dly_sig[86] VGND 3.64f $ **FLOATING
C2318 tdc0.o_result[97] VGND 5.49f $ **FLOATING
C2319 a_8385_16367# VGND 0.23f $ **FLOATING
C2320 tdc0.o_result[98] VGND 2.55f $ **FLOATING
C2321 a_6729_16367# VGND 0.23f $ **FLOATING
C2322 tdc0.w_dly_sig[103] VGND 3.46f $ **FLOATING
C2323 tdc0.w_dly_sig_n[102] VGND 1.79f $ **FLOATING
C2324 tdc0.w_dly_sig_n[104] VGND 2.1f $ **FLOATING
C2325 tdc0.w_dly_sig[47] VGND 3.09f $ **FLOATING
C2326 a_29203_16745# VGND 0.581f $ **FLOATING
C2327 a_29274_16644# VGND 0.626f $ **FLOATING
C2328 a_29074_16489# VGND 1.43f $ **FLOATING
C2329 a_29067_16585# VGND 1.81f $ **FLOATING
C2330 a_28783_16599# VGND 0.609f $ **FLOATING
C2331 a_28687_16599# VGND 0.817f $ **FLOATING
C2332 tdc0.w_dly_sig_n[48] VGND 2.5f $ **FLOATING
C2333 tdc0.w_dly_sig_n[49] VGND 1.84f $ **FLOATING
C2334 tdc0.w_dly_sig[49] VGND 3.83f $ **FLOATING
C2335 a_24443_16367# VGND 0.609f $ **FLOATING
C2336 a_24611_16341# VGND 0.817f $ **FLOATING
C2337 a_24018_16367# VGND 0.626f $ **FLOATING
C2338 a_24186_16341# VGND 0.581f $ **FLOATING
C2339 a_23745_16373# VGND 1.43f $ **FLOATING
C2340 a_23579_16373# VGND 1.81f $ **FLOATING
C2341 tdc0.w_dly_sig[63] VGND 3.61f $ **FLOATING
C2342 tdc0.w_dly_sig_n[64] VGND 2.04f $ **FLOATING
C2343 a_18647_16367# VGND 0.609f $ **FLOATING
C2344 a_18815_16341# VGND 0.817f $ **FLOATING
C2345 a_18222_16367# VGND 0.626f $ **FLOATING
C2346 a_18390_16341# VGND 0.581f $ **FLOATING
C2347 a_17949_16373# VGND 1.43f $ **FLOATING
C2348 a_17783_16373# VGND 1.81f $ **FLOATING
C2349 a_14047_16367# VGND 0.609f $ **FLOATING
C2350 a_14215_16341# VGND 0.817f $ **FLOATING
C2351 a_13622_16367# VGND 0.626f $ **FLOATING
C2352 a_13790_16341# VGND 0.581f $ **FLOATING
C2353 a_13349_16373# VGND 1.43f $ **FLOATING
C2354 a_13183_16373# VGND 1.81f $ **FLOATING
C2355 tdc0.w_dly_sig[87] VGND 4.48f $ **FLOATING
C2356 tdc0.w_dly_sig_n[87] VGND 1.95f $ **FLOATING
C2357 tdc0.w_dly_sig_n[85] VGND 2.45f $ **FLOATING
C2358 a_8895_16367# VGND 0.609f $ **FLOATING
C2359 a_9063_16341# VGND 0.817f $ **FLOATING
C2360 a_8470_16367# VGND 0.626f $ **FLOATING
C2361 a_8638_16341# VGND 0.581f $ **FLOATING
C2362 a_8197_16373# VGND 1.43f $ **FLOATING
C2363 a_8031_16373# VGND 1.81f $ **FLOATING
C2364 a_7239_16367# VGND 0.609f $ **FLOATING
C2365 a_7407_16341# VGND 0.817f $ **FLOATING
C2366 a_6814_16367# VGND 0.626f $ **FLOATING
C2367 a_6982_16341# VGND 0.581f $ **FLOATING
C2368 a_6541_16373# VGND 1.43f $ **FLOATING
C2369 a_6375_16373# VGND 1.81f $ **FLOATING
C2370 tdc0.w_dly_sig_n[100] VGND 1.79f $ **FLOATING
C2371 tdc0.w_dly_sig_n[101] VGND 1.76f $ **FLOATING
C2372 tdc0.w_dly_sig[102] VGND 4.21f $ **FLOATING
C2373 tdc0.w_dly_sig[104] VGND 4.41f $ **FLOATING
C2374 a_27321_16911# VGND 0.23f $ **FLOATING
C2375 tdc0.o_result[50] VGND 8.97f $ **FLOATING
C2376 tdc0.o_result[61] VGND 2.47f $ **FLOATING
C2377 a_22093_16911# VGND 0.23f $ **FLOATING
C2378 a_26903_16911# VGND 0.581f $ **FLOATING
C2379 a_26974_16885# VGND 0.626f $ **FLOATING
C2380 a_26767_16885# VGND 1.81f $ **FLOATING
C2381 a_26774_17185# VGND 1.43f $ **FLOATING
C2382 a_26483_16885# VGND 0.609f $ **FLOATING
C2383 a_26387_17063# VGND 0.817f $ **FLOATING
C2384 tdc0.w_dly_sig_n[50] VGND 1.94f $ **FLOATING
C2385 tdc0.w_dly_sig[50] VGND 3.88f $ **FLOATING
C2386 a_22603_17277# VGND 0.609f $ **FLOATING
C2387 a_22771_17179# VGND 0.817f $ **FLOATING
C2388 a_22178_17277# VGND 0.626f $ **FLOATING
C2389 a_22346_17023# VGND 0.581f $ **FLOATING
C2390 a_21905_16911# VGND 1.43f $ **FLOATING
C2391 a_21739_16911# VGND 1.81f $ **FLOATING
C2392 tdc0.w_dly_sig_n[63] VGND 1.89f $ **FLOATING
C2393 tdc0.w_dly_sig_n[62] VGND 2.26f $ **FLOATING
C2394 tdc0.w_dly_sig[62] VGND 2.47f $ **FLOATING
C2395 tdc0.w_dly_sig_n[61] VGND 2.23f $ **FLOATING
C2396 a_17477_16911# VGND 0.23f $ **FLOATING
C2397 tdc0.o_result[59] VGND 2.93f $ **FLOATING
C2398 tdc0.o_result[88] VGND 2.82f $ **FLOATING
C2399 a_15101_16911# VGND 0.23f $ **FLOATING
C2400 a_17059_16911# VGND 0.581f $ **FLOATING
C2401 a_17130_16885# VGND 0.626f $ **FLOATING
C2402 a_16923_16885# VGND 1.81f $ **FLOATING
C2403 a_16930_17185# VGND 1.43f $ **FLOATING
C2404 a_16639_16885# VGND 0.609f $ **FLOATING
C2405 a_16543_17063# VGND 0.817f $ **FLOATING
C2406 a_15611_17277# VGND 0.609f $ **FLOATING
C2407 a_15779_17179# VGND 0.817f $ **FLOATING
C2408 a_15186_17277# VGND 0.626f $ **FLOATING
C2409 a_15354_17023# VGND 0.581f $ **FLOATING
C2410 a_14913_16911# VGND 1.43f $ **FLOATING
C2411 a_14747_16911# VGND 1.81f $ **FLOATING
C2412 tdc0.o_result[95] VGND 5.67f $ **FLOATING
C2413 a_10041_16911# VGND 0.23f $ **FLOATING
C2414 tdc0.w_dly_sig_n[88] VGND 1.84f $ **FLOATING
C2415 tdc0.w_dly_sig[88] VGND 3.37f $ **FLOATING
C2416 a_10551_17277# VGND 0.609f $ **FLOATING
C2417 a_10719_17179# VGND 0.817f $ **FLOATING
C2418 a_10126_17277# VGND 0.626f $ **FLOATING
C2419 a_10294_17023# VGND 0.581f $ **FLOATING
C2420 a_9853_16911# VGND 1.43f $ **FLOATING
C2421 a_9687_16911# VGND 1.81f $ **FLOATING
C2422 tdc0.w_dly_sig[100] VGND 4.17f $ **FLOATING
C2423 tdc0.o_result[100] VGND 3.47f $ **FLOATING
C2424 a_4061_16911# VGND 0.23f $ **FLOATING
C2425 tdc0.w_dly_sig_n[99] VGND 1.72f $ **FLOATING
C2426 a_4571_17277# VGND 0.609f $ **FLOATING
C2427 a_4739_17179# VGND 0.817f $ **FLOATING
C2428 a_4146_17277# VGND 0.626f $ **FLOATING
C2429 a_4314_17023# VGND 0.581f $ **FLOATING
C2430 a_3873_16911# VGND 1.43f $ **FLOATING
C2431 tdc0.w_dly_sig[101] VGND 3.45f $ **FLOATING
C2432 a_3707_16911# VGND 1.81f $ **FLOATING
C2433 tt_um_hpretl_tt06_tdc_v1_8.HI VGND 0.415f $ **FLOATING
C2434 a_23733_17833# VGND 0.23f $ **FLOATING
C2435 tdc0.o_result[52] VGND 2.09f $ **FLOATING
C2436 a_22261_17833# VGND 0.23f $ **FLOATING
C2437 tdc0.o_result[54] VGND 4.3f $ **FLOATING
C2438 tdc0.w_dly_sig_n[60] VGND 2.17f $ **FLOATING
C2439 tdc0.w_dly_sig[61] VGND 3.72f $ **FLOATING
C2440 tdc0.w_dly_sig[60] VGND 3.97f $ **FLOATING
C2441 tdc0.o_result[58] VGND 4.68f $ **FLOATING
C2442 a_16757_17455# VGND 0.23f $ **FLOATING
C2443 tdc0.o_result[90] VGND 3.65f $ **FLOATING
C2444 a_13997_17455# VGND 0.23f $ **FLOATING
C2445 tdc0.o_result[96] VGND 5.08f $ **FLOATING
C2446 a_8661_17455# VGND 0.23f $ **FLOATING
C2447 tdc0.w_dly_sig_n[98] VGND 1.89f $ **FLOATING
C2448 tdc0.w_dly_sig[99] VGND 3.04f $ **FLOATING
C2449 tdc0.w_dly_sig[51] VGND 3.56f $ **FLOATING
C2450 tdc0.w_dly_sig_n[51] VGND 2.15f $ **FLOATING
C2451 tdc0.w_dly_sig[52] VGND 3.72f $ **FLOATING
C2452 a_23315_17833# VGND 0.581f $ **FLOATING
C2453 a_23386_17732# VGND 0.626f $ **FLOATING
C2454 a_23186_17577# VGND 1.43f $ **FLOATING
C2455 a_23179_17673# VGND 1.81f $ **FLOATING
C2456 a_22895_17687# VGND 0.609f $ **FLOATING
C2457 a_22799_17687# VGND 0.817f $ **FLOATING
C2458 a_21843_17833# VGND 0.581f $ **FLOATING
C2459 a_21914_17732# VGND 0.626f $ **FLOATING
C2460 a_21714_17577# VGND 1.43f $ **FLOATING
C2461 a_21707_17673# VGND 1.81f $ **FLOATING
C2462 a_21423_17687# VGND 0.609f $ **FLOATING
C2463 a_21327_17687# VGND 0.817f $ **FLOATING
C2464 tdc0.w_dly_sig_n[59] VGND 1.87f $ **FLOATING
C2465 a_17267_17455# VGND 0.609f $ **FLOATING
C2466 a_17435_17429# VGND 0.817f $ **FLOATING
C2467 a_16842_17455# VGND 0.626f $ **FLOATING
C2468 a_17010_17429# VGND 0.581f $ **FLOATING
C2469 a_16569_17461# VGND 1.43f $ **FLOATING
C2470 a_16403_17461# VGND 1.81f $ **FLOATING
C2471 a_14507_17455# VGND 0.609f $ **FLOATING
C2472 a_14675_17429# VGND 0.817f $ **FLOATING
C2473 a_14082_17455# VGND 0.626f $ **FLOATING
C2474 a_14250_17429# VGND 0.581f $ **FLOATING
C2475 a_13809_17461# VGND 1.43f $ **FLOATING
C2476 a_13643_17461# VGND 1.81f $ **FLOATING
C2477 tdc0.w_dly_sig[90] VGND 2.97f $ **FLOATING
C2478 tdc0.w_dly_sig[89] VGND 3.95f $ **FLOATING
C2479 tdc0.w_dly_sig_n[89] VGND 2.45f $ **FLOATING
C2480 a_9171_17455# VGND 0.609f $ **FLOATING
C2481 a_9339_17429# VGND 0.817f $ **FLOATING
C2482 a_8746_17455# VGND 0.626f $ **FLOATING
C2483 a_8914_17429# VGND 0.581f $ **FLOATING
C2484 a_8473_17461# VGND 1.43f $ **FLOATING
C2485 a_8307_17461# VGND 1.81f $ **FLOATING
C2486 clknet_4_5_0_clk VGND 19f $ **FLOATING
C2487 tdc0.w_dly_sig[59] VGND 3.57f $ **FLOATING
C2488 tdc0.o_result[57] VGND 2.11f $ **FLOATING
C2489 a_17493_17999# VGND 0.23f $ **FLOATING
C2490 tdc0.w_dly_sig_n[52] VGND 2.14f $ **FLOATING
C2491 tdc0.w_dly_sig_n[53] VGND 1.88f $ **FLOATING
C2492 tdc0.w_dly_sig[53] VGND 3.37f $ **FLOATING
C2493 tdc0.w_dly_sig[55] VGND 3.42f $ **FLOATING
C2494 tdc0.w_dly_sig_n[57] VGND 1.72f $ **FLOATING
C2495 a_18003_18365# VGND 0.609f $ **FLOATING
C2496 a_18171_18267# VGND 0.817f $ **FLOATING
C2497 a_17578_18365# VGND 0.626f $ **FLOATING
C2498 a_17746_18111# VGND 0.581f $ **FLOATING
C2499 a_17305_17999# VGND 1.43f $ **FLOATING
C2500 a_17139_17999# VGND 1.81f $ **FLOATING
C2501 tdc0.w_dly_sig_n[58] VGND 2.53f $ **FLOATING
C2502 tdc0.o_result[92] VGND 3.83f $ **FLOATING
C2503 a_14917_17999# VGND 0.23f $ **FLOATING
C2504 tdc0.w_dly_sig[58] VGND 3.82f $ **FLOATING
C2505 a_15427_18365# VGND 0.609f $ **FLOATING
C2506 a_15595_18267# VGND 0.817f $ **FLOATING
C2507 a_15002_18365# VGND 0.626f $ **FLOATING
C2508 a_15170_18111# VGND 0.581f $ **FLOATING
C2509 a_14729_17999# VGND 1.43f $ **FLOATING
C2510 a_14563_17999# VGND 1.81f $ **FLOATING
C2511 tdc0.o_result[94] VGND 3.88f $ **FLOATING
C2512 a_10317_17999# VGND 0.23f $ **FLOATING
C2513 tdc0.w_dly_sig_n[91] VGND 1.93f $ **FLOATING
C2514 tdc0.w_dly_sig_n[90] VGND 1.87f $ **FLOATING
C2515 tdc0.w_dly_sig[91] VGND 3.14f $ **FLOATING
C2516 tdc0.w_dly_sig_n[92] VGND 1.71f $ **FLOATING
C2517 a_10827_18365# VGND 0.609f $ **FLOATING
C2518 a_10995_18267# VGND 0.817f $ **FLOATING
C2519 a_10402_18365# VGND 0.626f $ **FLOATING
C2520 a_10570_18111# VGND 0.581f $ **FLOATING
C2521 a_10129_17999# VGND 1.43f $ **FLOATING
C2522 a_9963_17999# VGND 1.81f $ **FLOATING
C2523 tdc0.w_dly_sig[97] VGND 2.93f $ **FLOATING
C2524 tdc0.w_dly_sig_n[96] VGND 1.85f $ **FLOATING
C2525 tdc0.w_dly_sig[98] VGND 3.89f $ **FLOATING
C2526 tt_um_hpretl_tt06_tdc_v1_9.HI VGND 0.415f $ **FLOATING
C2527 tdc0.w_dly_sig[96] VGND 3.9f $ **FLOATING
C2528 tdc0.w_dly_sig_n[97] VGND 2.04f $ **FLOATING
C2529 tt_um_hpretl_tt06_tdc_v1_22.HI VGND 0.415f $ **FLOATING
C2530 tt_um_hpretl_tt06_tdc_v1_14.HI VGND 0.415f $ **FLOATING
C2531 tt_um_hpretl_tt06_tdc_v1_18.HI VGND 0.415f $ **FLOATING
C2532 tt_um_hpretl_tt06_tdc_v1_21.HI VGND 0.415f $ **FLOATING
C2533 a_24837_18921# VGND 0.23f $ **FLOATING
C2534 tdc0.o_result[53] VGND 2.35f $ **FLOATING
C2535 tdc0.w_dly_sig_n[54] VGND 1.99f $ **FLOATING
C2536 tdc0.o_result[55] VGND 2.81f $ **FLOATING
C2537 a_19333_18543# VGND 0.23f $ **FLOATING
C2538 tdc0.o_result[56] VGND 3.58f $ **FLOATING
C2539 a_16481_18543# VGND 0.23f $ **FLOATING
C2540 tdc0.o_result[91] VGND 4.69f $ **FLOATING
C2541 a_13997_18543# VGND 0.23f $ **FLOATING
C2542 tdc0.o_result[93] VGND 3.88f $ **FLOATING
C2543 a_11513_18543# VGND 0.23f $ **FLOATING
C2544 tdc0.w_dly_sig_n[95] VGND 1.91f $ **FLOATING
C2545 clknet_4_15_0_clk VGND 19.1f $ **FLOATING
C2546 a_24419_18921# VGND 0.581f $ **FLOATING
C2547 a_24490_18820# VGND 0.626f $ **FLOATING
C2548 a_24290_18665# VGND 1.43f $ **FLOATING
C2549 a_24283_18761# VGND 1.81f $ **FLOATING
C2550 a_23999_18775# VGND 0.609f $ **FLOATING
C2551 a_23903_18775# VGND 0.817f $ **FLOATING
C2552 tdc0.w_dly_sig[54] VGND 3.82f $ **FLOATING
C2553 tdc0.w_dly_sig_n[55] VGND 2.38f $ **FLOATING
C2554 tdc0.w_dly_sig_n[56] VGND 2f $ **FLOATING
C2555 a_19843_18543# VGND 0.609f $ **FLOATING
C2556 a_20011_18517# VGND 0.817f $ **FLOATING
C2557 a_19418_18543# VGND 0.626f $ **FLOATING
C2558 a_19586_18517# VGND 0.581f $ **FLOATING
C2559 a_19145_18549# VGND 1.43f $ **FLOATING
C2560 tdc0.w_dly_sig[56] VGND 4.45f $ **FLOATING
C2561 a_18979_18549# VGND 1.81f $ **FLOATING
C2562 clknet_4_12_0_clk VGND 10.1f $ **FLOATING
C2563 a_16991_18543# VGND 0.609f $ **FLOATING
C2564 a_17159_18517# VGND 0.817f $ **FLOATING
C2565 a_16566_18543# VGND 0.626f $ **FLOATING
C2566 a_16734_18517# VGND 0.581f $ **FLOATING
C2567 a_16293_18549# VGND 1.43f $ **FLOATING
C2568 tdc0.w_dly_sig[57] VGND 4.84f $ **FLOATING
C2569 a_16127_18549# VGND 1.81f $ **FLOATING
C2570 clknet_4_13_0_clk VGND 13.6f $ **FLOATING
C2571 a_14507_18543# VGND 0.609f $ **FLOATING
C2572 a_14675_18517# VGND 0.817f $ **FLOATING
C2573 a_14082_18543# VGND 0.626f $ **FLOATING
C2574 a_14250_18517# VGND 0.581f $ **FLOATING
C2575 a_13809_18549# VGND 1.43f $ **FLOATING
C2576 a_13643_18549# VGND 1.81f $ **FLOATING
C2577 a_12023_18543# VGND 0.609f $ **FLOATING
C2578 a_12191_18517# VGND 0.817f $ **FLOATING
C2579 a_11598_18543# VGND 0.626f $ **FLOATING
C2580 a_11766_18517# VGND 0.581f $ **FLOATING
C2581 a_11325_18549# VGND 1.43f $ **FLOATING
C2582 a_11159_18549# VGND 1.81f $ **FLOATING
C2583 clknet_4_7_0_clk VGND 15.8f $ **FLOATING
C2584 tdc0.w_dly_sig_n[93] VGND 2.04f $ **FLOATING
C2585 tdc0.w_dly_sig[92] VGND 4.1f $ **FLOATING
C2586 tdc0.w_dly_sig[93] VGND 4.78f $ **FLOATING
C2587 tdc0.w_dly_sig[94] VGND 3.73f $ **FLOATING
C2588 tdc0.w_dly_sig_n[94] VGND 1.96f $ **FLOATING
C2589 tdc0.w_dly_sig[95] VGND 3.88f $ **FLOATING
C2590 tt_um_hpretl_tt06_tdc_v1_10.HI VGND 0.415f $ **FLOATING
C2591 tt_um_hpretl_tt06_tdc_v1_17.HI VGND 0.415f $ **FLOATING
C2592 tt_um_hpretl_tt06_tdc_v1_16.HI VGND 0.415f $ **FLOATING
C2593 tt_um_hpretl_tt06_tdc_v1_19.HI VGND 0.415f $ **FLOATING
C2594 tt_um_hpretl_tt06_tdc_v1_13.HI VGND 0.415f $ **FLOATING
C2595 tt_um_hpretl_tt06_tdc_v1_20.HI VGND 0.415f $ **FLOATING
.ends
